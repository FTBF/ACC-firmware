// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:44 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DI3dNG/LVb5HLEO6UdaWDuc3FdnC6ZkFXlqyQaTyTdLOhCoLc8LQpePZr1uc4Jvf
jXAGusOpsjoc+G+EpxE6kpRUoNWfAZ9DNmuNspvoKXorP6o/u/Hf+jNLNn5YfPLD
vYO64i9kFCBZ5ANI6ynilUqRS8weRXwSmIZXPCc0L5w=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7568)
h4T1Qx6p/4kcTAH4vIaMaTOBUm1I02haiQoggHQboP91EgsYEwIGe4Vdy2FEXBjJ
cuYi8lSb2Sk7dp2935dRnHtB2DJ84s5n5kmY2dzolwCYFgP4EcHRyEdFaFSqcnD1
MdS5OCKFboszQxNzeR4ZVotTEjwUnPeiYnxGTvwtBFcaLOZmNvJfHB4zP1fsi0Ib
bmBICmIcicz6bvHqcvYLeKsLKFc2vUytDofp0g4Ebkso6Du02NQzJm/9GS1Pj477
70S7bAla6h/vQ7EE9Bjym7lv+c6CuE0Ayh145MCmO+Z4DVsdozayyQiEMZYAgs2p
S09l3aaF0zCASwGxT2jHx8Mq4Y8jdCfdCwFWOYMaxdirfqv7ZBfzARmffqXyEh/0
O8St+E9fMTVxzfWGWRbFsr3L+87kvhiw4H/Cs0AM1Qti0q0wEzN/vIx1wj1jDRCX
U2ul8n7kigaZeJN/mK0bFpSaFF0HAg/hYkVQpZiUoRsJpCbfKA9RO/UfRjgQP0Nd
CFsIIsLwDi0Nuu5uopSBu/YAzI8rVcgl6u8poa2IPznjC72e66xQrafBnOBWoLdt
oo9ioYzPBcn7kII6fTmqNvqEJh6Rdd9KkluvN4S58qKKy9YNg3d5GT23tB0JwEoL
wBjwsBCvNU8qPVBZ+DaRzp0NQnsO2T94OoB2Dd6OB1y5p9cMhfBw6avgxtTbZSXV
c7dIyu8FkAzvzIvgPHsZinHYDFL13RR2AVGHbJEzvaTn/4wi8JxjuOqpEQ7gOkbM
cETNIjumEB7HzsQT6/FcPnTPuor2wqgjO46T8xYPCi2dW1AFlngVvUiTnmvSS2c/
H+HkTDd6IPSf3f5xKZarhKmNDVAeBsP7FvVMJ5ssDQmV5LmNfLpR18lk/WGdOhI9
GB84HRo6YI8aVMfX6mcHYqKY+z1s9O8mzkwFqV5GPNYiyfxoLczPMyQOeLzz8Dxx
+3+TG+S0N3wb7AY7oWLDDHfgu974I6c7Ji0OgyCVOBtBFshAGAFYuVPui1WAR2gu
sdQcFH+sFEKU9yPDCEviVi8mCeddTmhjRUeWO9xE3vdRa44Dqpd+lEC24ROYADrp
D6Gc2QlHegRV1Nho5iDgmbZcOdIEFWlAL8GKuahL3Ewl2aYcJxszkcUfck7e6slF
n8y64HnETcCRWdmpIxNVP3hFyXRGTDLqBi0SuMsLgQMUJLLuXhEXCr+pC3Q5Z8aD
NOjve369gs+ww3LNAbvxxZXnVgFbWayIAWXvuXdLELncm6L6eAefPbM2Hu3gBcDD
Es7/XLpT03DYUg10meBSNQQm2RcEYih1sYbmlllo399NaWR77RwcIBZm7cB1W0X+
XgYG+PQfM+dyG3CfPFcLDe43NMcdbr8qVNqxJliUurH5ECghx0tq94VWRWzcJ9L3
gCEEHe3aMIriaLMVIgQvxfCwIz+BaGTpEd1wsmtDX8KsylFSwIIbpEKKzHAEfM0E
u9XZq3LyT9DyVs+RGWMHyuyNJ31NIMVINL3jFaAsOtp+vK8gj3bXTrN3gWiUJbwQ
Ug2E7kacytGddb97l4NFGlKjiSi7EtRQlnE/0e2KVcHWqEa9t0qOmChl+W4hLCPS
3CZ99UjUy7tt62tOS/8TpoRVSrmR17HG9c4rsnzL5qlR9hOByWIH45OBQQfR0P2X
Ly9OIxgFNzv7vs1Dz5235S5dN/WUNgwiCaj0e0AJRDQYwtM4sJgR8b2fdUjHVv/a
HMiqKZAOMrIwtl+wciwMearTYOgvfF+LZ57qrKTDmQoItosib6roLxfSTI0C/KgW
TThQVHWvxFARCXzv58MIHnS4wVCkx4dvAWLHSqwTYLrTwuQueWX4f04wdApdONuz
7luLyveFFMENFDCYsiVuBclYyaHN7SfcoMQUES9uwZ0Xz9wisDUBQnLMP8KxsI60
4hFhXaXQMQ8IpF7TV6J1FR1/gkYQyPNoJvR7tcpv9MzvjEp//nwQVRKn9NohOJ20
LzsV/ZCUgRZo+bRXWNO26SmSr3ZMUcxXYo//W7B0rN5K0WN18I6K+YUlF1zaoCQM
b496WiefZ5HrmF85SLzoNCRdbU1l4igbDTZ97fzX643TVaeFlV5rWYGJEIAZqcFT
TMhsslYdIbJLzec6vBTVmSYQIWtFF1kIdaEFTgza5V1HzdXDQKJ1NAhIbx4vKpSw
rQVlAecaLq4NPKVdwxnXHz3VN/myRgV2/pjH2VW7QVxn7qNJpvQSXsVIgjo3OOUd
BXSZ1l3R72TiQdjKNa5QPSobm/FIJJCV5+xfrS07GgGU3kF7BpyLM7dhSqk4ocWn
KlymRbQSlF1zStgi6xY1ztdtqTb4N3L81DlOsvg7+YkJqjsrNq9N+6xAzLPustVS
HF6l+t2MdNIImduW+MJqGf0nfr/ilMU7IOJE5iGqlrBEO6NSH8N9DvdwqrKyckMA
thSASWNLsfjk3CKpStEs1G8zjsw+zbRKctGHpdBPKlNbz5jfmIPEJxEh8Psdylqb
zst7HBr+dkE/ex7LoOMP2T/kj5ZO41nH+jmb5id6oe8h7pk0PSOBs+Pcdz1bK5kj
tbgDQT40eq74pcSSrnwqMu6zljtF5/elIRdGcW4g8I3hPT9pcUVdswCyF1bB2wR/
R0ib0DtEsWl1q2QWl7iBId9JF7bR3PaK4iLpF/4BGLo0AhjGvKf8Q2cE44m4dhxt
1X3mUY0wDYmyVyDoaW9hdg7rTIEPvYzeQ7uvsfKDQAGrQI1zAvd+zUREk9cnOYla
WMd8fn9oh1wHXk88yGvsRaMcJsKpE0m1h4Nub4HvQmem41qnxwKWqJh5j8W9ut2P
eXYWxWn0d9YiDKX9Fiz8/VxERJY40bYUp6tqirXosfYU4+P3Qy2bgVhQUxmKA1rP
pQaIXR9ARRR67RweP45gbmezjsb4atLPoU0PBhr+QfZLDM3Zi1+bsp0Up2e8JcRq
kCLnM7Z9sliy4FeEkzGsl/bYXHz7z5e8WZI7sYL+UQXaaJmcVRvy3QASJm8wPfj0
Ux8y9kHjvCwbNPS1JSxhEoVZ0akpgfHBFzfJDnX4qHK9jIINaoN2XY5ygxUiC3sI
DoqZjOP8uoA2KT1d6bjdMEanoVI9ofCWU0PcNv9ivpONIFpdoZZr0F2Z4hK10ld6
gcd6sxWl3sQ3QJXLytSWt4t8U37SavwS4nO7Kwe+PXaSxTmZpzohx3wzR0ZdpvDm
CBt74c+wyNJLk0MvNfTDX4cJp6ocN8GrfCd1uAzq67fmnrZoOuZF1R64l7F6MLOc
VSUjYA2ypsEHOEA6JXRTGuaGJch06ad3IAoXWx1klv+Yz7lQuVdpaNYAe/Snz8Z6
ABk1Tt/FRNiWlyOkz0IazlXDMPFOTN5mIk2E2hjUtpL9ubimv+lTpd/kxa2yt+Gl
zRxAIyj5McM/TI6euqTWlBVAdLBUmwRFuiZ+kNWisjww/pSQkzY4wikQJkTGyhE6
QBL82hPBotSiRToUAn82owNf8IEWQijS3YvFU+IXqfr929Xm5YFOvMWFQPY/0R+W
FO+OwkjfgxdHgnbh/FCYeX6N7bwR+Xl/+fgjUlEKPcbvBJbCDEriSMun0JSsoVrX
+qdD/3NxWebGsgl7SQlmQQXJHMszF2AqmtgWxq379khfo5NPI4QjgGFXj1uEA6b9
owMgj9CYJ5djHcGZ/9+xEj+Nc8RY13WyeJpoQhHgi0zN+Y7VJBzx1Umt6fdcT1vp
AERgWErSFbQsOmtFhXIj0OuaV75v0KwDhmLs3Lw2nhfqq6QTGr6g9veKTGjXvT2v
9ZS/Tl0HVu+uMBYaQDGiJq441TbxwTqtz8IzJNFLIfC/qqySsZmI3JW29lyTtL7R
mA6eTfEQfTv1b8Yoav0iXPIdS7AB38YmVZMMGiGFyW071agufV/Zo1Pd4N4pn/cZ
q5I2D/YsVZfg1Afn5tP9ud5t8m4Ds1pX+Ncfxd6xnyoP5PKycSU0lCIoA4etnhlY
ltbNQ1fmiqcWub1o2MZujlxDljRvUWsZCw1HFXbmkheuMU5OmP7dYVn5qqD4DBXW
muGnIsk3B+OkhftOuMqwbMTAo18/oTxZYOn73u4SL7O+CFJwy4fmYtqw0y76FRDH
9d6RiSqL2A6NEXFRyjWwRKYNo3NihDj5EeGhLNjjvy/nGk30HnlLw/Snb/XyHGGo
nGDdjRAwV7IKDP76RPI88ba/12768d8bChmYrM3/qsrwT2oS9MyNsdCgD29DJDgI
0yC6thh3txxK6oLG77Nw5H7GVUBYbzebPL231zCbErpAHjVLJ4el29dflgU2/y9v
sjEFbQgDzBTY/65PbVmTB4RESYENu8vXfX51OKEq6lt5/HbSHjzrW7hR1BftxhnB
gbkp4mOQXs9ku051CGJiovY0JU/efdFbVd5lbzvg8mrUo/CkAwvfS294E6e1vsxw
ucbqskFDxOyOq17ugeaugsgb566x6u0gpx3D6aM2dGJBJvGjxIxh0WVAuO/0zBJK
sF/bz46lqhMrz+eyNbtlki2BhX7n0An20klhh8FjenjGgsFkLEOOLixtMLMKCd48
c9i0Swh9sjgHYC6F16LktlVSW4M6Vbemf/7geoGuUz3nyJOWMUZNcqxeuZpxNSJP
2zYlzVWrokkAjJ2P/7cv04cSpnORLFRjWI3K0Dv2OAsft1SG5LRiORO7neLrMgGs
YR35ncF8xJ78DTIqt77Fha9FmEOgs4AVaJa3u9tDJLP1mXv3+dzXw838X9A2em/b
DVLCqXq74UPmtzVWo2sMCwvrcenhsAEFdjLtqO5Xb0T9cEoX+rX9U69MdzwduYWj
Lk0q95RsFOm53sA+Zv+I6Hs1XKeSAc5MpGQBUIp8M5ZWamKrooD3URHGwSHbczj3
opKq0T2yKv/YGrUai8t5L5C7CvMWVBvSdHy93K/1aOyxmmykyvVQ0mdcUPpumrx0
Ns/HNplKNna9xjDIjsP8TsOXaRLLgwcrpJJTbwgTahbLYDXJoe5npo45dCfyxTfE
YaakdVnovD3Iezy66CcxsBti/9ZKminoLpSjHPnzfftg469U8HdOK7/SEgfAWeUH
EWSgh0sSB/95/FeyYR30IJPtcBMWLKch/8yU3EAhHZd+pNBBmA2xWPlLC79uzL5+
Tqt5Fcg6wLVJF6gvMgK326fkpmiMHiVevYg+eqyHM+3pzzwo+NHsEdyzpQLpFfqj
qHHfcFfH/wPvAGppZia8+ggJqmi+u5PVxMdmLl3VsSgJfdvCDnhkXskF/vZOjcMJ
Fa0Vqz55Zxfb4xpqxGuvacW/mn5W81/zZlGOdsLQvEh5MSj1p+45mf300voVrL7e
xl4I99hLawaiCdIbXd9LKQ9V9Cr6ILbsme0Q0bPiJ7Lo3PjIYM2ECD8x20cNy2XQ
dUawu+uXglv59OVJBvC/rhnyMEMvDDdiPD/N32dZVnMX90lCNXX9UuJqzcYV90Zw
UPDjAymWGkqPa60qikiTqEe7tg5jleuyXfrkEar4I3MgeeOmD69v1ngGU35y2V4e
HWp2AA4GUgPQORze/tvdMurVGFLcrKchpv2EFcokiFmEAjqB4DOw3lrd37tQ5PEk
+noUSSerXE6R6BEKuEtTyTZUvmIe+8jekuJgcErGgKg+RTCnQyMunXF029MICX2I
S6+wRUNqv+gO6p3q7SuexWbfaS+hV3gw3Gzle84HZneEP0t4zc6Sv9ANLsq5qS1L
qQ9+RUJHvX6pkCh7410lZIjy6g73smuomV7LUxy5TkupLtmvw777ujVHLLtvqSdr
BxcuSF+nUgngEV9C7wP/8XgMs2007joLuEWYNYnKOc0Wqmv+3as5hh14RhU9cvrb
EiP+TCxJywcTFYm4Y2JLzPGAAIP1Kfe2kxPjwyCys5jXEmXo+WIyXFwaQ4G/kmZX
rkL7oa5Hs7r0V7jMEEMaNhLUTLnZYMAU3zIFjGslYGIjIbvKyGGaEIkNTCOpoTqd
OMBgV+z/Qg94CoNEPl9WldzkkWVswqPclf5lnz6eSa9HSUlpzc8yQQm5UwDv6fE5
6bUwFvfjJjm1ILV3n7TN2Vrq5NHTGezSBosxp2sDJevQlWOhhgJWx2gUvrQNEkXE
1jEGmckdniUPNiPd0Jsn8dMWbJRC9yw64k6Hc5SIht8ZO+dWNo+g9UynOORwdVra
UW/qjpHGaWSvTOe0aNdNfGCnCJdnGgo7nWzHMmp3/3Gni6//neDx/Swl4NQINXma
4mS+8InarjEArjhOfmmpSKuAXO/iM7/HzgY6mPit5IzhE8PnskJ5/Qs3gbeGqxSR
w/R/5dm9kulnLylVZTUgaWb9MOk7ZUqKnPehrJ0f0TOy4VyurQXhJ7BvLiANYxJT
oLJ3Wm5p7Gom+3HmOqQnnmRIQWAy1K2glDdxOF4mS2cR24kUoKSmYB4obcVwH/36
uAlYbdm2CSfpsl0We/i2FK5M4VsBO9lRPKd+V05/YLmqWgnouJwDy7wlQWo4eoJK
vXDnXUO1NSdTab7q9Iq1VXXtEZ/XQ4xBXfcvbgb2rCcOFgPRVzC4RiuJB8pQiUQn
e9MjY+YTgLHQgVuyHouh/OX70uS2NYMEvq5w6jKbSn84477wvxRCu2uKei4PTF+w
EUs44Un5JFcr/mmEWBUUZMpiBvf0n2BUQLyQZUiRkuQ3ZtNFXmJcSBKnocdkW8h2
3kFZgCaGd4W0MdnZ2T0KWbcybupIxJrN0ozoCyvrREeyfPCdgkGU5/mpytuz+h5B
3XMTRqdv+5uukU5ahUlo8DhZG6lcih5B+aADppxU0hTaKv0V89g4ndnj3OvBN0bV
C7OUwL/Ls23xNDyFMZSbrj+HpQtMKUU8MEOODoJJcZw4WknSn6Hhyapd7F0vN43D
4aej+PUvX5durwfEfVn87dwtDSLIJ6tSVEQUCmiUZShQAf4z5u/jbO7xREz6cSTh
jd7giNxaPWcfaVbvMq9QFnbBx6DbErU/h5Q/8/2N0L0sm/UggxojEQH0X1oxykD2
JD6YDxVaaehlJiomDBnS2va4sr9deLzYo6QkP8nM9EblA1WeT+/wAdZSYQ8i/gd/
BkpHqu+S39gVltIlbXx123Y0PHuP7QY94duR3yBWqicSNtF/yut0ucGIsVY2+wVP
HJKUMZCVrzKOR5OOMVuoAbkUppMmhppkneuBA+LkEocxsy1eEQkRG54JXQv/m5Gu
WPS0EZ4gg4mFLitXfvahq8oZ84KnsjSkI8YbHzdfQChrt9PruwHVfs+ker4O2LDX
ama/IYhdOAKxaW0lbMlcVnD4vWz8z9yxKzig60MSDyoLD1siDCUk2zS0PQwDOxQ5
hvuuYskst+ulykZmCK37shlE59wuQcNOuG0gtsxFLGyfPSsIQtOJkU3JynMf71TK
PRsbqAnNwYOtZ7Oemkwcinu0uZa1L+ajNKz9zE5h9GUWWqkegb7fCNu89pGYbj/U
Eo/ExBSc4eo3pNFX4boME9Lg/IMGdVwmc/VEpseaScfh+hmvMK1XpGSVVkx/2VLF
QMQbZY1agKNusIR6yTvWk5oXsJ1CQKipROE3wxav+JWsctrpyuaqVbAX8EdY6guc
FsPZyPVtzr+bxm4IPagtwGheBcUovY3kgD74YUNfyRga9ZSz8OYNRfCPInCIU7yE
kBOqpGUERaCnBMK6xwQC6QSJ1BMpt1x0HR+PdUQBBQjMdX7fcFYgbU6pCLWomxFc
jy85JXMS6IBEBV67914ef9y+VHLwykbTyfGVIVIZWvdu1v9/PYiFx1/HmkT1gxIk
KgHXAcmJM8NlJY3x4SzLQ7iSbYr2M+iB/hfgr9w5mwbtjfiKNJlJ11eVGUd6Ghrc
QOp+rrx/i38SY7fxBA8H579m+ijwpEUzw4XIp9IVZ40PYlUqOpORHPAnzLO05uPj
xy6Swfp3E4425r0QuClwnvdIa1tE46qDq8t2SrH6mG3hAHSDnHsagAyp2y8j/KI9
ZmG6TsRjPpbZsFE5OF9j1m87asEO/YvP952u3DW0fc/oFnmnjWJ3wMxEEVOClOTY
cFmFi0l1xVPKElGXDqb/4d+5yZkdjzCgka4TKdhuf4N1eBszHrODhCdoBpvAqT8q
eq+84ihD/INqTe16cSxyR2Ekwvcjmd4ptxDdCeJWhd4RUozLNOE94WVFsawTn6Dg
mqxOkApBC3LpcRdwI+603GIH3flKYXqJHKAazIxdlFb/fd7fnahkNsqbl0WTdGx4
HwXAIGF0U6BHIv+da/PKmlweQzeonz82KfHT75VhOPvCCI8g073q+6J0VYzan6K6
GQe9w63hNagzbYl/q5f8AbPnzwhn0gl7oxpXozTdDVV9tqREWbhh0vysUfQIgQxO
q91R8SxZWskI3XTL16blw1ovI3/Tx7WY5BJWfn/JDOQrIELpnIjoK0Edo775r8fd
vNGl0wlLfYPvHmoHSPb/VvAGXWnRVnLxeBpObl9QSITz+vHeIxrgFoG4C3+mVoVF
SYd+H5ZdTCNlUXmm0XxqllZXTdriq3W0KMnguT5WF/4yZ5rS13H0ewxbFkI6B3V/
1yMW4Fc2wvsPNc6IHdIHBx/uGdPmlNq2xltHga6xsD53c94AFbsCy73Fd1fZMfYV
A3ceDMR19LQ8r9iIfNppQ0Fk+bwz2n9Bjcr20iAHNvGTSh6xIles7rZCOE3/ND1z
oOej80GxEnv7XgCu+Xu38G6LsFLW2C4NgXetN51rptsdEC2r0n7hfx1PD0wsZhDt
rJjS1QV6SNJFU36YpDrXTIlEYqRBIIDZ3M8l2ulhyfKDpfDEyGkhdOD38PHcsB+S
s2F6RiwKS6kbwRYALwV+gGhN68dZI8p5/MC+JllfJeVciJdT+H51oWLZCd2JjGrF
t6rsm4AcgojT6NbzbSY2suSvwwZOL57G8rcfNaQhj0C2Zggf1mHpebGvmjhsdj70
WizyQs3Fug15rPYsKa1vC5Iwr5l6frNiksaSNVhKpXhYm3CCD41R06x4f3+kdD2h
Po/RUDjIlViGwhYfRpJpPVvZyfe4xJ/KOKJxfMkSRVAYsBx0x+TZsvXccYT/pvxp
gxGihrbkd8ag/RSfSaYvOPIxwz7WtOttZWpdmPxcKrVyO2eGZlAlD1FOPASlS10X
PMLRSXiRK67362h+oGDXAiG5QP2Q4DO1rF+pDUj94mWz2ldE7GijrKqAQ8INCATX
Sg4eSbhYuCW3y8EQt7G8AXLKQ7DT+QeTtYsN1nLKFH7jzY5IWrImTEtINP9e5fuU
QhPXJEdJzWR0FMQp5WkgCx1nC+ZfFScSaT7x/DHPZYijntqW10Hu6wjHd/4rUvl5
NPS14wD0D8Pbr1Hlt4Nfq83h2KWsxJUA6mTIS89VPy9P+RC0upuJhIMa+a9mzBqA
MvcFA4zmFixDtmRnzQWJ2ssEmwVHCvFHP0L6evRXHJMGrvVfpU6svbcnhcEaIJeZ
dC4i1rnO+HO3ZMawmoeps6VjqNKlJrZLcNFi/fC+YmXphM31dK9adohqiRuoblCt
aZpXZipLVCiTxeIwRvGuTmByc1dghvgAEwu0ZG6i1/T0Lq3GRYh2M/WmvDodlVJr
SXcXZQddiESIGYSuS/IEOSQALrWnguzzz8CXDkFRj1vBi4scfOkkYNPeXP6SKAbe
3Pz7J3xV7OKVVUqNkN1kskedvY6y8EvSfkA71/b1lbDCgbZSN2DWZOtD0k7F9pEo
d4Ha0QX4bXrxKQfB8Re2tIl8h6j/CnHNU5gU1xLhR57PC8dYbzbnZkdrbSDLPekR
1fOL0Z2H3qW4YY/010E+MIX1v5Tz6HbFSysW7r8Evt4ijSUp/7xMRdgwwjV9nD7t
w2n75IxnMaHacz2ZbYDVAgobdmZKeiB6LTDdoa/hpY5RXA8SrLkvbOGJOxbmQoE8
aMGT9u01D+RMGGtJThfhRSwVd/RlZwzjch5RP4s+1e4AFWOLDgQHfoBQHPGVz6F5
Bi/FwX4nRShsDTad95sglKMx+HJlXlKzRDdcVzK38ASmQ3QV3HfVYocEmtEsnP28
H5b4dWAevDHFE8RgzdXwDINsmUOHnlONVSR8WDBG5SFEW915K3nqrnP+vmB9nZnM
ssDqeMpNp6Go48wAMlXgW+CLwEI0y2zeC3/9tklO6DM=
`pragma protect end_protected
