// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 03:56:35 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
clwFTLeC/C6VXpZhy4HAsIjE6RmEY8gHPQdSAxCWgwKdDvyn3gBdi/ZTAUtPEe1E
I1IyuBoRjtJiSJTnvbv3YIlwoR0oL9yI7mIYzPnP7t/K7qybdpq2P1si6U1hhNtK
xFdYZXr1PmXE8gFAKU0V+/UHQSXIz7FWlLCUWq7Jj9s=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22368)
zpRuX6V1hBXwzhMOfKeza5YsZxv3k0Pcs3OO5E80zp1Em106Da/+6H/wHXA4wWOy
cEIqS8bcnFO2+8mxXWJphM3sKKukCVz1WFQG1XmyZQ7D0EGRCRV7f+tY/NJ40Pdm
37+aBXONoBKl7wJswHLr9h2BsniInEMU8stNhU1pYRVBd5Lu6ZXz19rGmo0QM2Pc
Nw56nMyWYUf+FX/GsHX0+knETPXgaYrtJ6dg0lgBn6sqM0fjVD67nKY99DiODg31
sqbKIcThX6HlXT+GqKLPeWwZ/fSNe+WtQjk4QzoUsyQ8zM7boNSKCTnPYhqMIlyi
SG25GvszTqAQ3jhCeiHxqvy7aiPSIajXH7SNXoYus3MiV38Mu4wV3W70wC3FfMhh
WTYIlbc9uRDX/rNbdm295g/MPxnar4/Yy+0TqCNa8aYrVfL7RX4IMajIQNQFlM4i
nbF0k7pf0XXKbtpr1ad7h3LlGFQCMeBgv5MULdshUrHFqaVhS3iryj9KSAgxmded
hl0vmRBL6iCYE6M7+GhBM2v+o3N5E9NzvXBr/VMadErNf4kN5964XiKN9OXUqhiU
TGBYtUpSZgrEe6xo7Vhl7K39EMBoYRm7BxyAMFSavr4GtpCRO7DyBwi3fPvcQXg7
B3ZPbcERVSDUDCb/LfHO5FJnfE7Ia0+hCEjUuBkNsT3OWjD6PRtleqGouv4syq+s
obiPj3xIxqoaz0+G12+C8EOz84hdT1YfpbwctV2WGfxkzLrujj38ECfN1WMi6Yjr
EP4wvV6KlNYJKuCECey1UeqrGux05g2BQqOXXdBkdkMcBHGKteVem6zoL438WU47
FfuOvgrRtKOgHffbvCXqHxbnfFc6wDnFLr0fsbnDbg+/rxZ2W5bm7cpkg+vpHfo0
emRyx0JqFQSDMInxlgruTBKN798EVbwVLMtzT38w7iSGI9SKRGjQyrNLzz/EvcrZ
+U3+riZhGjyJ5cfE94V1++Fj/Dn5i7NGwZ1CIzADqTIbzT92kzUaC6rY3nkrdVem
vpZTnH2CgPJ+3LHFlTXrpj8YHnIwByL8jrTN0T5j9iRYM2ODVnC9Ld6GWo7U5mKU
bzN545iHJ8Z5co8H+EdhZr4PsldGivrofs/6AtVGTMNilfJQoAHsjSYOxgRLfSvj
TbKpmFcAzxJ+PU7CPI74natTMupXClF+qNxQxDatKkS8eXRMUWDRLN8e0qk0743n
Ytmkw69dNV+xemh2kUUeledLq3x2bJezIsUSsTe9Wk9ekQ2F+OsRw25abrtAw7s5
/njGJEbbCtrWpAFvCtdcuEdbtO7daDkbrB4IMzH01vDdDfsMoASoFKz4tttRFpFs
fFlk2pdz+tmCyW7B1BM9YCkTdyjaYPdkHAZw7Kzm3XdjA/fKvCZy7/Y+I4JCbBsv
DN/+QlFSa5e1iqUgYsdGibq56O/6LXt244D1G5+IXzp7/YG4+VbtZqhaYzeiPRJd
ukzfYQblV6dtsmpoDdR2pXKx4MFazsG4ksD9XlWarjuD3n8b00bfpoNXc9OhB14m
Kub7VaN+2DF7Am5gtQK8hsXYhxLCTFMUbCEHHo6oSstyq4iWFgzwdqaARkG4jg6f
nCKyYHq6BY3qgiy4ckEkcTiMpl1IPi/u4WuhcvINaBockTjZ2ktG/hh8+qQ4aaXY
/aTXTr7AQeUN4M6PKNwqvkXr32qlfkmdIhYSayKRdUTzDGnYcf8K+z+ilKBVan+t
cg+nQGCdiIfgfa0n4FUKr3Qz5WfGXrg62RPXQ1Qf211RZ6MA3CeGYFwIgdZnU0RK
BuZ2h33ELiD0u/1oIkV10JJZhdsMf06NKM/xEIAzHRuu1dOJmucH4iszt2wRijX8
R3IpN5Jy1FL8x6iXXSo6EjJAzvMQqGLYAKyP/HL8hwhnEYXB81F4/tWQMsFyXIAP
pTLtGhd+BONXf9UMaaJSmbdnqpB220/+SgkyzFuKUGZzt8eNY7IDQDE7AuI7Uz9r
vO6T8Je3N8CuA++Gg0YvecwXiaEEO5rbV7bhNGOEYrrrJ6tmVC8SZKMy31sAuBdg
YhopKL4/VJ9DToGG53GHdD+qWQm4v7CzBN2P5qv2XrkpP7U3IzJAjIRj081SR/dm
F9tW3GYJEbseUgbt/W1N2DFalqyFzJQlb1v82PHnzwfxbAsJbu9dPGtlX+Js2i+K
H+JfGDnMWFCCGJFTJek5/TZukymvtZVEgDdlJukbN6xeLuI0y5bIDkNUJfnvZtjS
zb7qZaUjCzILhs2lD4QcZDzIbp/iEzC7FoC26yHfsmSkLaqDgJaglqbfey8rPbFp
GAXFHNHeABrId0zVO90XQ3ayTwLYYe6CPwURpHVd8JllV+vLGDdxzJ2Ay9qkZiGT
sjml+MfFbEPG0zFXplVV77snZEsxWgPCpD/zyYCzpiNy/ksuMkwly63zKKkcEcb0
3LpMdp1Q2GYCVZQvUB8hvbVqLE1Xo9QkkhfvKAP9nHsBW9b8Qfge4ULGck3WYVHf
7dDZ/GeN2Fq2hEd53XBYXzY2knrrUOmWVPxWBvj4jrCcSn/R/ijGG8fTDPYZVWJr
0VbMoUTczxxZxQ4JCwMEYKlrW558wdrS+azNpdeui/mRjrLcD/944R6e2UH+duIe
dBcy1q9dGFQoUjnbhLuOFtEm93zbtQIHs3F8eXJ2hytCq5Ub5cJ13R6YQtrAGFNd
wzsnSsZXyJjY7vMGAEtO2OyxC7GOctBnN6veQXQkHeaMHGWr3PGaRg1iUE8Nl0nT
oThKRwk1F7tPdRAFSg7VF3QRtYLC5ojBfLesSFX9qlV48PxSk6awwqFrDClJ0dzd
rgES+BH9ZKRalDMvonaPcjn6RfYG68s79vN4kbBvB+9xgiT/KUWzkXTA3aCsl3zv
H6qHeNrwdL7wcA9JhrVOYXEkhbYSEysC7fT+V/hdqzkvjshk8hi/Jz+JX2UfIPnb
7eqih5by7BmaK5fC3nzxYwZ8t5YrajFQwDP8A9Ekuu08rolxcvEmTy4rTgXgux5Q
zHYEETCMffnReiCzWdls5GyHFJ+H0F5QQRw9tPhvJivm1uhcS8z8w87b3TpX8E3U
P9hjJiZnQ4QyNUZuyCoKlfj/evVh71OsRNbuUuxOotkkDZglGcumOjC5YoiXwo37
nQi+owCo6eB2zVJbVcV1iw4qMOuRTgv/m6vFBZRAydgCa2dVXP8jDvILhLoX6j9d
FRu9+TeOdIj6pnnPBqfSFoIDn/Fe+e9ApimfD+KcACn9GT5JiyQZqjL1XpdaqnXr
EaMxkYMbQD6jiKdkY59JWiR1Bju4RPrzXuDOo20WSYwVjj/VoAUVNHR0y9iCva2i
0N+t1Ixjp2FjpAP9/ID+s20BgUsAvgWfZaPvK3r7ygVmgSrGVvleIHw/PRQFrwAR
qtqSAWjifonkbdMiYGnE/V+2TGyF1o4p+hnHqQJcNwUjALtap7NlYM8Pf8wsg8UC
i1+rsN6o795OYStOWFv4R2YO2gMVMYttdUauZPm8nmUvcSHbw3iJIKoRFnViuRoP
NwPzUFGSx+1pEazU9ZUQPzEFHVOp2Fr0kMnyZ1GfFZQWgSAsznbyiFGZkm2LwD5m
bruEd3wdJ6X4uC1Anos/hT0RmIFXEnV9wez8k/Da9s+rrD1gIif90uuMJ7DzYnLf
M8troOO/v31a+1HutJa6Zz6VibiuFMbOE3KCII8VsI2VDAEVQvckVRbSQwfBB1KH
xyrwb8Pg5rXm0RDgAd/vUNJoCfEST0BmdMFlOttbBVb57RJhnB5CZzNVZDy5YkJ+
E56WIEJtdBf4BiMyjfIkoQMsgzmhYNN1OnttnXKkm4VjCHp9ieVLDlv0v2Jpefp8
wvO0B4c0QZgm+lKOuMqIGW8BVdQG3fOPiZ+joIb9RJ+dL0ED7I5npsUY75Cy87xD
9TKByaX+5tcwzrlSIHDFTcq2zWdfqKvv/04IrPVEKnAc/qF48HiXkVE9SOZI2ks3
W53Llsrh+BgbubWdkrOjIOpDF0WM2HqyaRZBaEMYdvFwacPMypbykRlvm4BFmCLs
44m82xCLJp7b5XvJt1iif72UQP+/JGGUKROe/tiIS3ngPshceUvAyr79x/F5tx4j
XVRxGUd0c0kiRk0VAp0/C387YFQXGCEDnItl3dCvPXBIwA4zKeF94JFJ5y6kgjFo
WhKbkHaJqvgg7zHOV0OQNNy3TrYtJPZD+eCs6rDtPUUzOTRNLqllV3bu4148gSSD
voYSfWpy0rf0pd8Z4t6vetbpBOLwgbqsuICFKjEVDFZeO5cViheCebroe7kzM1VY
WGK5uYsEzx5Twmhd+C8Izw9aRN+/D/A78jk/ReexojERbesrVoXXXyzp58EjWO6W
OPq5yBKn+W6sZCiyQDVRGmjbiqHioVmByOjhGWZXIZ+QRGEKfMtIup1yuVirDVvA
t+un4s3ukMd5sfeHemJoCqBpOSEd7ZiEAiEmAw9tRJGgp1R9heXWfmllhXpST9Rd
COOzXj8JsRwPlsXcHcgspCkfvlf8PqYVKvVoL1EZVTAj5GPTThvE8i7XTwSgxJCI
OPPbOVuDR3+uFGEhdzSIjxL/DnSN0DUdLEawQlhR56fChl4l1TH6Rcpaq+ZJiGzy
+lppPOFdsOLuTYoqR2YNC+hnk1pFKzKZq1dUhKLMTw0JtNl/A/6vVMvwwkMHld8v
aBmJY2dZKmcteuRKVuZBM5cS0iLLG7j1p1zYyVRx/6aCkV4Y+GE7sTDhRRFWf9/A
Sxh77GgmKE+BpXn51859aVNAT5lqgM7s+we+mQrIXE1M1hU2RNXI+bs9zi6bBGmk
yT5jPDxvbX895+HgGBuZbxTXb91rO0VKsCWv+nznV+l3pyZI+iU182fgeRIc3jue
9YrwAcAfnLCKeXyvY09jrj0r6ptypGomPiP/26IyPs+Z4UGBdXUiH8bhqNAMMYHS
YPxAKWHYwG681PKLjuav7eh1HWumX1X9oHtO6cblqs8tDef8d2V+kIZu+Z2IZkvh
vM0dA7dStkjKwKjwtUtiXS30M7DOFWthvS6k4YA0HUIFoc+i+Cw+OVhlYA4zwJ5E
RTSvcq1f0uDGD7gwsQA+wfpljmzbkAYUrOV3Y4iM6xJUm7KWPl0VG6AQ3qe09j5c
5C2oQyoEu7TPkgjHZabAGIjCZSKZM1XeZmxeq6KzRUAm+/Gl6uSakbaKh5qhm9nz
oAdfcdI3iVBjohPoU4tQWo7rNuwHjjnu4NsYFXn5Zt9F4y/88CdzHDb7U858EqZQ
rorclscCaVy5tzowIHFr4BEOuCNfbc3+HNv7CC/1ly1bIpJDu96LpAJe8BYGQsOF
21lCLF/N48srokr6IolxDVZMGwn8B4wZFi4yv7MyaPWMtbDHpx4KcLgwSOy12u6b
ixgWaUKlGL4Uy75t+gjnpeeo40mRD21AbKwLJvOlBg04mRavK0d6RWmNQcPrQbGm
q0NsMUZOOuznfPO8UC8xpkoZpId0YlZ8nghBocoXLiohVs+Vhol/GHU6VgQsoJ5a
wrVBpjUi5FEm1R/SNXTGuFBN5HvFAjgp5/gzooUm7M8et9gUG04n4gWkafw7I9Ml
iOPWj+p8yxWCoV6tZGr/od0DUE3EImilMMsGtpOL6HorFbNilMQF5Y7D18uq0PUa
CFtcMDH1F3JohAQgdgSnc3egfwDvui2ww0Lic5nXsZ74Owbz+46pult6qKvSsWAx
BIjXr6uYA4F7im8vLeZwmTVIbjDVSQVoiYyZxYN+PZH+/9Xv4WZ327YobtGra+20
R9dLJygLVEn8BHlyhu/++YLMSK7pMMtOGttcqzVxeCCv5UbyrTptOD8QrCUKoUQM
YZ+EVqRpwuPzpkMybsJPYHuASbvXFl+5/JCMTSf/1zNZ3vDR54gGq7vNlocEaZfR
DB4NAGZAqakder3EZ8ri+pqgEvg6rJJTtV+20qYT82Nwct16ZrW2Ice/O5kIXRE9
lHZW1RMxELh25kq+yKW7g4p8lXJvEbjl1tKGJQucwaK7pg2RL5W9KjJZiZAdqtuG
JlYuCRXnJUXAUMEzXJXi4UQXg2at1OQxb21XeUGzgLB5sHRmsdSjHIF/EvpyIO7f
2ySb3wt8UYjTmzf2Kr+8bKiKHgyJvXEgDHNhQ/RWuWu9SVPyS3CXV2+j+WPHd4C0
7PvtamLGe0dOWJhSJ3PVjZPYrwD+j8VL5MnpItR6KEG86dT+DxOArPfyEVBXmjvy
v+fe8aChUyk2qZNIcmDXaf5/tKeIZKecRTfQ4LeEnhub/MLw3Qsj01AD+dTH01Rm
qe46r2eG37sfR3IwfaAX6EZ3T4V52yf/IGKNhKI3pojQWJB+peJEXDW8TCY/4JBh
Re3cCCS1225aBC/dNLHt8aVAFHYAAyBVbhx6W4RvV7WZRjgZtxycRU/5iYkVEJmd
hyYQu8x6AcE23djGPlcI1J1P+/E6RqlZz4jzuIYtP6vdk7zYs7LahtlyWIJB2aD/
Mvpo9af5EWWaVv4Ycfv+JJG4+MJvniCdsQ87lerY4ZpptMwhQ2zwqaZc796tiD6p
kYDkImQPSzP4cwuNqOQ/Br2y+Vvgh7aHMzkqPGo3aUMwlr2RwViZgEfK9BH+PvI/
XnGdHP1I7mzrxtWJTxrWYmekDoHRz8+vmRZaXrhx7i5c01nJCPLtpGu7fzr47PR2
pIXCh9wTQjBsI2EShUE1q5lHeNRYwKj2sAAGQLgdQ3Xan8YyzaJ/CpQmi0OAdrzy
zONCGYlMPM2lycmpvSdl9Pb+0+T69v6G+v2VYt8zPwAK8rWHdfpqn7EOXzY7Yl+b
zTEGYo53A2sV1FsNUigiltnWwRqBjUkiKFRfR0Gk5xjPjDBF3J/AEsUuvpNCAt5l
K6SFb9YgyqqynP2wGyueAX+jZRphnn0Z0CoX9eblwXCkUhahlztDp+Xv2X8V0FrE
AGl6GrZjfWLV0nGztBU1xOHs4EkDKSBQMIJHlqjR1JQHls7TaFzgQHBTmN4HoMwq
nn2xG7eN5DXmRLRDV9d73aEa7yiWUCVsN5ij0+84aPdLijz33OnJz93jcaYJl3qu
D6+UTc5EfMMoCynOMsjXj/LGI4Ipwok5nAgEONil5ymq0sVBuNeueY5DHuFfvZdr
HoiHD+jhftqMK1psi28f44vGlHlazMQ6XLUwBRgD1HU9HlH3yG8iLpeoC3BykLXe
AIIFz+cZ+n566xVT5lofhblYaV0CuDUGu/TMrjELBQQoO+IPDo2KBgb1rB3iOM85
PLzW+kq/wJp9oYsI3s56Bh+4dIhGiHNZu2n+WHAZyYhmKVelYnesmji9nKYeWyb8
2AcCaWD53NfT8BRdZElbIKiEqC7xpTZ0GOBNIk1SxvUzKBJvsGlmf7SkmUvSdQQ/
3YdtHY8B7xZyseS+ols6gUrhu77xX0WKxVp5fHZpA8GXBDHVYDHH/qHM8TJbu/zQ
Y3R/1A77XoxN9XoqPRSNXtZxSLYE4xyOJFW2KadZsf4vnO2tXJB3vizBqX2THgzY
L0/bfo4K+I7xuEp0DGh3b6V6Pnts/7TdgIYvA8K16nPeOen/lDN+Dv+fOIod2DU8
0ws+iFh2NC50Dz7PTPguhjwn8mbg/RTX0bK+OUY2hprBVKSTB8Q/uV4P+E2VUt2R
Wy9VWg8KdsErSEn7iqvTzs0hqgAm9uz5XVrrJVEl80OiW/wMJPDNB03lB9HO1eAz
IWevnjwTdTesyG7A+ErxOi1c7AsG/6SuAh3EPeJVlAnAhFKzC/T3t7GfZ1rfSaZa
Ug6iVjOreP0vktw8NkGfvrxNlXprbxSwLoddGjKsKpWvGa7HKw8oQCtviBxQyZI3
dRRvzDmr+iUQHe4SeBsKAAQrMOfY9P5FQddk5h+JdCXcav+chi1X4pjpNmqzdNsH
eadv7l3iNlsr6oMtVuQO/R43Mwfx0oPLdQpYlisRTwZVtuZrKZD2/Ibc4/a/1/+4
XYvdllu03XEMXcm0wmq9jBrdxkKh4/C0u/dInyYPPIg3hXODgs4Cd6ZH/yzaTnkV
p1JC+oqi9khMQ3b/vAlt8ykcKDhEwQLwO0d5haIcf8KiGmLqSmepBl2oVUVXhRA4
llrZqHOksIST6wuwWRb8iIsQfYagrLpgzsuq4hXMaS0a42UeK9w9aorFp7phJOeg
1/p79GRm097exCWpvmjRtEep64OWZBlT/lizIQzGIyzJvHUraObIPFWE13hy0lDI
9pE1CQYTWdVU9OwFHVLlPBKFo42vnzD+MdWXGMljQp0NVP6wqqa6PA2cmC0em8Om
6lqokvaK6PlDoLO7TIOOyaUzD/43BBCHNvot9YDyU4pGgJNDH+7IFW2rLtDKJRCK
zm5EvxqatJKjblHXiB5Ue1PtZTlb20XevuIttUARu1mfepkqt+VlsdYmzPwfJkOL
pgBuzzlRXEyk5hMezl4jv2c2+6vkN+ELdr5LaDEVli+igeDrl7WC9OQpMI9Us6h3
e34sfj8NwroJh5T7xpRWwxRESs5EEeYGQYcR01rIJGO23zeMqPGIFIaS9hKYDAFF
7Ddzect2FrG5+pbL2SDj+sx/p8P4J+u1QWprMvtg9ePO6UnTo2j+0XVzsaDYO1Ng
eytYzARBNS9SXwHh4YLU3qKoQCVvhBzW6eUU2LH1b07fuPs5FoJKqtgcbyf6Fx/F
JqZeQ/Vcxlu4ZzOCBgKuaPKBIbQgtTIrwXPsmdbkBdDEiLifYe6lBrUlbslwx88c
pC5tHXWPN9LGVrfL0NwsgpLSSes7mV3ppzsk2UqWIY99m+XPt5BpbXOsZgviNjPF
Tb7YVruDscQPQvBu+vgdvxKbtnfHYrjq6bXCl2SnGwNEFCeX/wal7hBZHD7mqytD
AY4Uw003RFBZfM7P6N6kKo5Mq0inKyycmsYyKtK+mMddF3VNyO4deT0tyFXy6/tq
1wbIa/cKdNODpLeF0ZgUqX/QfG+c8zXma7srDsuzUf4n4+3fGhjNC1R8UNo/jgTm
RvoMP8lrZleeJCc7g4agSYi8pwOazxwUV17dPZRe79DjL5jXtDCyEl01KEGadZjP
xCk9IjDiqOk7Zc3LXLnHchUXi61H8YJgPxROvmdQHLx01Y6HynCnAOcJQ3OQgLmy
g/jhcxrlkbMlhsjhYXP2QNhsmxXm2DUDauYBgbinIf/sJYHgmBqjHG2+sO0b96KM
3NoJIrbZrzot4SHw8DmOtfYTQFHGn9cJOt/eqdntA8Lijd4b4u0HL2kfoBmjBqB2
fpMR06v2UToxPUvdngIow89PIKI7TRsdVyXKYNMhF74pPleJ8xpJBMrWUQYT9LwI
r+mhR9qk+AGUq19smpeKQFDuW7N12gFaf4T+RFVGdmAs0tcxSYzCs5HVjYwnCAxc
e37+RaZ1eVLhdeIANmFoTA0DatU8vAfKFwS7I8HCBxqCe/OxBdDgKXEig+PKMR5R
KNB3rRwUM2CE4c7JoRHWkxMkFRaoTHQlok9bSn18KDSPZQIhQQPJDy3IRTF5Bge9
+TnH3YpsW5aY0cFkdtiCYW9N1MgitQuFqNEP4vlyCqnCUthYuVusBb3JAOqaRFPR
KGINZatrSCjf3BTslA1DH4JxP0uJOb3dzhAq0ZCr7NivaRdr+yRi49iXCqqdNvKe
wDoiSme+22iUq0ERpwGP1dx4KcSN9t8GwuxbefTQcw1zx8rKJoCRLvFNMkrGDtU9
xQ5XfOZ2cLB66p2MeVad3/wdvxs5guCJbkE1Msl7t7RiEQSNS5rgwjq+nRuRwuvD
fKMxLlwpc7K3HR+vsL/JZTY8GfWQLaItdNjyWmPnWuiFovALN0W/HSlUMGVU23cf
X4CKEa7KIa4+RNde8AwbMQBeIOk5gvE+tRlSIpq+vjIYd82p2zwNgidWiMbgbNrm
IAGZYW+cddbm1ZQ7YOCcnYHRlXhNQFcgxuAA2XwO2P47pieN9Q9T24vXvOpPo9K/
ZUoihZyAfGpZFSd8UbEBww9sDLlUrIO5MD/u+oknXWZ2IvuY5uYZ+ubHWz/TN4HZ
TnIcYcf7qISU1kTMWxtkE8Opkoaxs+VdY2aw0uEdKooJkMb4T79bO8EZCHZNRdaY
VMNwQDjCgy0gvUcZreQtEjPcS496pUkKpkW0Uoux/fXNrqGF3Qd0fbJBUYHGO2fI
KzCzLV1P+FGyOrmeSMUS/cZP1hecGTP74STYkAqcYsj6gXosn5mnY8bnxqZ1Zdut
evvDW0RF3yok5c/8xJCXXKb3jMrA5EC/LxyppaaFkBhCMSUapjeSAopdWDr540Iy
urr+CawUyJj4wIEQHCOVEVyQA1IyK+G0d7PNcgqcJGV3dfmeaRLwD/GYXtSVGov+
Q0h7zIfGoMESr9WfG06gBl0+XpkoxlioBGtCpBPqDlpCt+t8qplcGAKmx9WCtHKn
H+1XcHxoZULmfHPM6B15r8Dipn2GK89C7+sU7vPphbTQk3ZseZcVLtcAuIbzlok8
Xksp+UGdkHRdobbGyyEeQZu0sqVGY70w9XIEy7RF6qwzvo1H9GJ3+/2Gs5Pl0Ni7
W8V+eLl/fHkryH9xmtew61uALSj117yfpoGy4BCnYQ+cv+wQX2sPkit2EVdh/Yjv
vYQxuD49ckR7rIf607K3Er3dogjHlb3tT8V05dLpZrzAFbIpSlPY4Dxa0SNqpS4W
hQuIi3LGlzQRcH6qWOxFjlLqKsQVeuUiJUgQyKO2HMTzw1OX1qEaTq8UzE6ddRUx
+fj/dLYMZ5BtkXLtQCuXDp0WXojprtd4XvXlhngBbSxiZUnFnpCkQM2mYHbIsXEy
cVwnAuA8HEPVnyTMybeB+yWBuMqOPHwRXIJpQyGqG66N78texT4uWVykgFoZ56i0
5xMRrgMbYt2OEFe1/H5sXCJHbZOenVIXSt3B8ei3jgv32ia+ijE9w8BoiSMJj/Xw
WiZ/EOzXsXH+7nNnbcPAi9hSjibqwdsWMa5KHDCz9f8wgcacYBnOLBCCGMrEuoeQ
nGWKuikkj3OOuNcbmCbTHsBbVpM0hcfjT3sh6OvDme22R8RSRXRx4anfEGHv3jjv
GJNBW9uv0NSwD+Q7bHruHzCbdS92VXUoDhXh4z8aD/StYPoVZblagJPxjcGC4Ico
EnQVwPACiWlN9vRtOUeaDhXmbAB1HNYyNO6fxR9omxLBlpFIH1RenFVh65r2SQp+
93QyTWqWTfij4GKjbGdtetY98skEzUK3zegtn9IH70AR/6ENo4LmlcoFWFJ788KZ
XPkHraH4LKErxvwQovsMkLf51KOSMz0U5S8osbGz0kieLILxfhEfrnfMuy6+KVrK
0c+FNKSfPJaMOM02kCfakmovf2efyqOecohQE06Cc7i5tOaB38b4UOfx/y3kicLd
5ALfrcDyA3SMm1Uut8hTZT0eeJTSbTQNfeC+Srgz2m4EOZZFMHo75BK5or/MYGk4
K/aBDoYqvPz7gBzK31HGNCyrg0yAsWVQHjepG9sYNzGyCgtPpYULoc/smhhuW0oZ
V9dMHnHyV9CtxNE8/J8GFCxagLULAnL72La7RnqvsqONstHzqDR+FswLwrLxen5Q
fgpdOLmocbNQErF9e9NtulGVRSwnTuxX/dwyDwrRebJvU8yn70iTTT29KxuWcaQq
AM/vbPyfdTVqfyf8+YtOw+Ta3toXk1qYG21X2dUL+EwvBp5kAVkz67kFhfPPSzKd
l6BfI8s32PQsSGsNtYKwMo+H30Q12FChPtg0VFbp2HmY93OF7Jj3bqToC2gdLrMH
xPagIsODTEmGo25CTN7cRRiQvjvI2Pt/d2cXT/eOO+wybv3lFEulZdRGfUZAq+EI
vCljef6TcD+aI7XauTSOU+abVqKcSYO3a2+hC/OWvNXsWJvVd9hM7/EYjZlWYJza
gHZy4YuSs9dxT3pmIl0uQZjKJs7HzZskQXzN1U0ZS04EyxuDsjhh6Ha7IwshEB5L
XWKYMJJYy7WvYqQKfH12u750ZkCjM+pxr2e9vQ49pGhTJydtTPnKojrl1futce5I
J/Kchdfnt3KJtQqjRssVvfQVIsva20t8sIS2dpVmZDYMVD+umTw4ehIZjJ6gFzPt
ah1FUb9TCFhSTh9WkB7qpaRj4+kauBOQDup9b9KiafqMC5iafWUXbMQKo6aJo3OH
weURmtOy+6Zz8YfNvPgumV1KDDIsDTLQgYeKEzL5XWzlEZCkh9YcgvVEnYvbUb/D
McyljihtPkWDGUmNDAJtSnU+Ho74q26Jp2ij+JxRVe0nPgJOxliousM3U9nH1q/Z
aznTbYXP420/Ydg2AKgwT96On/kg3xTjamI7BU/lmE6PAIImBWKNl4b6cKMz/cwJ
wE1p5FHC8GLgOwEejbyqJP1mSQQUOVzUDIDK4Q4reNpkEVWIBFdobeDaxbCz61p/
OT8Vx9jF4ElpZzophmoUqWUfNWJpHOtzfHhwg9UQaa4xvzB6Fx/hyWHCIQjnxIT4
Ww3oJ6InHmX6uSEo0jyg8AkY3pShgHUxf0Zg3vAOTaDXfa25fYvJQOyKkoeGnLkh
Oy/uKxICbwi9qsLe0gnT9LnOfRR6c8A7krqbFGuxvep0bZl+7GMqUnsG0C++z+KL
bhbJMrH8HVhPYO4UxzihLWsgst8lbdxyyfHtj/FTXEbvVqfGUKN7xhL0og39wNNL
OqYnobP5yY2A19Aggxmkz2tf4gbSuC60qpEZXzwtX+cNjVqlyD2byQmGies6AIZg
vZEvTF8YZr5sLPb/8mB24ulr+1FxzKYI+7eSM332oJ+itbtKZPewVzCQxCCFJx83
h75Xk4CyqWmDuJDVorfx3brGkIQfGBq1PxJNFImJE/ldn+MvsmJ+jDnx3GiSO7dt
WTHDhQZk5XKRGlQslV47yIqZBqjBpl1hVRg1Pn3UyR01TnkXrNbmPjcKRJcgMXBB
UXoUNjXI5brV+vKjYvIg4krgrCPPeIQ+6GdKEUk0gGuC1WreESq3g2n5m5BipIVT
AlxLCd9O1EddpYISEeEZ+mC2dIScsPFw/TzFZLOi6Dswzm1wjVzBmwwBCwjk3C/s
YS2St8FaPkYEfRNZJNSygr9eBk6xds7xv+rPo1S6PlklREizrZzg9E56lYv/T/Mu
x1whyeFy4DXc1JguppFG0f7atLHEAuNqT+tkpViYnUnsbuH4yMRF8TXiARSs6Zp+
jc7vYLTentk2yNK3DtBxu4ZqfWetm6B7bNkKoVrbWpO0GiNY88Ppgw9QnOt3m5nQ
AbN/t4THkJURYuJJBTjQv3r/y6aTANi9DY4N6ZCHtckWgPDJSA1CblAvvKwspoGE
FAm+NNSkOtZS2fX7+JEbyPIjxnlsejtdOMg6T++SF/X1i7O1noOjeegALL48NNBi
52l6QBBOcbeYZ4u/5AAxfg+TA+InbAHynn7+8yQx4BU/MWuXFN/QB164MRrJ8sgn
iNECN6/UTqaYBNo3NlCyK2Gfpb0UkilCQit+nfgf0gpCk3zHNN55RaEotadBnfgs
PstEnRvJCY9pKgCcYGSc9NGszoq30XM81vaClAPB+z1Pxrp3bQHW/VZldAY3f7iN
5dC8pJLsAgrOLWFNkQg0L9HdrKIysjJj09NAmm3KCISCRcOPQbScf8vvZpJj3Z9D
ajm49TQCG+RBQU8nVd455hmGMHG3dxplx3ThHVGQCU3qq3e225I+7nIUcNWm6cxk
BbyyYIaWMfiJe00ax5Sg3XEKZsDiOq7YXSaDKljFoJopVLXq69yX8wcuQ2pnjB5k
lBW3pDeIfWtTz3I7mq1gl1KvgdxINjem3Ml4V7n8coWkJKum7PvZsiJFbPAwQsYO
C9gezPOSPf86QVISLQLpc0SroC86Ksn4yP0SV3OKMj2Hg02FvDimw1mdClfkumtL
e5Uf7VPltirtOkbXxMs2WYpLd1mq6aJIGW19tULlokP86INQfdpme2CGK6ir3A+j
CxXac1M2H8j384FDUzJwBzOiJYW6fvmjPpMtIBoMNbl3f8WUX03HMcyYY7tE0lfk
CyIQtFNYJM9wFSpG8ongqCylg8UfrR0lLt9roNkWvBLgqLgcPIZjtQkNne+Hg/41
Y9X02s652abwDmFtc3pJighjJ0zLlsFXaPiQrxEvFgkETWyeMcJi+q5WXhgqzGx0
qftQg9Wiq6N2OJKKJysoC56+nvq8O/8Db3p1z9jwxkZw0/gcUMaibPrtdb50oEhL
H1YfphqSD993tGJZRA0t9nBw+93QQVyZTrOO5YdRABefR6meQxWGZZzHuvp0U9zd
nmCBBvXD1LKsmc/YqwrYAZmhmu2NC18pWd0n/IrxEwxiZcop17MI+4waxiU/9dgI
soHA9EpbFMvlWlyZ4VGTWnlnEVtCOEMobtfN4haYORcjhq0YAu81zMJmPDdTMvup
E3j7V1ZPQPC4ku8W53zE0ZKDb8dKJlW55Qc7kNwiy4coaoU8YePu8FDKjG6A50bV
553nnmp2tlc2ScbKXXAlpdmkJszsWG7wnV5IP1gDWT4ASa3UTLTWXzxLzfjv8lRp
fTaIjGNAfskJ12nqnB1S/xFs+FL5U3HOfuK5TPMqYq73bes/VHUdsgjXNuyL/86v
SUusiFxhibKoKHHeRIU1z8o8RH+rjI7QFc2JJmLVclF09C1Rwo2MZNiFU6kibVCF
H026tHEwJtCyiRGv/mV7dUViAqKcCklseYdeV61K33zP3hbu7xSVIH2gSqDpXFe1
nfO+rzVAKdJLfut9IEy7QsETXAAHeZyvbrWCkpPEiTMAdkrDzU6r01Z8JMs2qs/O
hoFF8yA0mqGVmjrmqwwMog5VymmrwOF6ZvQ1dmYsRBkDnRVKVd70s/KtnPQbQMVO
tioAZYBZ1UplnJSLP6fSoDwLFkhGm4viNtw8LtvMmn1rLd83jTSj4+ZUG3OXudBO
8xPdFX7pemsa6Ju0qcauHrAeL2FBj9OZF6ILJ4XdpfVITgMSNq9StIr4cS4Oxhu4
f/RVSP51XE1n3Nb29PQdc56lEMgD3pWMqdTdITrcrsC26GveUrVy37bplq4tPUfB
XAGBr5mOFIObfCGlBayOtGhaAfrYGANjWVMCmonSZeKwDnrizUnx95c/srQZ2UX9
iCX9ukoa32s15/CkYgq6ZAXYkhUtS7oycHBjoU8HzJ9MFPMQqKDuB/ku1lzZJ7Uu
ipv12vRMItISHwozMJPt1Z/Vb5LT0DpqXSCrpvhSo6ucm8SIDYCH0eDufn1TjHXn
Z5iCBq23eY01woZUIBXUGrJfJ1N/mvoV3+uOvK7To7MCjrS8bj9078zolQRXIevh
L7EO7B9UED7UrH9+6JkFoaG9fyDJFxo45JwrtuN6RpsgByNSfFGrCfkeYfW+NlVE
URYjOxmmsc22oz6gWyIM+WWESBn2bIkpHniYM5AmnOgg//u92NTR+XyzOE+0lEai
4KLQHU89vVmJB36+nsJpS/7jGLIFWp0dllaxpLoJkyipyDwVYgFQTKx3fbEWZ46o
xAiiuBBI8CM7Idl54eE0zlLqIA8lDI+KicZ9l5kaAB1a2R6wRVYDkJqW0OLgI26J
3WfQu+weisG6JwwGkXYRgRBL4aWzBVQhNUrLNPeZcnL9DYoYNRUCt36tLnz2ff/E
WdpymS3TvbjkeSl88DMeNFSBy2agjgyN1vlRTsDoR/T2WVP04uKM6q3tZHJ6OHra
a/Oc3XRPo4Z7f4V/EB156UfpR8iIQrLBtkdlcolxeBVRNu1JnAGI3+tH6jpiIzzb
AuIDxRgsdURyPzJYVxwvWfF+VmMm6gBs6O3U82BH4tGwxLCMGBzcbWtjwwBfzwcJ
yzM4Wx7mlq2T+q0s9r4uEoD6TP2yAQEC6AZGSxoCZf6IqOnBVb4E9YuPaF98KAL2
UhjXN54l1auKTfV1Xptc8Cnj2e5WJu/TGlSmpmsvFqk9IcV+PFATqG7W0hcKu2mV
byMBBMjIxMdGNtyeU0FfJq7ZNne20D3bQcnaGd+S0SRlIgzhvqq8GO74HVJoyO32
4vlAdj7XFjh78nPXoLt2vsaWb59uF7cmvIs28iOqgZik7+21ccML5WO108/HKH2C
5jKr9DYwzQq+Z7o7jpfG+SEdyb+KfySIXuQB/dE9ymmOf8txlxvntd+mPU4+OtKi
U3afnNVkBjLPeVG0PpDl7e9LUo+P3ZqPV0IprsPZFmiBn3EywCW6/U0Y4WcjVxFW
Z0gM/HyVGuRVR+cCMdoJ6214EAcxnoOzClqmOhmDLwPyMmbeZLaRWJjR9p+thbal
wQCl6qClYUqLLD6VtmpnvhIBeBV+KCTPuNC1t3EElX1+3tw9MEZtSemizNcEw0u6
ApfYTlqLJduN5RL5WIFJRL67lhfS3wnSKENy64UCv9Enj/PNNn9tQgTWB634SeAE
ZVu11XZ/m4KA70fWo4CZq3Hs3KBF97KGFJ3cUmgIDBX+8wxEHYhNvVjD+bF644rc
b/Qq7d5buwz9Ku9ijqOtddNEOQjFDG3ktdLnsvvhPOU6MFh2vfUu0iE6fy9xlG18
hkhShioMJ7AVJ6nO9jLuxQ51V//9A4FJQ90jsN76BuVgp4W+T4XQD30RZnaAacxT
KzavYZizXGzt/jJ7CUcY6Ic+bAQPOTSLWoRKMU0wN0WIt3KmIpXBzj4fvk5o/2Yb
FC9CTXl2WSOPOXg2Vg33drZ1PY9XvcfjPE8IVgDhOfMkHktQnQ6s9iXPuD4qf1pd
S+nRX2UpiJzqxk03p0K8inQMfn6SOrpELxf0cdOf3OI0Xq+ugrplHB1UBdVBsQ3D
MdtZpwnc4ntNOnPIJ8XimpYZirtwL4Z7x4oHwFzWSmWnjnFSoQvq0D2cV8t16Ib8
LEJUICs4RRHgTdPYRJ/e1QukzZXTnqDLeAW7M7p92uNd4AkuAyxvfPp3gzr6qRAc
COPoIfs20OJouLoUKFtldUX/AtPZyZOJPyj0K+vc2FOnHMdxrMRD3Q2jcQFhH/zJ
1Mg9eR81wPUQ0Kf/EjWeGguXCS/0iYR+s2H0070EYWMWpis3iBAsi+hK9EHu4IeL
vN3bJXsoa4SLtyd3Gdyc7kqe0yaPe48+2YccgerKWAKzWxU/BAoGS3DzqNYcsG9S
II9X+E/GzwY28tFVwYg+tlgwLbWHGpk7pUuuEMuxGAon8MeQh6gAHaQBsf9/+a9S
OE8P40LawrCPsbvFP+DH4psIPsXCEGvVJmNSVXeY66IpXA/8BxZuwDIxUvT1tR2U
l2+BKoG5ojMje9XDErCGPlsInzH1UGzBe0SJbkJnq4Ujqrhsf6LpMirPQ1bqmwyJ
SFPbWPLd3E61C0qL2g2g63Sz3q7kBM/Qa1oMn8tXaUrpUpSb34u9LK55d2bWM8l0
+fUoAOq0a6z8wGdElXe4NLei7j4jTEKNqHfoHDovPDj7GIRZaBQuyaYT0ZtkwA/O
UOOZ2xmWDDyklwCItolr4oa/koF1tlkh9MXISt1iaGfHzHqBcq0BszQNSYJxO6oH
hznHg4N180++cw/VCeKcm4V+84qDo3tt1ZKJm4w6Gv7HkH+UxPdrh39X5kGqlkLS
aXpz2nrTw4sz/f7ppbVvxbm2wKUCUZIXy7xZV2MtR5H62J/AqnXr+RTZzIJHPzFn
GsEfMQDxPuROgGAKs6bg5Gk0LA05uDRHej6T0ahyOHCaBdILJHZvDAc9plJSCoM4
eKQ9uhJlSgYtwDCzYoF40bh6/scWqggD4dS1UitooRlnx2fwLWRdaHPsSduw8zTk
V7A+lliZ26JSx0s9HOerjBcR8gb6Zs9TAS5nXIVmYxfD6lRMjXsvz/JTSLPrxCmp
dBO46N9gJxic/PqH2nM81bks8QDlHCm+Q3EPsl/QuMYqCc9xzF1BgLTJL5xeaJRl
S1qM97Voi2SO/xtr3Oahn5xOebZta89VOB04hUXuyIVYcCDouqNY+X6Ha7Y4ko5s
rhlsGrNgwwaXUkdFrwQ0lPAvzgubJDOxgujZk5tpw7Hl4g5+jz2xhcA9GN71OMUu
oikdqwJM1QXhmBQUeXIlk3warn5Vfgvr3wy//PpwmD73L/lhoCZBGa931t9g92xn
ucBCAZl2AGCHa1uzVrmAvPXRLaLW4jJSQNWsPuK85Lge7VB73faJKxppBATJAIOn
PBUtiDBHtQ1eW8MpzHf8PNotXdDW8uvNXhbz5jGiEKYoFYsvptfkYqAnR1xrD2a0
du4TbRekxoF6PTc6JcdHqgxgKAEXR/bK8HlNTHoGdkwI+oU8g20kE1mLtLon9+Vx
bzVHMe7b/eQKZgFCZWeS1SsekERCOxES+2L5vS4lhvcCd19o2p2DFFDzL+NM8jv+
jf3XDG1uiA1qdRw1t9o+lxTQ/dLRZn+dozoySBx9HY5rQNS1eVlqE2be60eDgA9B
CO9E/G5mbuWbtAR176zkkJUOQfuOY/GndrLRTo4sD7UUAUN8PcLS5tDGDj3RMskT
bCADu1iztZci4uwkcu0cK38m2+i564yc6fZK16xz9Y0DGMIihIbQEJE0p2eCYjI7
mH4Iy1z1+BIDI+DaGMHNwcGSgeN6gw0UiMa3eH5RM8gYr78c0JcpNwPOGkdCWQ7p
Wc49UE8dH6S42FNw2iyON2a7xa7rFR+jkwXnoXEVvDm1De0OqobyTkWmI9vjoka5
WfhnnkbegyZ4zylXxzGGVv5yjCvGdM2F65LKPajhL2a4UqHflFpclZsUB9yhhg5x
fu/J6vPw/rpTEJGgqG/uBQCmkLFWFmJ4y+t5I+XNuYGkVQ6K8bc7T/Vn5W7nxTYr
MXoMscTLqm08xJPpRCMLCU8/5Sl5dONZlrVW5rrONlRckcsN+R1ciSteK5g7pII/
SrU/klMiNsJf2CAbq+M6oUmP3eBmNWrAjUSuPHDTnVeRgKmCUXCpUzV1XOVjJV75
xFKKeqKMP0uiUtobE6gSUJNo4kKsK4mdvCnD7XVTG0e05+WK8LVn0O0731UqQEUB
ojRe8zt8+7ZR/rIIDFKAkZzbBCdxMCTvVZz4uLK60G7QJheAIGQtNkunaa37IuSW
N4HzQ84N9LBfRMwkB/MqIjFJLKdG28oU8yqR0JfeRGk3jgaHGsonnjvwkCt4Imxa
B8fRaqQbw9ysQIXArSaFKeh4uPoa0VxnUVxAYHyS9wuQGTeEs62dAV7jVKdPC45L
prRrxfDwzk8DmnKPVpOD70WPita6EE2/zUTP4WOC4zriW2IvzEBLLPaBqtVasw5v
jWOQ29rxorpoJVdj7x9dAZMCezCyp2T97s7yG6VKjuWZo5FddaXmGbpkwll20DNR
htS7ie6TqQZbh9iIMBk+tApYgM7F3yzcviF2tTsIE3hmz1T86NL/kMCeD8gHAoiB
U5fHq8MinKvGC6mLRBWuTQgisMki54e+OFe4Nadm41RdmdJ4ybzq2zzQwChwS26O
PmYE69fHJniBDd4Ibl6kLAXk10qi006ZuVW7q66MNP6XG94t/CPXR4PS7LS3RaC8
mW76MwwObXF4eCHDJ6lGU5LuARMw+KGuit3Sb/iZPyNynUNRPkAw9CgXwjutqazS
2hf9MV1BpM3c/DL44p/uAdcWffYJbpnWpGIZU6C03we5DhXmQQjKfRBXFTPQxZz/
9oA5noCPfIjFk1OTQRJE4RL4fQfQM8UrlHihxx9qvlmJogdDMZY5B4i8BKmosI5/
u+CdnyWSHjQwIL392P4RsRHcPrs3/vahYeD0Gn3hMHltO7swjZeKr4yGKgt2cAL6
PlNP6LWmS5b5+ZhnKoKOALB76iJEWGfhg9vLN02DeL2clKvuSjzTUpYO7f4aFQq4
MOiwZYSfAFUuKTUqeVJmy8iiU5QZBUgAa5vdolvrL9oxrvsOI/P+nFjCLnDSJWTV
WbYDbeMxv6xSdzPuAxAWIDyzX6omfjOpPUT0AYLhaBAfarF78UjQQivMcqPqKHX9
jdSdtV/CGwvtazcoTMFZJx8egwWubkQtp10PBCXfkOvRmr1+/U6A9slb2LQ5GPK8
uS5hXQnCctaul0xG/DBbDlof+ENqN2C59aMoso4hmxYv/5+x5BhtQoNM9asvC5qW
N9G1QJLYOQ1eSaDG8yEGz0RENMgHdCWb6loyvNONvkCAGAwRhgNkliYby/5mxfLT
XW8xi7CU6hdQydJyuaJCpfhDlIhSkA0VuiIdEc/z+pDTfiF/p5le+pg3Ub0beLFZ
FLJ4YImDd+mPG48V+MIU9G2Gc0d7SGceBodJTszeCEUahn1xkmMGl8CNtm3iiTsH
EeChufSHnumGjUryaOr7HzMiPq6MnwnAQcZcBf704iimwTP9rd4BvwTVQBIN2LQz
09z88qdx5MS4wbRpaR1s0taxqZCW71DbkzgEk8sMMeqJqLW7K9HUIqAWu3lcZ49n
8kxi4Sr6v/JbbuRG9atq/GitUFx8g5imGx28tsV/+VaAOCfL+XuykZkWxKaqkuZu
hOliTEEeYcOUCuxNSsMHoVNlHXg4TNeSchDSwXD4S1E88xMXlVoaowfwVV/4OSJy
QPVcBQ/wOyHDVHz85LiieJbuMOmV8c1s9kbnPkE6nPzYhgbZm8UTxnCLmSDcJ+vl
dA5j3H3bhG5aPm2zDNKAOy73cexr/UuxNDf/EmVffhUHikNz5tqBQnzT5b4PvlC3
tg2xRimTPzv2SD5zr99QQZfoXsPvPDpZYAMi9mqYAyKNNPJP94fSBkRW/bS11k/z
FnYaIUEVIFtUy/pW3+0ZQtWH8AAgbIKisWKTh3LL4c5Jvhs0deTecZfZV9Mmhkst
wvwrdsNUKI7XbgM4E4F59Qj2jF+t6FY8rts+LP085u/4tVIJCcIIw84qIEXSsHho
oJhbYd8+enRAHoBWpuZnnvfAUTd5l0M+fh7BWvV3saymLrvnsmWvm2yBEvORQ6lr
Jo60RtMbArGtSrAcIYW/gUTCUzPgpmvlrCE1w9I9q1I0MV6O6pnYYNvyeZaVyU7x
vrF3tNJTMo2YjFBzlTKMOF3/rrBduPxlXYDXCjo4DW/zozbLIycH6TRqQweAxQ+V
JThPgUYvePjHxSo1FOmmwvzHsYGkrN1RhSNVJPSwxqogx0970vHEKBmLxHDF3NuU
CUGZp29npqZ6fFkb33AqM4f/KM0T9RVmto8lvoCtdxlTUTWaQFi4SQluPJfKrEoT
54WoXskeZVm2MrEEUlmedH5Ryzqaz84FJBa7EQ1U9M0/g7jvjpvaBN/MubE4JW+f
ZsDldoI4LmpfwhQ6YqA7PiC7ghPn6VD9BJymYV3Xy7IE3BNqWmUGBDjEBibvD7Wr
yYVuVLbELV39a823cKM0i65INKqDojTXcI1SGzskiYcSBc6HsitKPLyYX6tZPnSE
0qj0oeED5HS9+J0A5JXdg0xdetDxV7tMQrVFhkkqAJuCIRq3MYzRKydWJklFe4pA
WSnfPpny8L4Yyauh5RvBMWdug/yKb9dnMdnOV8yesaTYwKmVrM2Is1eDUK+UvXp1
YcdPesPyPSyo5/eoC/jbmTjZ2On3sUdqU2bMBgnYTe13s+pa/rsZt21wyrqrMNQG
QiGnJVd8aXBAtN8Tzqq3Rn9Ta+30mj7iYA2IFwQCKl+RnGTZzApPB3HsQkCe54Ku
V9GCalCDnBvrIfy3QDQe+3ywi9ymubJf/lNseeLWlwS9ntsJexdBblKz0B4g9t1k
7L1Y+kIh5uEuKSQoFpFFo1Bz+TCgvVh1ZoCaAwnAQJqIFQnkB+FnIi2xBw7nSWo3
zeC+h8Qr+cUdWKBDYVd7U/vQ4WZAcDtYwopuUnlcx4rgdUzN6TkDd6EJ12tS6X7G
3hS/xwVuzX7s6xboB4tc5UO7f6QW64TYj2W/H2OIYnlcsR1OO4L54WjMsWFZWUK3
HHWDIce/7LXvE+GCBp6XVUoljPzS/4iYp0woPjuya6ithiX7QJEDCURgMRrbQXES
wMPRGIMfybDVPxhv10jSuSwq8cfTqnL9saOZLNqo5zShYeoipkp3HUJ3P+nhsEZa
SO/gCyCahIDc+y7zdk1gywKZ70Lp6fyQ+xjNvbkJcXNCNoOe3vT7zxF6Wn4Bu6OE
UUvfzRzSATN0WRd2FgtnU6VPYg4DtKb2PcukHGWOEvLQRWCxUKqGbYfN8Q30/CF4
8MCJiXOqJS9Kwpelp2UNAvrPHDXFq3r3W11VbhqQ5z3NcBwSCgY/kxCjfiPajB+N
/3DKiYJqeIIO2v5L2OnTM8urV3t4GZXoeJI9RyFklZMdrhY35Kivs/hNSxx4zPLR
QmvhIde2TvWUNExWh/hqgIEFxM3WVM8l728jcECRWvqSqHAsMxYzoV95cGvpeC+w
95FjfqBh/c8GfNnpA/TXoosFS5C21CQYQ563fCOLwYlDPmnujAWmAOY/d40BhsvZ
iSjgVhNdx9c80ddymCSiJBH3o7TIuDe6mJFOzxCsGbqRWuZCQdn9CIb5fytFOwAz
OGWMn+Aqt8v5BysgZLDQK4N+ac8n7S71P65KoYYpMs9cS9i0H3JgdB5jyg0D+9eD
OApfsRlFXH24rqP4muqYpaOOUvwfFd3MxrDXTkffuIejeG2W0q0QYKX2LEUuMQh9
HfTjVcyU/lXtpSlQzNYAKLw8eiwGbOMPzDghgwvCbrCCH6GZucZht3TuvFzKG3rh
GmSiOTcAlswi+RnMwjUgiYZdbP8FLKci4MqKe3gDce1UU2D2JxIIVzTMsEiisfyi
xz6iTwOaTfo9GQGsbOBvOkNhN3JAIasrKZ6bVCwjJYYb3qLMTqew1G4fpCfZA09i
etbW8f0Lo32t1TdIfnBZqcvvnr0uVvrjoXI0yydI9ya8swqWbNBIbFA7HAFXEfWW
osQtACvYy5uEdKvJ6hnaSfRD6rjc6/4sPwGoe74l60gd3REYe4hkRRNNLPKSxbbk
Mt/lQevmeYoR85+3y5+4b3Yx7MQ8qrbXQHuHz2Czk14d2Qs2tGZ8coJP9z79rfff
bnYMsvPuQjiBdR7ZHdOQMUEDFR0vuCzx5ztHN+IFspTobfQmqFucn+o01UIroXl5
vYlgPs11yLFN/uC4QUGUsC9cF0Dsvom8+W4jjjzBQcT3srdr2NpRPqCPnpPr6EeJ
9TeFuyzJ/1XwLZOR2KMqVVmlQJEX4txK+RxZw85Jk1iSueMV6XDsn/WZDwgC45BL
JAJMOHcdAlA5t8jtH7fHpDRBoLLYYqNAOig2HRBhFFS0wqMC5DjWQW24ko+QaPZM
IKN/hpJdgItPhQHTnqECEuA8XTm/F+/jbgJBOQGnaNM3Q43SkaFEaI2SYHu/Ls/g
ObotuGFapeoRv6Lfpin5rjor2XC8JP92Wi617nglFqoHwWQX311n+Fk8bmRP9uWx
WfVgIEaROa5J8cV6WAvVhWY8HhNr6NdadA6nZqZLzhT/5ddp7y/xmK52Ph4trh17
XKXwAJmLjsDaJDTBP8WILydmTT8L64tyPWUIsR9TR9w/KAWCa7SV2LrGBmGmHanN
Y5UsMDGvu3FOB5TLjULqlRSMTGVly5B97PutVXYGDsxMBfrTArU6u7g5vhj+oib7
DbYySjZqj9iFZqjZpYIA+txsV4g6M6gl/nz9UcX5pQfJIC/EcBU/f762qymt2vIA
fQNmgtOB+O1aFb+2Vhw4WAiiyHjk8erhoFYHZowYQtjewnqEZSu/kKT7+QzclQGj
V7vk6e8RCPIZ1G1zAmg6UlLuy3nehPBWApVuBe/6IYt2K6FgdFuGusgpVIpgaDIN
5dZQXls6xvv/xbgSaGfK7+yPzTRaS4jL7jAsUu0NnuLIks8+i9YTkT8nyogVVRkf
FRix0sU0JcnzgIJ6KheT7LZIxDmMv3DvSQhkq6H2r+yPfH5cEliBCbSZOde/wYVs
MpW3zc5ZUrAkF2G1QipduxQVXlkCJKLantouvegNcxwodB3aWYNemk9EXuqOULmq
gKXiK80bR9OLORkOlGIGZZ2d9C6fKJvNtvaB8JMCuazGjFlTCZN9Rbv+iz4gZQZI
Zfs0+V7gK2ZLbvBa6KEQddULyLduCaBknszuYY4UsUXJO1oEie/7R6uYd8v7GdEC
VoTFExBKJ1CJT2LPdYvSh4ikjdFkj6csj4YU/gR6WfJiAwrfDn3gr5acqZa201t6
tPuvooyZf2a5S+AzPVoSusfZGTPoJvwu6My72KqKVbA3mmbRKX6Qpr+8Ap82tHIC
hzghYxKl+QVcPItBpf6nxxG+KchQ6KHMdLL2yNtM1VgRjn0HCoUEWz/iErDkmvnT
TtsovZlxzhIBuu828L8pRfaWBwsxmqRD715bJHpS3QC7pcgh7kzOXJRdZxTQEDmZ
WIcBFCZkSBoqat3Ra4mDr3NDLIWrnWixRA/CzIGGdU2k7vCXuqlWWfqqErUglU/s
lj0jiMr3Cn9Gysyys/Ondury/FRAXQYfD3UoUwUFDrsE8NNPZgFI4Xu869x74Rrk
ZI8pUsYsJ8zknJeiXHSuFC6FBt+CYf96Wn3Yht1Tt/aLlkAllE0IDG415boN9MZP
BcKf53+7pif52Kzd7mMKQ2RbjTgF8iEgLlpUJj9BzgHhqkA3ojf0oMzJ1F1361F+
BbSLhvy/YRsLAQY+1HKRwdNohDbuDr2MNSpVHIgkKTUpkpPa3DE6slPAWX+Qvfk0
ldcjq0b+sf6PlVuImyMMeUnhyxqsig1F23IogJ+bSHTe3dgoBD9jkvgGZ5G/9ZMn
fgyMeLxIuIuA3yU1ix2WsEZwmzqo14RMSY6RbtZk5e5C0NMxZFKEyJQwNKovnVED
eLNDOcftDxZtWT+dA1Sc9uMUTo2A1cQxzfy5fybIm4UXk5CQEsu8kp2I9RC2BykZ
UnG30Nxd2ZYL9SFt/vkiIARz2OzIjdIL6GTZdFkwNup+xP+8yR+hFMpxDMuXIN3K
4NKsHTx/zv6S52UgQk0l2VKuyK/OcwpvSBoKCvZSn+hIHmh/JjSSyjsM72YyS+I4
NVZytqlTI1Woarv1/r0k3vPCKkUI7bgd2w9OuSPN3EQftyUskQMxAFIUGdG3JvQl
vBfk05KKgUsCfnXMStkh6yXvGoA7ArgN5diiFPNLsfe1G5OAv6ceFT/EcwQzE2xl
AV7j4nWAj+VjMZfh/i7ZP8z0+E82VizP11qOh7x3vJjutVzrHBTmT5iCtsZUocHP
1fpUoIx+hSFMqUwbMdqUE1lvWgkjRyc+5qSU6gDrJwB/R41KSDs/L1EsO9Sm1FHQ
QBSC0I8LVEPsSNmvDUuQXZWEFFqpoeXnRPIzw1E7BNVoxqeqK9jz/+hGtRoyxJjQ
RDv9wCDbUFSxyAV8h9W0fZRSKEzgl49OQM6pYxSf4/OfLGx037GtBSN6xGa2EzRU
wuuR8qKHx4+cK4fMtqM0ByHJXwkU3eexMPbwsEZGgbLSvi+x4ShyH9Av4ogt7VQz
gehg0BP8ZjIE2n30DUDNZ3WhQOlZ+jdn61nuBBJMmNy38bS8yOBHAdLxnvwhruD/
/aEy4oGW/kU8T4426Ol19ex8RP4yHbfRwitHFq/kieaiUzfnAq2YWZiV1BdkHwxU
kTlr2v39zOGrkwIvxE3KD9kvAGIrg1coxoECy148O6tFI7p/F0qbjZv/5V9Qgchk
xEh+UQnwIW4MmNldFygzCdRhFB4RvHoZifRJTeNjGy+cPpdrvRL5rwN7YW/yTlsC
ncKnJrokSFEwvGrkcn191Mf+ntLPVH4VADaWTVekm4jPJUabU73Q4k+FFmThhTz6
RxRehEmQr3DYJJmdU+pFpkMIWabUmEqCDjqZxPBh5QoP+wCEgdr6p+DKSFZvNeFV
mywoqGt+WrFxTuQrVgj1EUvl7e/kQwaaMx5kqIZD6dZG4a3Mvp8FXE3cMy0RGQnK
j4b4rn7x4hcCfxfBvEVNutk35P31tgYOtcbQjkcxYglngewW2bJFU/TJ1UbXSMO2
Mmw10L0qRbXI5jMUyvmmRygFDfFtghftv+fWV1npxQleohRNZ8n2Lt4pCW6XpeMR
ZOGdJk2SnC1urtGlg2uaa6U0YeCf41mUqEcnwG+465YvS4JqEYz5t5BHIGBWyVXN
UyAMhANVcm+FR+hEfgEcLKj2vqm1vjbmZCzE8LaFCip1oVzWJcOzyG/CevtP03kp
NltigRjAp/waIWlwljlhIiLmbuDEFtzygsqaTgmLONAlT8X4wjREys4JWHwcAh7I
BRha6F8GNwzYi+CY0lroyzVXXhDTJJZAzJGYHHAu8B62p7TUBGjFmx1x5y3AvLMN
NEltJ+x/UX9Wjs2yUdBZuDbfl/LSqnaQviEgLnzgPJUvHuuzCogXo68xTDVg67R0
isqUnIVu04YvFIfT9qHATGvn+ONqB2Remzw3zrLOQASm09Un2IsodefGxXZ9UAoQ
TKiRr2qu0pzupCdVVFoYZOcZK9KOUqQ0GGfM4kqYMYXagO4Jz/ZneugrktfYPHie
eiQDp1eitS+G+ZPszR1T6hzk5w+I+bLc+yxjSbglbDr4ZgykGQxJQEgUdElW7AN3
EswTTLUIyverHW/+5m4zIFOFQFsrsZ8N/XROyYV9vegrNAsbook/IajdIAO+lzz5
7K2uoNh5oBgrc3Qn5hZdhdpi9hJyYMf2EfavlITpwaPUCoyf6qxMguDW/xHSijq5
S9GxEEN7HYlIxy7Z/7OGznVNx8YxzjBsVe7NjbiTO0VXB9RjZn+4E+8NvLmZcmmD
I50Hh0Z8GnHJoHtbSh6ws5BbXT3bAq7COgc7VFnsu2+apN63VPph/5LkkCSUuomr
HRno0yXxhFK26ouhyaQKxvpuKNdEVHqXBnbKzg/8O8vWxARWB6K2K3d1qfTcPtM3
OlCQhnyWvVXUkF7ARNwoRfyjWGy4bb7JEFr7aThgwPkelTlqt8rfFbxuF0X8WtGQ
e2tvHah4YGzo6z1nyrhzb3Kb+R5VboveUla147u8kMNc2lBjfYejMtLSeYk7Pl+Y
ISQADHXdh1YUAeoJsbx1Dy/LXmDiyU0IPcs/ZkM6ZHtBM9Cgd95Tq2e1Vsdbs5Tn
cqEQaUyX+26eQEk1dmawARXWwq4RAkDAE7nMQ2f5ClMRWyQp/2LzjV/6Csi76m1b
3yiOuhN15hDhaDbrfrKiDShxGfyEFnUz528hsMqQhCROhChXJ8vH4yDkZTE6clch
ugmWTHOXRbXDtH28LtpgOR3Fno/oJfGh+6TCyiHLL6eFo/gdYH0uuqDHlzCfA07H
uIVAnM+sVrVfMIXjTAJKukBzYDSFd6cNKs8l0tQE1qA7Gi9xnDUqqC6/g1/E3tR4
LKWz0+XI2oZDrUhWB6GD3UflCxodNy6dlNl9cYpUOmOrn63/q0EEcCTHOVlLbzm8
ZrSmlgqbmUNrjEWpZBt3a4sch+pcODGXera2RjQFZdCPIAxJXJ8VzyEXeuC1amuV
+fDzfqJqWTVaefoBqd3QVmjzqlOAPRbrzYjNTZrJmAr6BcRCZzwyooHdMq7utQek
WczX6hwP+kJxVoFyyXdvzY+plKZmfa/59fZJL+sGihwIqVh4WjbpywLH02ARu3Kk
ZXI+WlmIR+J/DrkAAWhUzTzFjV00lLRtXr1pI+Bazvpu6qlfbyrdKbqbssOvf5s6
rhsg12Zigf6LiLtyV2zxiIS10/EC+zTwQj3y71pWIuHUT2+fg+OtOssNrSBRy0MY
n4rp/mkZqFS8mCAodlM0XmKho8IXP44SMJaEzlo4TTQXQQs0AxooYienedyQv9wK
Aid9NUeXVG1Cq+8AuJ4fFJ/ZF2Zl1PvkfkDVX4P2otO0OHpui8gbbPTZluRC/9Bn
xBECpu4LYIrIoUZ5XEOjSAuGYdBBMxQhcH/Z9QZNDAL/qESO3ggKBB3eriXDkhvl
1oMQM6kzscLOqyNoXhwscS+sb0dyumEC/C31cPpnNSI6PpbMWc2g/ztBNwxOtlCk
r9n0Q7sgV/a0hrQYX9Rj4dlsm8zfd9F1/Cjdhhs5osiAcHPQolGzNMKzTOEhOtEe
8J2TNx0TiIcEoRrKKXta5PZoo5AtSTEPu3hvaUSbNqrCE2HCArIRqDEpJ67gDLCv
6yI/68ZVsY5HNiGUuuKOpxJAlVG70a3SoEWZquTuz3qC6YuI5jFJuMU/mytJcpKX
7zCp9UcDi7001X8nq7KF9OoQLzRx0qlSWNtdXbWCjzgdIaKz/JtYi49uBqfpHbLE
kI7pQPXAY/osvM27bdeq02EI8I5i4Vf9kn7Wng19g+JZwPBMa/YkvL6a8ssP+oFi
kpnTr5hhpBsMIgIQMr01ylKhpDx6esHPtEohgn2IFr7h80t5Il2WUGUYws00EyJp
7cJqG8cSTl6VEDFtqVPsgsxskknlAgv6eLxXz/7KIADMz75PLURFUEzeOLUT9qQM
TuhM5hVKaX0qOJMmD1vZ3o6mmDDSi2QtAQgw1cXqO9FETxo5BrfhKkSbsNjkFwgB
TtNxZ1WLkztxk4tkWOni9n19QLznnUBDaUKhytEVSueLQplyQMvCurPk7/ZvqEL+
bfY4dguMWUOjeZ7WKMF6mDlVb4cRbc9sDW/HWf+7kezxtc8EURxb/wDfJaZGBVZl
TDArYRB0cjWHhYH58MzvK6q8r979ozb5BhbLRA2ENw91alPgk28ra9YB0QpVoFvO
j4c5raIi/a6JMHxIciVzGXxS39qUM45H37Ndt+/TKMzCg9fc9fBOf5/WHehH24Ml
9lSUAlXjhrV+3aAaJ2DyZW8D27q7vU83sk9JlKofJLmR/45PCamjQ2xfYEm2WV54
QmyAZylUokLukjUerYPMZEkOrmtxyMT4HabyshqwIxk/RlNllaPWS+I7tvOD2VT+
bYU+HlRYCgS0A/TrNuKfWhDtMWt0fnUmMwszvGcnhuhtbgwkwz2eFfvBHdBlOOJ8
6aXpIa0sAYLKEDhfRroYrSIngLQ2yBcBvHasaXUPDrgHl55Pkmas8LOiMPOWMlo2
ARqoOSXZjD6FG8ceie1I07LjDPCUrO4lqTYVyEOPQlvptO8bwp0Lv31AZefM/9nR
XhOgFKJqOITEx/qnlN7sVUv/+Xc9wJSgUeN/AYk/VXZlMjaciVYGaHshktMHk1zG
fH1p/WGqf0gTkuV+95YV95Wtuo7B6H54VE5K4d4xRIAs+jABtosMJEmC0VE9gfYK
C81frosatoH5e7vhsztuCfkzlk14paywkvn1ep3sgC8eeDjUoCoZ4UBgrcRuGC55
D38npfI9Pp37Q7/DsMsDRs6IteAFDM/BICDTw1Ax5xib10uW3jW3vunOtyM/gIAu
QCrvO4NiZFLOeuQ0VACa3wlyemxGIQNhz+3457i6rKVvBBV8I0nWVLBN7SuqXMd0
cJ1npQO0u2U487rdBNx6zU9Ak9oP4yYz1Jl2XnHKcPbEaHX2l6l4kPaKZAYg1mEI
c4skGDNV4pRzOkY041HWOlKOCYpxgf+yTOQwQ+Dx/WBgMWTKKj70qE+ktDn9agol
+MnvtsNxz2l5LazjRCE2f5lUdBdSq7wD5vHgkoAwR9Um/jA95z1ZlLzrJJP+byU6
5cUh8aCEr9ZN8+kvPHeTyklDF2mjwy3ObONJgxLO6/DaySePZsB367RHzXwaRYad
t8vZufuxswWgpvg8Y4Vu7uzsucAYbgxjDBif2t+zIjOWQL0knZhvAQot3a2mlX+p
3fUxmJ7DcfVCIL98L1gGZTkvCP5zb5QBWhLzqYvShEWJYjFz/KqhGI+9uKsdJkyW
RRwkfULad1m6f/NjELFhd4Vt59Y9d5DVwrKYKGGcCjkN6xcq2GRyHQPP9KoTqroT
ZgN9NQm9PLnej1iuZd4Q3PDRsl2+OIww8vjktZlZY/72RHjm+zDmQpeneIpAVHD5
3A1S3X0qRd/H28RfsYnHcYvh9UGld4Z3G0HSLt0uFVJ24FyVDcQwKJ9LI7WY72GD
v8RGRaXZDiPVs5jRNeUxJeRQPeS6eES04Gje9X9m92nyagiVTIZbZrWyzD8N/9MD
`pragma protect end_protected
