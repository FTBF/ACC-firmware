// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 03:56:41 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NKLX/Sz9GuR43eC2uMmxrqGMtkRqT+m3chem7/Z5MLFaenKe3w2RCEpU6OopcXS1
NIIgdURt07G2/O6DNKEcnJd/h0TMfsdyxx2WVfnrOo4jBnzj6yudu1Hj+L0uMStz
gc/W3j3K8PmJWm7PWMGIX36uInAqPTr+nAsIQp38GIc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19936)
t+XxjHHPyr1eIe9wXZ0evvYvUVsGobw65tlJNJWIUajx108A/ma5024b/LY1NfFN
2ndwHfMXaKrx6EMHNveWU++oAv/+owwbB6q4DBmBfbSE0nh+lM8p752HKLxNETek
ZFJJWCcautRVzNj13TMdnCI2rvrjWus2xMLC1uicxYYJWdQe27LKohcGmfQERVLz
YGbMDAoh9rTgieq3Mp7yK1hAIxOThMErMzDf7izWOkHv/f9KCDSOAxroe8VMSY21
yYIAAKRU3giHKqRRln9OpmCqmUBrJd58yATSvw8N6reKOCdNF9oVz60h5xdSj7IM
qYE1xhZvQGoDELTXv3N0Rz3IQJT1Xm6GdLAkkPUZD7iguDW9oIBWZeE/I88WnLx1
nODCxFbTxP30oFxrL1ajHXTp4DPxYykzOllIrex+OfkbV8yyIVY4aA9JXBwAqjcU
5P6yzCA9QVb53yDAZAql9c+U8d1Ua44/9ZSiuJhZ8dhxMYU8R8j4+0fYSNpE/Dhf
q51pV47ucHcr1l9dLsJHHboHsiVZfh6xooeLc8vjHpmHhKN6kHe9jxkizGobCxW4
SHNn+FzmUWt61JtIRdHUEk2dPyrYklwhRj/doDUd4ZKThlAvvvZMYMqhygkDIAAd
Yxvwy1n/Kz1h0AMDJg7FJhSfEhhseFsCWowCYIhJKbi9kdzmKTqB8W236nAq7p2R
GQjsrxECvkZFOX5nqHNgDM8FRG7bOFQsdA1KCuQPMCOsNFcdtr+ygl/URVYg1QjZ
RWZo4hI1DUyCKQV3iRWnIlhsrmn34e8gfa7FQSU5qSa1WebSoTbhPQEuag6jxyvK
EYq/ZzPk+n2fimPVMSQ7mpGS5G0BlBgxKJ18SgDrxw4Uh2OXvhTJuanLB6EYjXc1
VXLrKqXBnY5o5xvdII3CTgX4a6C+CNKZZYx2YAuEWIwzRVq359AWBFJz7ynL7iwq
1W8pgrXHs4nUaVHd8cwtJ8/aYeUKYpasfGyGZ7c/qMp+2QFNmqHQClADW6W4tr10
AqLKNCc+TAm3k6KpZWh3tfxmFzt8exOTCMGnhmaeXpImk2wmWZUJOmiBd78btxK8
zrzfqt8+qFS/oK8FnxwrU6B5Sm6nBr2R1N4LvZryeO7iKyqZzhKji3gG5URREqSw
o0QeOfYZzr98FuTSgCN9gJG1PzChIyKd/kdUTOnGHgyeVw7VuZMhORiaeIWIkitn
H711mrbEtKEyxiqgXCfAgUBeagO/PAK6Ny+eVGG/t1TV6q89hD3vW6Breh+Aa78L
bWFO2X417e8ZgQRhuRw+wNB5KkV7qTLUlOwmLLmcrz5uW5QBIIugY4FaIopd6RdZ
puZdTqNEJl1n2pnIKSqp8cqarb6n26hVtb1Or8P/rFR6aZye1ACcd/eJu//cnkAn
c+Rrm5XGDgZkb0Krs+trjvoGfJwbRw2RmBGvakUBUcVQh+DYZ7x7kupTKyvnTJm5
uixaS7OpVMKKW++PAIflwIPUkoa686MQwcMK5dwYPdDRFcwCsPCoTEbT8PN/Dkyi
Jdf4/C0k+DBOcYhyYj74ctesfUihJDCK3ne7ZwkaHfqgqksG/Dvkw09cHaEp7YGJ
BF5XMTWaJNKJVMxtsImylMl+/PqcN9u9fCt7jx9c4l7y0vF/QJpt5Oo2wXEbkMVr
vJN7Rmz4ZclUQIpsEDuZH5vgW4HsTfSUpej6F5oZJAvRXsDeq2dPtKx0Cpt2CzKy
LzwZOjteC5640dNCZIAtvwMYEATEBW1iNkdItpjuN/wtm1Rz4icXwLaRwhHxV/5q
Oppk/1nStPD05kNRZMqHcFnOeCMbYpHmc2jdfxZKysuxPJpFsaGElMaiqtUpaeng
TwbdkHIPjPNQUya9zouHFv5cEvcUFh+pEidRVidLaj7w1MWv/CiG+povJirmdh9h
RY/QirqYhApT/JU+HvudHDFd1heZd4JLXM26kBxcptfKF9jKETZn1uZM5Rc3U010
Qn2eALr8NVk9x/2OZR0L9Nm7VGi6rd/5PFb37lOOXmEPbpblOvGwf7HGAw2KtPFj
2r6JnEFMQbuET6yxV+6ySbvqr3To5AwSniW1CsLG3IVkscNbtloDFF7fGVRrfFsA
kevoyMVgulnjpSMPn87XO4ArCSiftFf2fio6J+MV1HH81bWAgnh8weMrw2OvHU78
xu2RPIrPYbE1FKcefNdnGgI0d8qq+Iqugm6k2s9HeUQdEfJdD372LHGc7KcMDu8z
taCaGhaMk3ACqGLGxQSHqqgVKdyqU8bY9X4MlpBZf1fzklkM4KHGYFJ+bYAb6xwC
pxNc25HDXwYOjm4cOS4DT/S3AY2BVarFyaBetNekhhmb0A0XHpUda2Xvun1FnvBK
8SEXRGDejcEThfdcUDbHrcylW5qQrztZbWlxQpfmOJ3pZphZWKryASXBa2oJ8vvS
uPooBPrpfAw1d5LrdM8RfL36Ws8WoBzy0OHBVVQWpPXbNYXdZN4v0z0pSdzeWO+K
g1rLYJz6VGtwTLKyMK88Ql5l+iJ9CVHW4YIERhaV1j3n9kTmB3LqWKmQNvHUg5+w
k5eeR/LVScgMb5kAAw7vW64kMC6fO69T+6HT/x+Iwv7OnEPA/9vbb3qE6+FhPJa2
mNFauv5xQYbzsfx3CdVcqRYuniBNbJfvOOg6qG1Kd10C/oeHt8qLBNmaC6DIW1ID
4NRE/RHgcgnHJ2zcYxgrA52ECtmhIhIoPQFVO7Y9WrXMErDy1rjWxpiz9ONDXBri
mIyoIe0kBYi7z4jflAoIKdWxI5rIYrlhuKsFVkQYBBUYEtsvfeyfbLvbIs2NESwK
83ST4NKzAcjrDqtF+zy8esZivwflgEt8RBZq7lxzinakVQXHLbQf1OVRWpJ4NJDz
K8xzTfXKc4polNixsZ46Vvs6T2J/1d21+05fVsX/JJ5LkPTeYGWHcEHgWwB4HChe
J8YX+EbYlirprlimPU3zGEZxo1YRnqtzCEpwINr3VM4vM7n2cro2VHMQzwEiQR/P
ZHPZZEx59JuPz7X4b4HZpL7UhEc9gMiDGo4nYk91sGpFggO25jf8uvevURJx8Hia
4ddAE4uYN9nMa/hRZ51cNS0MaX5oJfwGZPoJyBHwMTg/iIfF9688r4/RyqhZIcbH
L/pfDaSxpn+ImOH5e3DB7cWV+7cK4vds1VohH3NdCPJMbvvTAQG4uqS4LGoCluf3
FpyByVZIGeVoeNcWyb34tSflvfgDWe+SoPZzT+r7CJM9ntnXoWQx4fg83A/6o29G
QbU462IKi9TS2MooLeMYLf48pzqe1MopjzM+UTIUHc6MKRtgwcyOXtm5cElf60MZ
mXYJOPH3me1KPY9NedQsmwUGg/JbbTbQPHOc6yN2lqraYIozfBZ1SfEpbD+ZVJK8
UYl2xabgJ8tQlHpmxjT8IAFAp8Gq6wh/pKdkyhmh+ZlJmsoL91KjsLoErF6pLdxX
vs6z3PgvAV0mBgH/5z5XmOMlatrvpqQ/XEj0jg8hPWvX2aMzuVcuc5PRUOi5I5d8
xgIBByXOhHZB0kSdfTCiLOBTz+fG4TRfmul37DrT8mGWurjXl+JCzYTnd9dpBAhc
u0xuJF+PnrnBPJ81mJfX66ipVeF+QufGjcPm8QXoG6JRIA7D5LH9wVhXrH8hN7Sz
EHcI/aoTntzCeSNms/50xJiBqcEJEcTK/K8z26ArBB4vxsGOOu1kTYM7awZ63rj2
40tfMuxXmRBIaf7oVnlMldu6YypzkVmvlOTuiRBUpQIuvglBJJjbYp9CXYFxqOO3
f3wViB/IQjw2xoHj5HZgvxZBAUgKmUiMnZGsWhXf7zF14nYrgEqdEgAardjySrb3
xrFd7uyvsR7VLaM4laX1dRCyPCYajrMePVreEIS+rIN0KLLg4mGdtP27LkJhCu88
N4CpxG9lqDlurDUQwh79+s5RgGHgCzllLUndSJODU5YCNQZ2WFK/fRSDIuz/+bOA
zMyn2spxi16cR2OBMK31nx2fc1mA91lFpPsiYQdfiflIiljXPMQX70PWfBo93Vyq
9yPoNi5lO9xUpgBUaLkK7FUtsf5WibnXrqFA97ex6JdKnAgCRb5SRMHsCqZcCveb
26lK/ZkXOlRqFOv7KX2YHgtuiGmVVrPLEn91r8hVbqUgcEIo9Urj23Hg7u/6RNAI
JxTCSfT9L1DRR68LyP5mWfDjVSurXtSZFaK1tk8iBR7EwYlCudBYobeWjp8NFL2D
9ZimQ/B5XJYAVxVfEDzxQMBA+xbonAUEin9YAFDZxiL1ovaFqI7If9z73ogJfECI
+t47cKwbATf07C2OHy8Th7ZkpayDfY+tyB3Y8nTROJAWcVh/lKsbdUlK8zOsJKi+
UkyKKR0ypW6xhM5Z0OGhwax2xOHIeNNfT/xIpfFqdqxJ3c/vbLEcQkQAIZs/7kJi
K5JJq/tMS20OiMHgwbh8QsXBuWGFCZBik+LfEGt01K9vA4dSzsh1cxE8ICxAif0G
Yvsu1yu6q+dbj75iWMU1/1QhYcA+NQHdCT8oCGPZ2CkE0NiusO3OLlhLZOjL+t4j
9fQ6RgIn6Zev9LctamiusPP4MBq9d3XixjEhdFxHlSsj4FD+Nanm/lcQPrFciLvA
BExVwRQH5OEEIwYZF3efHYPSev1nNrRGsOJtD1Y5Xhsmsz9S/Azdb07Pn62+CZtm
+xsD01L/BTK5VEuQJVPIHWE3N6LR5PpYY7t3SP+HUvS2z7EQLiO2it5r9BD3ZU6I
7hbyI8lqfSm1x3rY0ndmi6NjfBcOtcE2v0cuScc9anZshnDY7ztYwSWMUza/WyyT
ubRZsQ3gYxqoHcKRnyx0sJAia1eoKBemvX9Z6tbgrmyWjPwR3exOOKppQZfDi5RG
XTZ0SW0FhQ3EpWBohoAAsFXgtvdfhhXQS88jf36fOONc8R4i87+T4jtthvtm6uoX
Yn3sOLzJ6e9Pka07F79Gxhlb7DpB0N78lFr13xo9kpzTmVzy7VDldC0wDcHNhuGB
S89MiSE5jFT9SLjZ74ynGBvYP5Cq1AZOeIqh2G4whdUqFFHItVvRpAxDC3JIZKa7
pre+vIil+1hm3ghuMLNTiZ2mOxV4y6Kl0lpNCxPo5AqrDNMnKy5RaDPAUFbyMt2f
K074OxVocPj1UKHiCi0lJDnwgfE5z2P7vt63ZSx1fTnkmXKp2ZZ32p8ZVSsVo1z8
shCOZ6qezhQlPoJ/SlVmKO6RPeBuNad4AxHxtkPWO7kcow5+aE6uhyOMm67+U9aU
xgUSS5PiVymA6XXJ1VRrDa0rTxYjrruuePZvJEZVHLaNL0rpShMWw5s5odkpf/fl
HPW7Q8GRQvUUxx3Go1aIdIeMcjmhQN5WlHSHBHiqNxYKqeW1iDpBQ08ScX5F/1un
GmqEpjrvyZQqzYoS59d7Ox4hjD6eRcENWY+zAJRSbf/vInN+D6tfmJCC9DOdRboP
e23ozBPnjNtQqJz8rhOULZVV6YTPMK0vWtu8jCZso+eqGa0nlJPk3B0MZbw8/whP
ebSUCttdOlhXp4Jn9AIYFOpeT1ErCE2Nn0QgMtTmLOr69OzP41vLXE+/3+dVH35+
zjV1NrdpyVs9eKK5ki+4mMoc96DWwah3zFTsyp5N/TvA9BsPEKb7RxfxtCuPfdKS
TkB9taRm/97U9emK/RQQ0Q72alDW94zZwi8E7iG70hpGpyAUsLLHVwHaM+w3jqnZ
w2p825rNrdoc0mjLj7VBoCM+JZvjmAy0b4wUgezzjQGfdRQnKhgTON9z/D4KYneJ
G63snZSqO2Zcbc/zEZzmGIrBYHhiOfTxqKj/d72o4U3yqWdEst6fqPiYoOiH6F5s
Rktttal0S1HtQ4V/9EdLX8vYqbAogkjwSRRt4XM4xWyYqsrZC3DcL0qHoJJDVyOh
b8v4PcqL2+zVXlvAoLUrxWv1JClrM62waB4PEGrA+vrjGtzNGEjr7kBa6JvF2R7H
fPbOultGl7078IS2Wa3Go1YTcz6ZmJiQcYPuDbokmr1cJe6NoehBIbxysiXD4C+t
nMdIQ5lmaPvxlKswZR230ZJbSACVUPSkZCHzxEvOR4FVTn9XzoOfRPc/PgI8zHCe
D4TdLQjojM/k0eQ5OCf4YSm7Up8UBA/KWCdSPp/QSX9wKsdweL+q+I+0XG9wn3/V
suVUt/XR56xWS5kDkvORhSPbeqW+1gFNwUXocqnnJ/LjEXGlqoS/G3ubASYy9+zo
LI0Zi73b8C89OX4y63lKwe5k9oU4v9DpYzeUQU/Kmi0QCiaaKHCqQOriO/6SHEkp
Jkls0JCUD1Kj7+kM08xj95bod36D9FQ5PS1ABzFG6d7i6KbfnCK/d5PRPRPnHEB4
Huou2U6u8IuR5hHkXT87KWdf+acQ2i9yxrdXoIf/ODj6MhgwPmI23tmE2RnXz7XK
f4iQZY4JcJasDkFo4b5HyZ+jbQcQUFz4dV3AmAe2kxh4wbAyjuyRBhtBpnGsnDK3
Id2hZPJB+pDSzn9PUeBn+zTzhZD/JRyh/Dy34qDFpmTfPQl8wsX453kWVgHV+DVu
GPWsl4naxdw0HSeHTlWhSAxJXQpGYco61Pu8nahoPi2rZURozLn9ge3W1OtOr6CJ
0HcKezWE4tO/2XUOrk1onbK7TnsHxx03tW4la2ytmnClfhPZJbfx+7lvnh+R6gig
QtHh0ZqnTdnbKHiNoxz0MeUGQEPUUq9h9FmrW8dTAmdSFlDyCL3vExkt0+gyDduG
3j0YBo2ldn2skyEKhTDN+z/JWR1lKdGSVEywisDYNb5EJa+l7FQUIkkLoq5PA5am
SVhs5TP/FiP1O1rP8fa3aIxydq8TQ3tfwuBupforxuvGDBySlnZK3GcZ0+fE/Sll
ypef2QKaDbdMPDCH1uNAOShYqS8ZmviYspC9pNgmfxp+BeB0IkmKNtJcn+TAbRb/
SOwX8xodkWQ8GjE4gxsf5oRESxmFwEiEYKCSJrhZwpxb6NLqkifKz80lpsVicgY0
mJNTGbc6r1JqNRTjCPb08UUpIdEUwSDFur56bl4bBQ3RNaLRi6NumqWtE+ybwkSN
rTlSwUIxRVwDbdxZ8EBQJk+jG4ZBEf2sp1TnPR/z/lCBGE/VHLIHDmkmMBI7hroQ
15kYnWy4QECcV0MhRosgVh7mpktGHrduakZP3BlQPMLMwnXOoixY4sx1CzyoKdpd
Pd/1g0x2JqbSoQHKYRTRsSg7lmcSudVtg4iP692EIhoK9fbo9EAyqmQNmRCQS1Qv
WO1JZOBhVCHRzOrYiTURLcOR2QtUb/9CbADGxIld7JSC9dl+a1MxjgjVHJkqY7f0
fDQLab6fLSBt4DKINm+/K2i4L7p4JvE+x5ehQe+bc0psN15IvzvPili4eLWE2bl8
WlCfrgr4PhuVCR93D6jP595yerodMXYrz3DlUo12rSRr2rFI6vzbLoOXn+38Rm0R
846HclMZFLFqq/qJVbJCdb78ztLuOvazDukXQg0MEaUqorlnggJUWwLpYJsc/bMk
Mlv5xGVJjV23TKDcDRa4R7WZGqqDUaP4aDZ38urEeekvQ9dS/fhmNdamRBtMCxxD
CWG7f6pdkovG5kd5JidFirrjZ4Tgir/k4uMmaLjqRFo85/rPu+R96Rz4gD76GX1C
Vs5MKq1a1MnwwGubhr5lH71qdmakxgXsVvW2+OMYN5/GDObuDUvTzoiJavzg0U7q
UpWce2fnTPfPBbV4T397QPFeZ1cXMSh/Fwi6aMnjCzPStM/zxdlTiwkPKtNIqhk5
3b83UL+D6BiGelEHhO5yQIfUo60Sz1hbY45AfQ9bRgSeC+p+s+P+kDJLDQtCk0zg
9+vzu9LRYOyAH/zJJMBG5eyexyHCtWbjKrjX4mIbBKmelfGyMh76Q5JhN7Ld/rf0
/MZsWwOf2yb3hHZct768OWa29zULFHI4WiJZKF/L/kJr7PnYDSR4F1mea7S+r1ot
54xPd8DTFetm8EM3VULvTegG4LXhjcvf+uWFZFPUTIcgjpgApDqOmqgO8gPLVWqr
KcFFg48Tlgksd7S2rw8RO7yIaax51oKVkQcpMhL4MM3j2fP2Y4uZW0JDPQyaDTPt
0p3ZG+5tFq/qvBzO42xsLf9f1ZfJUhd3GoFp0ltKTeaOmP2zryK8r+CGMZAccEid
33JGD0z6nJ9VWm2QW3j1FPeUK1LwIVtWG9xhiIA4H7BqBnNJvyS9fLrRfXbLnZI/
gFrDRfKCmFaqLsXi202nXsQPE9nbDl2r1JGSo4Tof24MGSS8ZtwbceAbUtt0YCpU
308dd2lNo752jj4HN6AEvUVlX37HJLfxynN1fFESoFXnLYilYhEfFHQjRj+6NWW6
UvolmKhZO45yQk9a8nJpvhUAWbJD0deJxv8Ta73jOuNVD+h/U+MRR0V+bQvO4K/4
BpBT3ZFIvfraDd1OgHDX8kE4dATeYp/sqPzq0QR3lnNbNreGC/apAUdYrM5fz2QG
N9JAeog7a5sjk006xacpS89scQq3PO4TBBXEjV/8pqZ8HPiCqKZL2tIVHjA1HqQv
4toxEM+1mLrXW70wUWkTaI78I7iNEVF8HCsLmtUWoZ/2U4zXL+4/uYHOTafz0oK/
hICCKjvKa97ucPxNU68w1SCgrzWCVpAEkSIjf/vbnZOu9MDcd5TKRdSniwezLUN6
qnGpE3iGUvt/ebMpiUEjssYlPHSwrS/fv7aRCL1Lnhp6SOKRi3V4jG4tpD1cSVk8
4u+g9CqId6niwvX7kafgWQxGqCj6Fx9CyXrKmpV4Gd0xw4N4lkRY0qDu4zwWy1Uc
4J/hOFjd9z01xUqOuXjxt12EWuWwhYGz3pxkXI15ObrjrNwjCJi7SABPXOlXhL4q
TrGdlMF2KxopdZFm4t7M/ZM8xih0mUcJUn7wEG/APauVBprJf2fWw0eW3SaEGtdp
EaH6oTKnlgJcwvHWI0dckuUiKlegD3IqzI+laQ22uSFoVBwprRo7a4Jw45moUPcO
r+Ve+nwxVwTsO5LUE8X5ibuEzC/7jui5Fm8rHqZ+31cF4/bfPs5SjC56dvdYiqse
uisBhuXxrzc9jTV8oN3vkhKGattpgZ15YLALNDOCsDjfjroZrxGcamN7T++2UuIN
NfEvWg/4W05WizeRveKhGEOYUi3I7XmPI8c/53GoB6jXvSFG0qYA+USWHoMKaizx
inz3Kt8HALue4tXvOvD614HWQh9GGoljKHAuRgenuT0UCvzUgC01k4gw37THT/H2
8mv7p33mEgp4i2O9GYovt0y5jAb5pwybI7xwtPtGwFEVZTDmToxKt77H4C1cZjFe
YudVY5JNTWfh7C3QZ03lx4xYEGLMWNqCKmvn+Jklz8Cf3SJFgMClrV/bAdGi9jyJ
DW5GGdsQ1J7SUZ7D8gs5/rnv7QazI/h5tVZANNv314JJiRNVwcvBd3jnXqHMLpF7
oiJ4gdVqAp+q8qHf9AzLjhj/zwr70/Cc/hv3XmDp484nS8aM9PisKMlhnC13hP1M
VE482XzuyyZgmC/TqFnsBjDXhgLViT6Nr9hba36cRfMkJNnuxz0VAsQrc41dv9L/
kcjUlWaRc9x4sQ9uztLetzeZVmUrxb0c5t3O7XET/i2LezM/cO+LZEYxhJ6Oc69D
1COVaPrd/pQ/Ve4YoPXpwlpu11rWy7mTZ4mhQzjgitARMsZ2WDr0uNsowbE2I1YY
SqP3phbricqQPWBu+uazQvtncpxFSHGG4rT+sj6iMN2KoTF/fNSfhKGrixA6mPl+
49cWMJrcZwiZX5t0/LT75JoCdx1REwHafz1Kq8GDgybuL9ZlqzKKfTmCSjPW5dNZ
S/VRePg02xoPPAm9uhK/F7Hi85miyn4F4M5VU9xN+IQpURHeoLB/FL+XtWwZtd7X
i0nrD9PL+VGH8NiFbHcJN3CFjMAEvVKYS96Kfg193zAk/oeFHsqyLItZG2cdnLQ7
l+IpEvrrRyPOq9f8oHFGt68zOfGShVx+yMuFLBdVhbNtiBIoMlhTRdGZUSZqGWGv
H772oSFKmFLtTuJt9fCRyg/NNPoUYhiv9kbVQ+PF3xzm4t35O1wB1RtjnF1tTiLr
w/5F1ANlOc6w3BTcJBjyMMzrVKe/ENRynzCuXFhEBmeUEzG+xTOW/BGS85rIL6x5
abclZ35+rS2ZCm/2qu/tirDgA9NlsNyr8e3FdPAGIc2wkTG4oPlJ21JBJODuLHmf
yeuNIpZdOiQUIjrYHsCrQWbb2cOKYhjPStuQD6tEJyN9hnj5B77/ZPIcoOSN82bG
GQMUQ0bSehHxm+cC/FuVFfuku/4XT2DVEQdWenlmWDUCVuZMaF7m+N8aBUpHr4QQ
ssfhj6avteEYm9gmsAUy6lXMgtMzhcBW+DsYtPF0xzdB+ecYFl/RD0Ov5bH4eQfI
nJlrgykysH2mqPKyFy+9OhpY7NYhJlKbmue75hNB6XV7j2RQScDggESF4XmoLXQv
adn8YXGx3QyVZy5spzq7BbHdtlvthTKpZ0lNwZpl26zmssJ4OAodDzZjWTj95qHd
1DFV+gjQ4gYgEGMdJnxRpRXwWqE2EtWCD4g7YAA+1iNCHL1SR8ynVWYcOBcbRkJS
2T32xY9hkdyZ2nMPpWqHk/A7iS02pd0QCxGXb2OpQOSC9iFvZhf2O53QQrBW0RFG
09DJWLVjyHcDvkBNgIMngo7xib8/C5vGg9V8PXfEmYdDRF6s3Vu6ExG0dG8vOCFc
CDQirZUMXE/I14CXxEVALN96d/ajkpBcii3j0RAv67aMkwnRCW1ft7Rg7XLL1JHZ
aoRpARFUQUKNYVwTIsEXf7YbLCPKqVVPRZO9cqRMdRw/pp6Inly59DqChECx8BqR
FWfL6NpuRkqP4hc5/oXftySWbGmU+9O6HGtltU8vSe2PYzG+lr3jVyYAv6hCVdFS
oI7pQM/xOIUgs06qIs/XbUuN5I2T2I/o0q9cI88g5jdjWZRb2kZK0fE8xsEciFCI
bHoIIGCJp9aD3WBnJF8savx3kuX5Lghn3ekxMlbulZwFfEGLMLZOqodbQZdBkUr3
04LAJU7ADMdV7z1Ki7DavQCyRtJNpt7DgqU8DiD/STUJ+VSjazpgLBv55aLx7fBt
u0qS/1VX71CTMlkM9gO3hBBpIelPN9u9ZkjXf2s+Rjx7h8rVbNUmUfupF44WMpxe
yCEYyslmKs17iTND9RwF2qnyzZlF5d6RnE9jsAM6vUO8de/TWd89f3IoQKJXcwem
hp3my0r62xOhucjtAjJ8Tdep+C16vIcG/lcTo0auvdkWs0NezXYGbAQpPfe9QJuy
NWztMuIX/4voQIIfrzLFDlFwRxxzB7AHm8IvTy/yWgRjiY2J9PpLhqAIUNTdsZ5E
PhH+xE9S8UHLXDAfZJPW93l6otLGSmbTyaozGlEUShzQjQ2tm9sOHjh1ARYq3YAw
qNbP0JL/PXmSpee+viKhE1+sNY8A5fPSwFbjim83EiNGFvKyDDfOUILz8HV5qeMt
Omv8wzBs3h8acnT1apAemsHVVPOVzYK2vzCOoDXCT1yMUznplmWEhj27VHl/frtW
SvYXtFD5VC70vHJ1Y2HUQx28B7HAGSdleTJyytcDZTicdKxumRUhux5bs8XXaiGa
mLQILlTcwhvSYkx7IhzMgOTpdQrWtIoD28W/2EvXDJrKm5KcgCDlMDYXCrZcJU7/
pdExCBkwnE8kcxAsrvK/sGki+zRmSJXKbFLmKq1Dq5rDHtjXhX0wdC30oJxJLVV9
jc4zUpIabSUbbinzjmwLFQJ3MS/Sv2JSUHIpj/qyazOWnGuVx1UAOsN/yqPIN+6h
a90ID1WHIRYbRx58EZIIrjOHfgyVEdDsKVI4hVBEFn4rBBE6VImf2J0Nj313NXiU
Y1g4Ft/9tJEAikPIVUqeOlyKHjlemTBJH6HhmSluOH4o4PlhcdFi06aGCogNvEQ4
A9HxwqQwwhiEzj9xcWJqnVsB4UpZTIVLNqQ/dr3Li7WuxBb2AJ3IXe/3gFqr21jp
4tmpmb3XqoKk4YXjPx5sv2CDX9EAEl6PWSCX9Cw/o66U10hPWDVSEHQMD8dMJM00
a79qF432SN51L4XaS6o3W+OdmCWXRddEJonUTy7kZJA2qm/ULSma5sk/fWCpq7HI
uwj2EujCoAMYypxFoDM8pbD5XPuFk8aw7nArknEdIT/CBliRE/A4oOm08qJWUJpE
AWrNS3hqC5iIfFDOBXEgs/n5ja2V8XIVGSQOW0m+1FHq7VJ0S2Tty0fcE21NDUNa
l2qJTDsDG568Kbf5oH36fDi567BAfkwOjRfV/hI5h+J0S/895BO0xNp5RgwhDPBB
jmlK8o9+VTatrQHphlR9FvC7QOkQqgGspQFdo9/OrCtr+AMR/nnPXL1dU8qjBuzN
wFeVi/SlXxbwkZZn/a+Ud1LDWXhA5/bJogWxMAGQbbsONT8V5wN4OQMPcJqLfHaa
n/cs9OemGHN046HSLxANitkNauSawcWkvqM4xCk8C114bM4eevWrZf7qsiowFmO6
h5xSGW3nBfA56x3gZb+vQv5I0Td/JApRuoaoCTXGDNnXeYZBXsW6/zVUxYxW3hQe
HaHzeqzogXwaNxJf8IsVdKzNmAaxkOUAOL5tBKXLD1Sb3q+CByjsifewtXX2EIb/
K00eQIHXsB+5oQdY4lnpM94MJxKSkj/kph8bnuIhX2NnNIsp1ShwgjW6TfC6hQ42
uhzlllnNqsrluWSTY3HHHr5qvgN29HioBq6S5YRwT6Wp8OOYDyV1Ai7YmUdkwrU+
U/T5BA/rxq0sR1ZzarH6tWgnNNBdg+ONjZuzOmNbB75vAgWUYozk7zkoMn+rmpgh
fZRNayxqBO/+voimS5UV5l41t7rBGVixDG7eEAeI9g7QSyOfJeU8VocgMyQ/6nTf
2CSUc/HttJWfEx2TionhKo61YkSe+mYbHgf1xR6hkiX/KQgmiJY60jAwzBB5Ktml
FE8nFOqkmC39GxJgxLWm889rPy+RnABkWg//H1xj7X2ISDBaEUea9eKLUfo4cfh1
lvAGnLaytWRPC4BGO4Ud5dYTWRxD39xya8bxgcgdVuqc4DqZPNDQ6biQbMH7Il9s
vaGeC9uF1nb9DjaRw/KiUMyzmu5KzH0/5KFL+pZZK3Sn1OQMj6PZ/kWZ8pcelxZ+
pkU4ac9LZy4GlsIFUGOfswWfgS93/CDqcg8hGP5J4d6hdqeZ1Ps8ppkKeqtTXvaj
gHdTARbrem894ClN78l0FRvErXm/wNxrmt8GFxLI/S4M/qHDpaSi7HCBeXJDMgkU
FvvI2uFQCVBmV84mOSzYmRv799aPngRH1MgqRixyACBs8aUwenwepfDFS0zLTKvl
xZObBue6tqPs1gN+OnGBmqyMmEhZd4922Q+K5dc5g9W+hpEP4jlI4WeOpCtNPs4W
ad2RzvzXz1vk+FozG1YHOmLSktuc53+5FcfZhBtrfV1BaCVXQTHXFT57ITpRsvkM
1GvCttUF/DIkfEe6717826MPVPeRRutptiMHteC+eOqD8YIM052xss3b5GYTcJRB
YcWsWbCLzkHqO0sbJaOSITrRcGhcQ6V/9JloEYbM3m5O3kJBahFrQ8Fd0B38TLWL
YHFa/zLh1pWHqXqmM6Xqt/ujPiaEg0DLEwt8Qdr3nifOYIjYUqJjA/AIxqRgyxhv
APPNUdBoj6c+wXNPVgcbTC0Th0NgS9HuRIjXo9FQDZOMA5xPRHSgosPjUMNf/TBA
o3BXrkSAqqxu+qsaSoC//fxS4BN3hVKKt2cZWBjGujSC5F2A39XuzPcaP7S5yFXd
0WP3aQHmLKWZ7/nyX7PlToTSqJjlCcmviZ+5jSYgVN2b5SlGXgAmUiWUJuiBGczW
lBVLjttBIi/baYAMX3qAXVFQ1uQc/8TnDiyPDKjJI5R5d1RC3DPUduKQeZLOfedu
O871BbEzMWmLPXaezL9pkIpEzZYkQdotxjEtRFc46jppNFjdIQ9DviStCdtaO27+
0wYr8Zb343sXWEBdILWdwHTs9x3zHmjAWl0BnLUNxXxlR3wyn5EOCts1JInHdKp6
R6wmHKFLLUyI+P1E56OA9spGKSUUWZMjvD8JQLrSbPjFVpQ3JFKefK6Snu2XPvVW
gyIW10C+7uRSOGGTxwdRynoAv6Xd5Fo9pWjXLDaY08rQuEVnwROBkFJ5dvsjsFvZ
jgLmLu7XAW4yGZ+iNbcz9BdK5RbpYMn08SAUQcV0URlB5Agnsg3EI5DDQYJVh3rM
5VBUnuSUtpQBC1GfjSMZYMnLbNbykw4xwDz61xRoxX3wdNyfWEAHpto8J7yFGX1M
RjJOgDfITnuLNJLdR9OdjWyx+zeXlfa79EQ8I8G3dAXbTTtkBJyGDy3poZ2zNN7p
SajQ392mgZ9U+ULnWKsmzgdvq6VZxfGulYJvNAPPV0csdS3JhK2D/8GirAy+uEq3
OFTklZzEpNizimpJvrCDXCFIlnYD2i228HePl7zS+eBUfme21rVo6clnlklU7SXT
LjOyU2JW9AtOwwNexgq2f5tOWZdyTVyUPFpyZiIOl0PZrBsZKlv7kh4Dqj1eBgw8
xIhsqlqIZCmGJkaxWVWCpTbBg9ziocZcrNiEicZdoxOyljW308L3N4qi9NguMW6E
45R7GILFxRrfc0UItE4NIX++WywnufPJDE2oAQUEaiZTLPqQngKJfpkeYx8xgP9j
90PpJfl9arH5RiaL8Jkj9jTQIkcBL4M6VwEQYMv+XRkfC3oBNcbNroazacBUaLsY
SGEcgykPXw/1PJSaiO11sCEwkg07nOsdRR5MehZJy7PwndFTMIaHEyphduFz9Mp+
HXBpXR3l+EGZhXPtFv2SjBugnW94wRGvxFrbVpI8dbKqHXSV/W0FcWmnqSL5UFN1
Yxg1h9MEUryBKVOrHVoddA8Ic5cCzZl/45PSmksJ/PZ6WbbFA36yhv7Kh6AONxak
IVGa50uAbbmFwF7aiD/9Mxc40JQX7Z8bcgUXH26DgJDN1cLrS5bSbA7lDHj/At5d
r0WbP3CdTcs+Bpk0u5Ypax3CzIO9c4UDFtLnLeHmAOdrAwa1IlmbmMQXedeoo8u/
uQ2Rp3R1ISVmRxj86rTkI5JZZeQFNWVzMRMUVSjJSViuOzOi/BQ7Cp+SbdRYpckn
CaR9rWjf0tC1D94NHRH5IMCP2UycVUdOiOeJVVTwvihc14UbMLSbk7QblJXkS2UQ
eqd4EROLzWEBWpQr5/22ynDk8m+CLYeav1Dl6Tugvs3FoPN5Dwf8xI2nzVxYY/1q
cqSCgony773VpMtuzpPiqDU9tWkc5W9FcVxctasm5a1js4Go6k2rIAzgONAJff/K
OIy575VgL8/iQgoKDOYFxAnd6wG6EFAttuXJu16KzR4GYeEHd3dXm6ZpV4YG3XCy
xQcpOV10ZilqFBfgJieEslbb8sfpgAz9n5Vh5bcfI0rVs0KJkpaA6o7PqSyzcthn
Whcuynw+3GRuphwR9Y7oz5zRuNJCSLVTdMZebljdcU5AqyDnHXZBRzZ/Tn9klXRs
BLmTT/w1zRi7rz5oqLlBgPPaSAtrz8tRV/gZiwBmGS7DEZHQzUxHm5wANEN6PZfK
l9tQ6QdakNH2Lxqo5BJC5b+2b0SYVtTPK4PPPiOWU/tQ5ZNuJ301/2BWrCxBtCsi
333fOIA0+FX060FocT6MnIJ/f/t0VI05Yh8UzGI8TlC7jm1E7V5pAwozXLZGNmNH
0fHePTuTareWedCyT9xnNvHCZOZhibeCo4DkMmXY3H346yBvTon2Sq2a6v3smv+L
q9wPhe+D9oWM94Ai8pu6YqbsLZkK+5Oyvw/zasKpHTtGlUnhljg3W13UFy1RqN5J
b6bU2l229Pthh49ameI+icU0SiM9pXkHPwZfHcF3hKua8y7Xmhspy7V/gh5WfNTA
yaHyMQIxTHF/37kklZAbLr8bWtQ+8w+f1C9iApEspkT1wsm6phPbjxzL289FNkZd
HXz5Vpqm2fb4eb2BVFOmvhSXYfulBKHIyRkXQeoR7AZQ9jbiUAtrbTsUNfiF6mxo
k/0vaHJAFDC7jb+c5j1EBniwIK9Uk77yNdu8XJhwODOlNFEh8cugWuTvXRvywbDC
yq6GspKfl/dMrA0vh6D/YeTykzt3+FUerDEhTAluJPPQ+29RuEzzU/OkY3KEAq8E
jMzCelOgbNAHeHRC1YZcjm5fRjh/WW36mWMU3Vho6+C82Er76uinTixExl8Qj70R
qa0XRDiff2u9iCuKQcc4YgT4scrEzEr/AghcP5I3hnIjCOHNHVgbuF5UFrxkgmdD
/N4M63BTSQjmGpjxh1Xb57c0HDyWbVCuplPVDeXSSxU+sRKQTlTicwwNNouNMuYZ
YK7wmkBJlHoOdsrX54+8SkEceXyNJz12p//GGMk7mHo4bQ3Wc+TvlnC22zf91r7S
0CpUSY7KgKctS6z61+C08fQrQ+r9mJcHzFvo+27KaU/ulOd0gtVrRT89yEEtyHZv
T1/wIf1RwxofTUlzsmkT1sO3eOol1wNJzy93wYdCJDRtkR0aOrZJBpOT5Hj7EpkL
O87DY/oJcA3djPevTgP6Qd5TF5/FYD3A6tHJHmLXChV/uq3qG5VYejyGze3MwO3E
P9qlUH7tFhmXihsqJwAHuCpvmfNqOxCupUhWST9JjfeDbiuJV9ina10ptjExpvpn
YW2cs9SVtwVaqBFOskIsSCJMJ3z7Aq8XMUOI1eZNf7DMd4bHHqutmnU9osvS2SVU
9DZl2G1TG59AI6e5HPVpZboiuzBfI0wq3OxTI+82+VLrWx5TLnNCQKSYhGO/FF0w
V/iiStwRRHBzWDajCVM6d5YgjCMVrGJAtdqet0UNyzF4pVDNYZTAcyJ9qxlC7l4x
ag6BJXwptYABN9s2mJdfGJCZ6qrngxgG3N38Ey8UbGh0/S/+iNCJPlWfFBJDruWj
QFfmvzaZip2ohECDBjRjb437f+uxLnWmWJDuy+XQMJBAR0T1d8Q628zd8wuMCBIu
I4aAxfgaKG4m6y8jY4Jpdnvo7MyhFnurAdFjowLXCe79VfHTwlBgDuo/AF1iQoYo
FWzFfyllKhEBChm12LC5AE4P5XRon1cj8yZ7Rz6+ipeV7Gzz/31aJfVxl5FQ/fnS
3wlyemMLDrfNWBW/pzIdxyeu4zr5b+t3ksn1q/WsmyWuQeYpBAJ44Qx7IxG4Iw5r
bRRNjtt46MZARt1MT5n0VWs9fZuOHw02VKU052lDS08D09QrDgsDuyRMEFbeleh5
bZBJg98h7fuBBCIUBlyOQOi9mKDfHHBWRLXX2Ss0vpOf8FAA/O/xm/SoDwq4Y7YE
fxVTBP6A+Y9dENBCTSoyeRjXqxfKFgUh3+/JYcXeVpBRpVEIy7MQ2svoYXVg6B45
t4renDz0aFfRvx3ShCa/HEySE+9qXJ6VGvQTVpGFxv/q8ZqVH9LAGVSKKvxl1irL
Fu5h1sssc5QWa2wdziMpziu3duLPw2QPyf1lW5SAhxc7ZQb/pSALSzkPsixHZwSi
9kg76dB7N9h9NAk53FG8wUHdnfjGqAAbPLzxE7EdnRRdsd5IK3CzzrAxnEtATXSo
tm3X4rGTiT4Nm6u0gnr+EI6Qj2zLSC8IDDZkNYdwzd7aKDqqkhSr8ZyDDyNz4Q4+
UF0fl/cfGkRnIG+5JIIp59JJgEZKpm3Jalslich1TIF50kMsJ+FWVMjDhTZh5NfH
oZjE6JP9gaoLkFU9leWwkW6jjvJC0wU/C8eE0gB1UhQXlrDSP+591TgipjgiIj5Y
qvuzeApgu9d7dn0SEUMoS4aNu1zZ8TuqUKXriMcr8BbQpKIX6Zq4BKm2IdujIMza
AZAEYNQCf05+vIJymvpU2mw6zaa27ftYrkvwh9Ip2RWD1gNKxpfUAuku/lGTDgrW
FcXNuT0kPqWHclV2w/ezFlHGPxOt6IZ0ljHQumtcaSYTa3VA23KuLMBgctVBUuwP
q4BD2iUdpsktW86hSoAxPnFeuVURfkhL0nLMWwRDNrQ1XXf9wl2QFQhRseTnAdz+
kgzRPjS6VUu5zX8h1J8dDgWMueX/1I7XxyjL8pj9Pw/A50nSAPacqO23v0eqNKEa
tWHWrdHAEehOcRa+xlr3aOj6p3RdHj2HSmb2FiNzypNnX+PYbJHFNahlNRYnkieQ
u4zbTtl3k3eTu9SvjTrCz8bLDi+2u4ZRH4ohvCQgVs5ACxapCnnVI59Cr+QgE16F
Y5704nisV9lYSr4JIy/bTHGmc7fNc9WZ3FDZk2EHYsE03AAX7ZPDuBvkMny1Oar0
YUCHeuK5GMAXuKbbmx2cmo3dyYIQ7qqfDceUOmxpBbTwKBm3ddgaGZbkjT0wk4V0
wtZDAKwmZuInNxKMEmXAfpvB7Dg2eLV17nSOR1OXyOCOx1tuUSutXFMfhZNGOONz
SuZx78z+NBh6WPEgJ6MfX2pXCwoWp+SrVZnMp5CoNCM7a7CY1jxrzhArwXUU13jN
L1xB7M7LyWr3X3V5OlBZ1fM4oFZYWOWHmX71QXdA+GoMzJEkwKWhaKaO4NAirWxK
UZr281T5ktuCog/WCyuPoyZyV0Gsrb0MZF+jYuHwPPPw6KFXaUoORzWWcNgGsleA
jWzvss5+EDTLnVX1ii32Ts26de42GN9Dyt23vxQWHgs/aBopzSzY1bq4YOkk68Kg
h8iC4VJV6+zOvZus6Qa4dGR5O5jE0SPjAoAUIraKpD5cxp/8E1iq9oR27apCh57X
gtJNSNe4SuGndKwllwFek7UnpALFASx3InSRjuvLRIvNZEG95xF1ICrXhEBXX+Vd
/CLTn4Xg20SunuGx4J2GD17Ud82toRk36gtO5qU5ujROz3t2CSG7zn4kCnmy+eU+
vvtfijCL/Fd3UDdYRuhtFHPJpoux33gDEbECLJsZB2bzPgcHS0uf3L7TQqxbIEqd
a/aTlaT5MYpIHDCcZH4O8l6EXYnP6L/n1dbvITxhfBplMXucudWrHz4DSxhYURm0
N4WTZrGjemawqiupU4GBAkVSzRthSVsw+oT8z/YdZSY2y+vgQzTcteCsAGHCElrr
O4k4KomAnDBjMhHiwtwrGpbHJjJwU/5g6fRsQqsnGZliPSronO1EwaGCwRQAeahw
uIfWNCMYQY/zVvrl71GzTsP2bnygA9g+ZDlVTVeWsl4yRGNH6Qp1Z1j+wE8ABYOR
7eJcs1fnoC+dHptVej8Zl0NFaNuoVVYah/TR8p2ecHJvjkyDKisxdBRvaIg41v8B
ZO0VJzl3FR60aIFi/8AMw7lYsxNBFG+6VlgLB/LtlMg4GZrm2pjsKtwlOL/YU2t5
SNfFxTNRZhgtTeV3soLLbKbFQftvZi5XO2w3xI/CLN2EjXVbfeE+eB9c1rc5dwMh
E1KqBjVWTHTTNXHPYkjmKz0sGNuBJE2m4mZjK+lkV2XQB0ukmw7Mdpvx1+MeSyvC
GDGJEdcTIR5g87uVvYz4RULaaO3WgU37YUrhUFWkG42QRgWUxYDdmAg9vyTyams6
tDkKu7qmuHcqv8GTSLNkZpddSiHX17WneMr/B1w2ZK40LBZbRPEcWcm0lWJbjxeI
h3QWndeXhehh9ZxH2d8ME4ylYL8g1BjZwJrI4X3qrMs4MIBWZQWd4B4SFRnF71Xy
4LsuTJGMrirO645jyG8pnM/ebWbDecaEep6O0lD97Fc+7FqT5Ss1ADr5FTRgTq66
D7U+Ov30fqGDEFoBoWi1USrDNjz46fJUucSHQSVij0gEyqgmBPm0JvKRdw400PMj
Oe1fcbdB9480A5n/5DPOhdw1hQeoZbJlFlv5XtW+7NhPPEfJvNGbltsxK5S+Zt7Y
G8IxKM7exVp7psI0SkpUfddbn72AKM7O3Rtkv7J9ToTMD/71ELx+GGWHS3xEefei
E0YNlDxZgkMd6c8IdMncUQd2IvjW8NSP9NgMWqJ1y2eeIsd3k/jS8X8KhdY3nMaF
N4IK4Jr0WImLzvcUj8IKyNL0vwPu5kQyBhq1C2ClfbFTaow1eAkkpN0ozXcgU3f1
VJLpiPlV0Y09MrUEC9yTonPMT9FmWmOaf+6nj/3m0VZ+GQi2wLMUq9nSzQ0eBOHY
9AAD8ygIx2QdiFmBPBW8OdowUQ150nmxys1t9WW6F5g7OtosNlgiqwpRXkPaO0mt
/2I/4YrMk0vNwOiX+qWg2h0EiOfeAdCQ9TAS+yjDv6XjmJsUz+SaPYzq7lfMUsJl
2uHRIYRH0dTCDe+wONNXXUKuQwtBPvE0p/eB47OscaZZMazV/dqVOWPPsAB66KS8
ZN4xweV5oSLrkGKhoAwE3Vt0flLbRGII4q+4KspjPQs7u3MVadGzv2b3LNXzj3IH
yJIeruKKN51ayAo61AQy559ergK7Jtt41/miFw27pSNDejoYFQ+Tfklv0sdq00wR
AqBvhotXViYWf2z5vuX3rsP63JVDqdQKIUhwcR8SGoq6AsP1rh/f7YR26LmpFlMc
kjaadKY/ovtCPaLUtY2Hb37HQNNqYFQZKg8snQoBTtxuscfe41bzrUbSgjKKxCiz
Y808uvf29DBoqk8ROnXmOj1i9T2SbIlUX01G2Fkox/Yk+5tY5WvoP0UVr455btBr
ePMH+6I1PtPHAe+BM7u6CFlNM72+m1nNk/TgXV1rlXL+MWn/Ybowwxc2e+bQLTMO
IrzmK42vNanJ4MyqHraDLMFRMo60XfRQQfB1qO0Y23dvQ1VbDTDEj1xqHXVRndpg
J3pNMs+o/BzdxTeTm+WAc4Jau5el4kwOXG91Ov2Epb1lL49ao+f7tjAT3QtFSPXd
xBRlgQRtz8x0HghrR5FU1k5DHX+Z1ks7DWANoMShYjw8a5sbnCoab8GIckAhneJH
0aifjy7eYHKPSU+LjnhYV6feWryukUboCJW/WiclhdoqUAlmN/iuBIitJYqOAU24
1mOfTARdgVfhRxcVBSmZ/OY142t4IH/RWaRqRysKT8l8nmuDlUesaYUvdTwwqKhJ
7gWqXP+wbHEXSOfWa9nBX4MnQoQw7kCdA+JZjSW+ygAp5riR10XMIc/oqVVeS2x5
2abkM/yXy8TxIA+WxXy69ofMet2+itVfp8i/TGc3T5R8s5Xcl6AjsqbWfboQ884E
5wVjtxxqoTImjrMVORuqWSerYWdeBS1au9hBU1Wwa8y40Uf8lt+isD5Mh33TNF7W
dV/Op/FxJ1mkm6/ACncl28bpKZDW0xj1YQqL/1BwjW1v7Hy0NrHZBvVXdVxheHvg
UIrA3x7CyQ5wKOW9UphGU/GFx95AMRyeWhVJw7bs1YPp1qX67nM8DDP8c/Pie6Lk
1GjdaI8JMR88GYSxpxOb0wuSXdE/+dMTUYjw3mfzXgB63qrCXrhMV6jgxsGwCAfL
9/2PCaT3/hXQ64IJE7+MlUUTrHuKS4fyajzJ7m1bMh0JY52rl/2qnWjfQNbb/ZSy
tHaq1Ha2FQwBAf4N8TXJWtgCoIp6VOkvNe6avA8Y0u624xFSQWT33jdtJjJWzUs/
FzAsgWuhM/J4ZHTMs6x88zR1dmlVx8xLeIIvb5sfOsiytRixXi7wQM4O3XG5b7F2
0KPx649kndzJZxagHc/25M0hvhSZ8s5miwu7Ic0lF5E9NGJFHwgAEDoKN14oq3pI
xW/5QrYv1332vdK2aSVspmRnbrhZvjTxSo/c3akT/hjbMRHUH5yHO9HlMY2vvW06
3twZx0TllGUqzCSHD7jhh3VJToc0tcdDCqm6BrfZzI/TEyFxINkD0YgqkjExutp8
ogGqIOqca4Z4j2kH4x9BS8TDoHa9p0BUXbBk9uPWFCpYgquFK3VOEOmNlKIaIDIg
48vFnGT/Rny4l1qQe3qCbIllhqlIDx4eNyPxcCDgEYPPXkP8r5t0SCEEXcngTPRp
vMEv8eNbPov1czJ93eTDBD5nQ5vOJ0dWvbdZOEsqNBav6sYBgXj7EAu3VlT/HTYQ
yoeObCZnAgIngKDvPPD2vmvw5/OvGlQ8sh2g2k2f3LfuSmwnoEoSeOeE1x+IKlKi
PFI3U712WZpeaiH6uhKOYlJ3mi7Vj+9hvPD+qyqKMqVa4DOlwmHR3sKUeX0uMtM+
jdWUYVhUOWwBv4LG9UgyAHuwmv+19zHt+HhyMUJ+bHf1a14Brt9L90vl4wQLtHih
QjILixEb8g6NBWdCgAekPTcuJe6GrbjB318tOUuHX8mgb65Biah0Eks3B7N2extB
4yL2fWCGzN8T+0cJWfiLdIVsmcJ/kIF25Vt86vfzoKwbustTYnMnOhcRn7KByZ3U
TxZYx0nbllLmb93VzGS+SphfVJYmjOZWIwZbiwvdUovd2ECBnVkITiIy/GQ4LqNx
EvJA+a7oYggf+n1QfclpQJaS1vYy2T95wtSXvokf75pFUOvdoQ624SMWrgvhG3QS
zEMHw+GWJm8x7F+/AgtN04FnDI8NgV9ZYZZNnDxKhGDjxu2z4Gxx5JLw3Xi1o+Uz
z0Se/Aj8mb1x72XeF3j1QqEq8Bv/hAWl90trpHwcS1eV0DInLpkbGzKtp02XZcnF
Fpo+bMx8tHl6JO8HQGTubl6Ix1EtVgu0w5pyTijkhqGP5aXthzQIRrUpoeQOX3nA
0Pi7kproYBYBIXeQosF6neO8DGIe7RoFlscbAoU+xlN+nTuCqpDLlc0daiyr4BBF
lAt1vQQhnWzKiT6NDAtmLDLvZ30g2NjiS9NKH4ajm4pg0xG/D2gZUhX1g5D907Ow
tlnQaA+n3NzR/gNggn5WB1lI3DiUT9bZt6PeoXBYzNXdN9cCdXd2St7LjXUMaKm2
WfaysWeufQ7kou+jRtXROiPQfXypoUOGYChlfHiab32x0Y8uqR/8g7wOAQORe2wg
39VN0j6w8/JRct5qYcOGWDOcSBylrlQIcdvzWMLL5HFbNE8koKTFm4cPVdLuNPGM
Di7E/jSenZFSp2jwG6es3hz3dsZTic/DvOW8VI6te1aLk453laftXz1C4aHnpw2J
M3cxq6Iga52FTKLowepnFqLDIV6Mj1PPAYdA33cllxWyOBfIo2Qe8LxrWNVnYSQ4
g5j8NmoIf0uPaZ68AIDh2dw1XmtTO5X3tGs4qU3zZ1zbnP3rE8Awqtegq5dOHHNg
VGN7EVpXXCQoW4T5SktYvZ3fJELEosqX8scchL7ZaU1pUyUNVKGssqRw1O9kCW0g
L6VUpxtstuRmJSFZh+/L20/fdYQl4wYRbfP5Dqr3ZbwmRt1X1e/gWF04mVUdXpHk
/807sSM/ilAZscvzCi5pR7UoGJ8EfdDIfyC+AaDdO8gcao0X24Z1G7ydq+6xnpYe
Rky/dA8Qp43vV1qQGVRiMaK8ZmilwpS7szRCckx+IalNfPVcn4++OMibQ3J7Thyx
z5TGVprTKelg+XAPiUv1KdKx4aiRaCS89nlQeDCYanNncn1vQppwXAnvktzNcrz+
qLba8wFHGW4aFHS7vdsrGFDjYF9bK4qPSNZfzPDYU6ii/OM77wKOdKTL/wxh/Mzv
Gk/QzOkB68IWhFG0PiJbcTZxJolh74TriYwkTuDeYYQqGOX12d3D6TkFj2/Bb1Cj
gQlzWhiikuw9fTcoiSgAQHBtCCzWThZy9/oDiBz0t54cwL7YH8f4TMMNoxalQZ46
omZduvKptsAkLCimw7dweaXu7uaEvyM/hMsZoBn2gbI7KWA8/VRZv09rp/F5+pkj
TLAM7+ZsmOARpQQZ10HKtXNM80NCiJk1zlAhA1PZSZsXc5/7crGmnEYVIr3WLACH
2AtvByin6KN5u/9GETYv2p1UcJQ9Njs48WW8k6LRj2SlzPRial0gXeYL52MgCBv6
mxZGr1lwhWTIkNFvoFPkbzrxUzay/+HqazmaWhP+KyV2U+ENCpY4+ZXA9OdDQfGu
2ceI7xH8F/7SMFcIULnGAMW4UBZP8k+raAU35najINcnfv0vsaO6zyHGyZCOGaHI
00i0mMsbCjhgAtL/17dGMeaeSWqBgcxEbVg762os5raEO+/Wvth8KO8bv3m0zmm7
5x1SxL8ciYzCjZj2gny6oSSdUDh6ApwQRH+DexSDqBs8pnWNhWIn9lfL6Am2jSth
o2yfiUTIzwluKFZYjFuTLHuEoXqPuV7BC46d9mFWUh6dvHCaM/yk8Tqlp7fIFCJP
JL6of4C8pkJtP/AiVdBhXUx4/sK3CYd9XZzXcs1MhxwMNqjGv5iYLw3XGL7uKpmg
ujSHj5NAe2j/HMmQFUvc9eXUIAYvRoNg4d+6/r4HuK09eQNjH0T6Y8DNFVWJF7Eo
PzsCrsZMn96gJEPz5bK6kcNfsGeL7JAmhO7nURuZsT2XETTMLtu2shUfJo3MNEDQ
O1Jx7Ie/Wo/jwpWZvDipc3rpcHccD0C3/pSBogCXarvkJuxAxJS3q/X3BMzIw2Z8
kXvX+y4iY6I8UaJLH0j2EjyqN9JaLzFls9hawi8s07ImxF7Qv8l7+nVgnqlLkvvu
zCYI1GaVkrTwIjD1edXR1TOl7XuncVizj493/o1TdPuC7XAPClOg2Pw/GAuNVS1R
3kYhSzmI1SlN19UmCe9PptJECirPbS24C0z+6AQPZgmL46lpEAR2jtR3qTpJkFUp
V0YL4iEJctUh8AqJdbro7GJPRaZw8W5ZNL3KsQLigV/T5IfYpR8U7tUMip7HsMv0
Xj8DNzfLRnpTFFXRuGnDcGA9RCdgMxbOpxbx/ipTayvZAVXfMSZLXc2z9Gb5lx95
tkkhuNk1ljPm9Usb+DiuAPCUaiE2Fn8zCNoNEBPgq2Vv4+mqwuBQFptQLyHMbYVG
hWHLT0jL1TZ/mkVou1J2VX4ODIklfUdRaIcCE4mkwCNUDr/g2rHx8YaSEoxZ2GaA
cntkNsCQhn7DJ3bYCd3JbDERpz8TjAuHy2DUWvapo6AuMMksJG9rAFGdfGiSAGnO
phrprPf5/BhCtyfhUfd7oMI5kxfjdKr54nukGrDO91XJc0lwj3a6LXAbjNqGuKvZ
AZXJaz+mdOXEDC+xVaRSUMURrRsd5bYObrRVcWb1HD2R98yfBPUQqD0QvuRqujFG
tjHbrDgXaAir6B+A6Gxx44v98YObN7y0rGsk/11zgJODaqmn/QEzVmbvCMx65tss
xCx3icY4X3D70HlkC7fBeK1YnAxrlZwFzCKyzKHO5paZny6wrWX24eSpnzEZvstT
j8WPsh8d/E2HXO6efk4e/w7kg0IkfH7RBEQknoWF4zOGR5BDLY7ndoXlY1lLJcWF
pClZOJYGJx6rx7JE9W3sV0xjbQh4aDaFumGl2Q1r0JUusC5obcKsw6EYoQAnL+qV
E21GUkUElWswWDZlgDxXGcvAWX64oyWtHVkYqGnHO1wkqZlOBuB+TDz1HsyCQvrq
3IKtu+tQ+x2XsmaYjINg/HyDiyJlfB2VRcm0Y2cxBGZm03p/wCK3RT4grNcDQLg9
cRIRY+M/lQX17ahOPz1gEpjFVP2y9qjwYBGZpjhXpYwGr00nF235GR6mDppmfP2U
aJcJ7ONDjaOGEkqEj6uPn3RC+IXwzbc3ucrKIS7GAoVk42yR33EEgL9Wf5qEHMgX
JkqW8XEooiackHMq+6eggezzQrwYLcgloaqF73QdLKDet/FXEERBzDaxD02rqDUK
V8z1RSehM5HiVxUTgurRuQRqzxzeC5EN2hETtj9H3Xdr+zx454UDTBIUvFc/YZqW
6vT1fL2gpS2MIsnpG8vcw74pwIHKK0AxJXtYY9aJ0eRFL6Spq9+NrBudITB//iJO
jtvCiV87q+PTDNUgtLcvLmPKDUqc3WZtJWdmHemVjmMfDg84jAamgYopj6mITh3k
HqwE/xPrwn2zi76q53Miaj1UJZ+zTn4GtHMNRh3kNFwhIR9tyEnGzkAAkxudERdB
MUeZLuq2v3zi6MU4WNJZNydtnvHveqVozeAHmcNeUumTsSSwMcBl/gxbb0HSTI1O
QAq4WhK1qxalF0zL4WNekSyvaFceDYrsEcsP/IYWweVOuWcKtuYFqRtML2e34r/O
VMgWgV60poWyOwT/bsFWwQiOUE5d3vUqhN2QxVBn98CETBbuSuR7rQ+i9jtMHMan
1S6fqlIvVDY4K3v8bcMdzLznXfBnXD56/3R58ld0Y+wyLvaCtL+6idX5sv6ttEhf
uFEU75Iijm4nsiJCYjqpt0izCf+keRitZA0kuiO8zd7od8mBwG7w+t2nXEK9rDL+
y7BPTSNIcy2FUqqdccZ1OzHqf1tG08NERVArCT9/yTKDk4Ky1+3OxhoKzSCtoVyL
kIx8XiQMYRGJXQoG879kM53QK0qtHfrUrlsGvGOaxWiZtradYzAyEpjY4dIZelFI
on+FNrIN3rGiTcw/pCSjafQlI0Ewp18pm2mgOVO9F1/1YpN9OLg6H+ME6pWBJrt6
dtdtmy5mlijwowU5Hijv9T54JzdqUY/ERvSQwKUti3ou+P6U3ryKneEJAJ0eh/G5
s1dJUHsDZ//mRYNa5MFz61uWKQ9lyK2p+UppNjv6TXZLP1scU5Vw7/IP6fgTADhq
FP4+WgN0JoUk1wkJNHQflAWvVG2Lda1ZPuIb9rwWpTvmmmubWBv93CLvosmmu9PC
G/Bt2z0+SxVUPZEHMOc/khpfeMCff2N/W/bQEcX2MwzbYTfemgV1CVii5YkEbawv
6A5u0imIfFmqKReya0U/jQ==
`pragma protect end_protected
