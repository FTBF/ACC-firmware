// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 03:56:43 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qeDYN3+fc7p2lYo0Ai+Bt+jVJt3yI5RF7sjk51htsGes1c7JWGw4ACQIIZql33Lt
IzX/W2rIEjo8kZiDVf5+e1sqteaz8Ilj3A1uqMWMRShU8p2mHQQqDj1nyQaK7eeI
wMpDR3/nhCwRNfQKHyjHX9nQv0zFgnstL+ag5/Sxh+E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13344)
eCdKyQlyWo2OLBkZE0u7T4HuLcAWVBi0QQawIoU7wj0twA3xMzcLdaaQyie/UAmd
x5rGgXmFt3Fx5YCHT4gWkeKzaeJWpAlGokjxRoB//Rfxu9l2qTAdK7KuTAhb7+Qn
fuiYdwqAK571m1XwzeFBGMH4X2pwesBrv56kj1MmZHeUJXr1fM224tEUyC7R6usG
+tmg2XK/CSHskRSSgPGzXLmL5ecks8/+WqfwcSkoD+/PFYBtJx7G5bdIkEu3HyXV
NKd8TAPLtCuvPTm+yuE2XhBg5Dxke606Vjr4J9hmN4pwInUMvUwABN/RsoJFt9AV
ySZ1zt/EnAHI2v1DKqnEVsxYUdlw1RjYXlnfkOTt6sjnrkh//N/pXwaa8IoG//Fn
3PftJp5sKMvhJQzmm5+fFvJIFFwB699fooIs9Nc10DftIWVBSIdEJ08eLBgAwIK/
c/kklecpn+sbVmmFTslDv9sfkMkJ9DF2kTiAQaJh4Ukb5A9vHIFBS8tI1U1uwEj3
Y70qQP/3Vv9QdxspWomaFACdo5NAU+FWFa8LqReKWRF8a/Df5t4XE8ZB/NMsXggy
YLNsZPNJqTXDLsengFfkggvyFeEtrvVkNHNhmC0Vg/+3PdCltu3K8bM3/gf7oI+t
6ub1zxty2ZVBvkyBk7aRQsOFG3X8pZJjOujYl/naySExnvU5BDSU3G/8Bq/Lw7E7
jgcWctSlKuv0570jbeiy1MEFAB1K5UyeAbPwHfLd6hPigSS60953WuOiop4vEDFV
8WFHIUPokpW/96mBgqjOt320cjqowgjqVUFdoIISvdknRIvUA6lOBT/fMRQnmF7Q
Z3QMRRXu4Mf/7o/KobWk3xRiBb9UYu/dzh/BCQ9H1+Jd+Fc6E87cWurXKTMXrznl
Dxzu0GtFgqTrLlk7qL8dUrxu6MruTmhb02HKVqTzAkpzckRZNpxbObqoCiZLkKak
QRIHMepVoHla5MjEy7JCCkH9H0QRDJFy5Gy4bZyB2aAhA6AvAi3bfT46zxIlE/qh
RM+3GEoYBp3cQQVOJYgpGDs1xS69j/gUJENz9YkTFAAOl3jl6idB5/NS/QiMjCsV
Cgf9WKzk0Bp90eYpJGUeLWwOoMVSQ3OfcImQS8qxEsLwMjG2kdwl55Obb9JhKnZv
ene10nlxInvI8J/uq55GzNwI+uT2p3zFRka1gaFXtmVgZ8YFkm9UQ2dMQft3j0nF
k/55XhkNDcLXQOlYepjcDr7SvATMq+exN6ApE0JWDTjOIvAv+/P9A5MbX8Uu+hr0
W6puVc50FIkNGZNvJAybxq6UPl0Y2ogKi9FJeJIxnbUHw22Ri0AcIJyEvB8BnrOP
emDQGlcOIJLId/xiFZe0UsYNGlXhr7kt6F3uqtlEDFnjZ7qxZhKhL65qrk6NDfR8
bJkJWEWHSiQPwIBLrChs/Eg6bsnScKdW/BR840Y3BgF2GUMqRcXvtWYe952/H5J/
B7ayCJ3ZqFkYhxGSi5UqoWIgXfzLRa1r+3KrJm/rWs5tEbuGNjLzD5M+LWA3T0sh
II4aTYvpD6pVxV6VGSeidL6ekAICXAttz4X0fcc/gGAWmhj24jbrH45vf6worb0G
+jfh6Q2GD06QoSUxiiZbEIlLNiBLeELODGO7W84ffkrw7Dea84fyTUkRG2YWUEG6
QPU8EuhshQIF/RBooDZWYF7lqGDkVYSoxNPfk3b1Io/MKx6rBZ2+uRkJumSh12hG
/pva2MeVa5QhpeG5wSUZh82bZHgfg78Hd9XKkvay9gIJFq6XHu3ARydbPsrpexVB
XjMFJWhVBHx2mbQaIhq796JOMbIGOmzUJRy84tGnT/ymVx3Lf8cSaZX68SrG1ppv
qCeGVjSsZ3hqzlKy9Q/angshQyWZQ3PE1wgC0x8SAbM0HewPd3Lk5C7BXjBUHOPj
pvC6E7ERGkEJqOunakG86iqQ6iFg/1o1A9Vg3ilUwDJ3ps0AK8+IzIP8xjBPzw0y
WwaCpQ3l0+Og3OQB7QkJrUJcWMBJe6j8Y2PFUbr3NqgIfSng7svt7R+I5smglyMm
VT4nr+j6nGdadnJ+uEZCKj3m9W6rucGZRnOaDhqKj3hrTVRRbpXIh5VY3vWbbqjX
r0immmLyYT6nmH4ZavDtv0R2OznQZnmxPnZ7zTiKRnWXlzSVVuWvthUxycQqnefx
rMlq6agkOjKE0jr0HOKmoGCmjqBpRR54LmX80kMCwG2ItBlxZ4rR09HyLhxQAGqH
eeL9JgMKXkn04WC9lr61DTBfC1rjmPqVNlRD9+vKwKD3LaIJyIFj5AZ4zAqJX5sA
JTgxSL+/hivFG46JFmN3ynPXdAGlfu4dhiDEmWpVq8P8xmM3LbbH52qElGz0oD59
7O+obUzZKanobHHbyS6ChHAZsULTJEvYhYyxcfwyS7OkO/xjKEEKp24Dls7v7kzb
akdOPbjjki8ei8mnNCQET+x69M72NkTHHfjGHfY6ZoBLlTGX0ufRdMSz7RTuTPNa
eXR2i0P+DJqtUmrWgVz6+gqdSNsIMzZ9b8/il4mhJSEs8aDywGW2VX7xiW0nbVyA
PM+FN0UbliqJOoPL6BfwRL3tiOYiyq/J4Eh/PYlsVXs4WzMbSLnbaSqgcydQZbyg
Y0RPTBEIAmQLwqd5erFrOYsas8WXcwFF8u7o68NVM5SoG6BJqu1gQZ1LEyHpMbuD
IjllTkxzxWtB6RDrJOwQLtJLp1Fi0H4WOOFgdUErDB9m/h+tXGawqpl41vq4BTo1
YrIwiOSB3f1cW1Q5YQLsgHqmcqNNbKlqevQ+jPGLDRLR2xlRjURoDgd6xHjliRq5
HMUxuSIRjFy5lh11Px0UQcyfISQ+XMOC7+Yni82AHISUAe4Jxf8sWSCHBSKFru+z
64KqaJBAvscNjxS6XUn/pf7cMMtt5aCP7GqIVvxn5eRswAdzEZHY09cZnO3kTNrh
wEq+d2DZ5gEx6yuGfznVM14DOawv3TWCpZdbnGu2OWweqJMX1RdaO+TyymyzgdqE
m3rAXZFrBwC4TJLZXcOjjZ/rwumefeyGadetI5ovMPnB1sbryU1NFJ1SEMO95t07
lLWVBwSem6wjRt8+bnY+jBalOphpfFGU5cqafhAtFxHxwFT/00nd3+QOW324VZC6
jncOJL0wKRKqym7iDz6SW44qjVE/AtN9m5K9KeUBWnDANztF2lEQc+x537L4zCbK
ntho8AwX3LIg7m4tel7xvT/xCTDGI8PLIWZ5PB8ch9n38PBKKjniM45z7dWdKjRc
ym4DhULbBk4xM3U+WMkAs6Z5FkY1fRm1iA7yHIhsOXC0K9Gl8NJaDKoY31a05/IG
bJrdgasfYPbGzBjqq2QkOCAgbV5w9H8L3eWRpPwE7Lyj5rAH9u62fJIsnL6KH/3k
nHIxgo3KLvFJj2eHPpJEoBtCEQumRPf/QFg/m4WC08wMvfOm09PbBOEyKYVOgGqN
mry6yZKTHeyA/xod7NvBU/IZTW6RqB879c+TwbhDzGXn6RlTHbsBBeEVpO8SqQun
cwKDnVpQy+X17kamb/5ZUAz/Ir3EFCMeJEdsrv+Ime3XiwOb0F1c5J4MWbjQKSfG
hqRhYVWw/X2VVJKZ7D+bTDoiqqye7rXQIbwdFFrSNauk4VlFhFeF7L+fdNRouebE
ysrsQ78NzrpvsrD31qRhMUNAfW5JiEfUIzmmVL3yJkm/iK0x8qxh0Oaz4SnfwxdH
kWbKPAsJ7ez64mS+Bo+QhgB+VYyxSBqVKmKm7kPo53eMYwKqZj9Ppgm8f7uVF8KF
zB4q1K4I3OrIztQ9PbroxnE6/PGTGRDp4NId7beKpEVd6QGj17NBgVDfr3+f2VN3
qKAROrLxl60uKAt2yBfFeuOPnPinqpHKJo//BYmd4EGMMzHi+Wehof3UFhBhaFVi
eX9QgVWPhFd9trC69hHHIYMUdjLR86M1XiGZMRknf0799oBf0Yy7ijiNv/+BrHL4
4h1N3ga+HiTjEXHNRjwitHmxrqjQIxmuUPira5NfISzr7iLoU1VJtFSAubgRgARM
B3tuY2Q0g4OVmbssD735Hu5kxRQ4sZx1mPP/1F8yyIzd6R1q8hvNow5FH6wI8Yhx
lh8HslZKSJBkYctvo2Y6v2E+H+tqNWcSVmO9etdPw3Hm/MDy9OAnk4KJOnWTO+eQ
DnoaF0WvVDJYlvAYRCfpnqPSWPsuhIMFlY8xrSTR0VZqPA76tpO+WMC7HyAmJXaY
5pPT/vBOzAZJIpYvDM3zvYK0kVoIsK/6+fCEhUrrUyiXJxJKxTRuYV2n2Bsmbbau
VecNXXLWtSLJ38gTtCUcXt8Q7I840FbSqzaLswQk5wR0nZoRC72TdGXtntElOlhA
6SxBW+IIIeQthhvIud+WgarOZBX2XT81U3ENRba93CBRR0p+5ETxFTE7ujF9Y2hP
OI5cNq0bMi8b0VB2WqwEgNf+N2Ya56Z37+TxqJVLBEaSzLnMdzGUghJswo/klIRN
qEEr/37XXgr/qf+6HbD0VeoqEto3bGJLseopC1eafSTSgHk4PnbpQ78WdZIvmmgj
K47lDUaNaw0PiG5XTGBkKOEVR5EAbh3ajRc8coeDlBgUic8u6LLqN4MXwhcYI2pV
XXpohFLi19RGjjLsTxpcCssnJVOdrk45CtoyqXmcM9VQjUnQ5kDbo3iAZLVAuuY/
eJgQe0s3BjPHTNBcie0vMw/WVOxC9s2/XhH+tey+S7WhCctcrrywwwa4I9j8TTji
Yk3Lb7o84pDQtgZnOqATcxpX96of3/tAYlxxYHEWLS5IyafeblL8ZxIab52Jk9Vv
Y0mufYZ/Z0RtKOLXislTaMwgkmTDbcuCruS6FUlUuzcCClPGiVJQWyfLkLIQcn5M
pP+9Bc3ulKdC1GNCtVDwhoeauuc/cnd5V9HZtgjVK7s1aV8G7QnuUemrP2oZPm64
iJCKa9pFBn+vyVI1S2u9GgTc+n5MdAXcqFbmk9wqFQFtFOeqIEDE8OZC1GK+cPLv
wGoRBNk8zYZtuVdBAZst8IB24fWkz0n6itKVcSkGBgCkpwg7yeiDq5BczOIuJ8V9
JLcagCVOknVcZ7v2lksKddrHq9Df4ygPqPp5RlDd4yztWiTbCa1EtOjimAD8B3HA
erYEIW3XoEBQM+6L34hUdmPhISg5meU3LqSAGNtAI1XoYBeHFzDzgxVy5qKV6Aq+
jyjRQhy+907JOgRFB7IrvqhpHFmmPXSd5Zl7PKBtYrych8HDxs9jqjAlw+/GW6G1
bNuelT+W5N63bwVmzSA43o0eIL7niOnrMcyg4GYTdn86ytR+NSZ5WaNMrcc32qnn
J/XckeaSKyQKdpZa6YdTPqwqIVo+TTuAywqvvKTfikPjMe0PSBZ5TgEbkYpsyl1U
PLaKEXG95alCueYKOOMHqvdOzfYTHnfMbx7ESVBNCTKvWx0RVsLFt8PIr/54zVK7
SsYgfGGeaLGmFJ6VhOBAyPmYphaCNFzlXqCXo5K6eO+81DtzQbVcaq8xDG6+OiMn
MLTLcCIyPw0R94kJeh9iOI46oTaw819Bht1e7TSfq47d1HRFih1UYJkEUSVqall0
QGjjMUc4dfUd5SraOn3cdNr/gYBxNLCa/wbkjZII1I9n388jRZiwUQsjOApxOMF/
Ei6sRknx+bWiJgFkAkXTdVRWf4RI+Rw1dHYea0UhzRIopuwsWceHyd+tdysghWLC
aSr9JmGnh9y06W1Iv383MF/RVSsM7uMhtCAnHq462OerqNWo7nLjpH35+w3ABzbD
DkbngTl/QDmAA0LLYOLBLh9OxQ8lCGCMASvMWiqdpmZiBREBrd8XCurAQYeTSX/G
ELiQF7/vRErgifKXb/raw2MUU2mcgqACFueVdJ2Z0TGlv0SjBuF6WoWuhI6UNVn1
Y1I0R/+z7vEPYTGtdCqmBe6T6YQx226HugH4EvoIZD2/SsIjcfkHYjAU22cCKDbN
5pkDq0T/czu+ewuBx6E/ugntnITzm5o8m20uwtfbNV3YOusL4SCgnrzE2+IUKaXU
se7bNGZA9W8tnZWOydKIZ+ruc6SVeI1C3JL+53GDyEZSJAEEP6ti0f6SZZZT4dyZ
/XTG+0+rjOwe5P4Ok4dTZFSEOVNrlKEKdxiI5IPRmqXTdGYDeWgTbrV2Ea0mpF1g
eVaYJMN8nR+CrSJ498t43NBU/NN/XN9qRus6aU6jbw1Nr0dxXEa/qTExwjVbR36k
HcR/gQn6Mz0CqxzS09jqrX1IJWHBuK6+Yx7hMOpSqmnggnoozHkDePtwS40p18jb
OwuC/8u/xuPGvM++v8eJw0svmaG83ifgA4s8CCY7/pZErefAGP1FTpC3V4Th/JfQ
uU9wBr0dmTHgTx/HbDToJa4hVqN38W6QRhyHjED24vayZJWiN61UFj8fXIXqovRD
VawEhcW1kkjBxkbUzSojiVO8JEMOpsCB+BqCEl+6snOUKbUcRYJVGxVYnQd2gQvr
YcvbrQ7Ghn4i1bYRofL00uGxfj1Kxo37HxGtFd9/EC/ZngAb2kdps2vip+dVPSKj
AqEUaApLora/r5A3FgZZpgXzyvHvvD5NS8fvgx/jdL/hzYxvgOCN2/Jfa2Zf8ZHS
iSubURfUKe1eLSvWGTlPtPmygqPFkSRhk+vflQ3sSKdop5gBEKzwkDMUPhjRucke
qc0vQEKgerKFpOIDD5dvOBEls6Vui7dDOOwLBVFBn6P7jCstUJ0oAwDQaJY1Sava
EQUadGwkJeV40tlMqQny1c4AMh0PDyxX5cSOf1hgGysS9ZywPGl0wtqoijFYh5Pm
KS7aXCML/w6OndZwbLsmWDPJwI0scUHGGQ5Oh7iZFOsZmFyxGXDr3VbwFc3+KGqc
imtau0y8nuSH1g4g6GyCrbIbqfDtIqz2K4g8gg5u8Y/G2ERKoSzMZn4gpGhqjRdO
P8UkPe4/ZVaf4xVHU4IU2KoUodBvbOCgT2pkBg+8QpdKUme2pJvr6SBTKrszILK7
uwQ1fx+jP7vPFTFU4zUyJn8J4gdpfjMPwZuEv2s0XiY3GqEFaodPw5SNwLgLT/6m
Q/ydb2myFKSwEW4yaZhuV4Y1apczk7MqPfLOIh0TE8l3Zwdovl8aSbu8TXHZNVbS
xlDoPjeBr6BMl71FRD6FNZc/6+mF8FZiHtr0lJL3nP7vhrXT5W/fjOnxRhhNHHvh
qyJCNcwZSe/ejssRu0w8v4bi1P7b1KH1aObTaFbnv0MZodcSLbtHJidXm1DV2ao3
bcKfjLurl4lX7cWMkU9cTAlJi2dMh+r47StJ+Yg8VpLOslzsdwy7uk+Fzd5hLwOq
sJkiqXrU0lSqLCaCwPuUNgEGc53HOYJnv9uMTHSFEQJ5SO51k1ttKjalT2mUYxjI
uKKkCsNnAdCzsWU15yrkth1Op/RXlFW/pqq9Jzwik94bA3E69KrRPivQ+ihP+U51
BIjJnkoX74T3OEWFmk7DX/tdlfvN9NZBIICF4MkMYbYsOw6j4UyLCRrwPh0yoMtS
gxSDgDIspzAVWP9lIU+FQk8xzyn16QMhGZ+QNaNfg/QqnBNfEWjnfidI5Jrsg1Ym
9M7lMNRlxBt/aeeaKE0yNdJJZ5IHEOe0dIR8tWXbtmwnJX4B/bXvcyjRYHyzAsSS
ANICAuXKb0fryjN6hDBaoQWgSrp8hIb7cqh2z0WcE/ZoE0WmYv+czl6p/uNTXSOr
OQc0LRCJqgmUgpJPB5bxcWrOLcg8rUsH0m2mODMNTvQeEjVV2o/IJTfKESwMkpu9
hpJ3iAczjcH1dBWDKuP/cm3+OgOkcD2QQBO13TFGY4b/FxQ+mCojVkugjiKwNECG
0jH9R6ryxkNBcP9Lkuq+8jcu5XkISNW9IgP/IBaq+PdjzEXuyyM6E8kr9c2SyKvJ
pyIF2oMSp0/NdmMJS1MrwamXhwPEYP6KWSFPmcmq1rjs3oZJUEDA8ndOXVubzdB+
jL6EJLcS3LdNhUg7/LLJOqmH0Ki4N8KwquYA7kZzr/a2EwUqgF1HyHtvhk85aJ7E
8c7cOYd2aiPp7NdJ75wBlhYYhhlUupyjVlvS1NnTUMr5KRhvTnCRl/MeMsVgMq8w
VD54MbUJ7qzwCEn+M898h6ZWYGVppTV5dUEYKbIOM7G6XNKxcJrYyOfxn8jgXkR0
yT91vGaPs8sFaRzk0Y5csvBz4b73Si45aX/9qOhm2xMU3W6/kQ6lhtYRVJy6W/YR
9/L1z1vr4SYh32x/Oh1kj6/kRqOPa5BL0TPRcgtiyB9dDq05XLEGVcW9Tvyjfjka
VuFgOeDJRz1MtOGJOGJIbqmcRTT840o2fGtC9hUPCabD6OkCNTfn2Qk6RsOlsn72
AheLERW8tGsA92S2zsADg1ey8jw1qjFsv42BqgfSryuvfLctOiLMOzf1Kx2ONM0g
uqHQVWAQANTuKA//FLlg8UWhdI/KUUF4BLlUYerOekiRw3qsBYx0DxEkOm9jW3+Q
Mu9cQAvsVuOHVUfvpHSQGx9M+gbI/1+NGqn9TDxrZZJ9+cFVoMZtR70mfEFfTovG
iZwR2EKglSqBeAAIrhcQjfvjx7r3r054iaTEdPEdz++fYGwhz/X8H0ZMim+jlEtM
+8yRK+D4lWBY7djSMdc35loUn2g5A2R6uhdv9OHeJbxfvMMhLDH4ECyyF7tl4Jui
e5Bg2JIhwP0h5oGf/UDWjjiJI+Pcj+9rJsnu8oSmzoSP5KGOJMjFJGY5TKeHW+Fr
SZj5Kzzx8RXpT5n20vVH6eyLIRDGn/pif1EyB1cC18MMWpfjpMUEltD7VdeA5vr9
tPRUhGkAA2UpyieWpqhqv2KOUP1y+i7Qobb0K7C3bm67bJ5qYMwDD091A0r+oDv+
8coPz8xRr0ZxIPOE99H18fvnbQ1/595pel8d6Fep5gt8NGUrXPCdW9L0vcBokxda
DE01T/ZjGWKGpZ95ragBmgWwH9vfol63mWb3YilMYhHUFxdft0sCzH+fF5GfHbZF
guNTcnLo9sxRCNun6GhSqaSBZUApFrytRMrFQovzSNwS3s0ChWw6iw6ODgKpPG7P
yIESL1+QANZUC0mLxZJteBMZLIsW/WRIOjV3/f0z0ULTTM3s4cmDZTt3XSSJ0N+U
EjzYqs+aaFY/poT+wmkMOw1J5GRHeOJetg+hech+AA+O48Bi2chyRmSvoF8TUuhn
yUCXn2wsoqRXjN5VJ6ZjaLEmYqq49FGAwoshQwmGz0l6fGQSPZBuVubn5wq012ye
S8MPc10qcJ0v3ZVSZpELSQOZNjEskU7295Zvy1KXnA+YCOf7DY2bjKT6fQ+lP8TZ
32AaqKz9LUfSQJjSoZSSd+Yf6Nl0BSrsFTfts95fs3bXip6DfKd8Qgpatg8BHf/Y
3kCRj2k35OKjPf5hV6VfOpQjOLnvipWEjIiDNPGB0TApujz3nHfod4uZ+DV25jiE
8LZWe+cjpoigCecWv8Kqd8bkOYlLUAzjxw4blfWaoT8jr4RypFNiTZ5SmLrqzR/U
ATrfPOTP/5pJgcTJLT0gVgZFzK3+J3zspE9df3upQ5US9YGV8FIT5JexCuarG62v
+MBraf7+lNc3J+IgvV27cTrakuPVD9Cfku+4AS0+umq81lqH9QTKZAQf+gBSqDXg
F58AIcWey8/DevQObFbepHotOcSDiNhb371igKU0zNLJeVi0yCzGApXL1pSuKTRw
dENQDZLbM5wwtXEwhBkHZhVZ4/xJOYMrdFWNhp+FyGe5qKfS3xCUe8XwYFA2G9uT
KUSNh+DCOZcMeGw/Gp6U7HVBLA4RYLi3soUv62HzidVXTJOOqYlRl4DLNzJMUEqF
4j4n/kQcc+87JwOx57A0wo7KifRx1AHim9WzbLQGFcfW6g+TeOFTn/ko5XNy2jwK
JayyjNgbigahRogS1oxbl94y9t9bPG2z8fF1PexpI/MlwVBvH4Leb5ocJZivl9BB
9erQornAIDca6Xx0Br1pIFUY7FaQvLuucQ3kwtMp85Wgj7CUylE7aI6Of3dStqZV
YXGOt+XC1KW5UBwD9icxpA0W7Q3PFrf6W40WsTPsYgbPtGBFbwYqYBKnKm0JPBE6
VUy3Mf4BKAukBiYy6VFEorkKVqujdcspL8Prz02oCXIo/8bFmkSnVo9VW6rxnlzj
5P0DxCkt7LmOLCvzQR7y8afAWhETntxCdut0K1ekFgsIpevt6geL3aacVgHlciR1
JK+HUkrnsmCjmKSz5DA86IoK9yDf4Toj89qQhtvpTXwzkFJeOm8XHLTo9zykpalU
j51oIHii4wAynOZrfUES7gUcPKf1yViN4fHGxfPh1pxXUC6mJOmot+m+X3gAcd78
QzqiLjHx1bBs2wxVDYi67ypOq33OzgnmqKg/mk7M+Tvq9xs3UxU5sy5u3B+d24db
vFkE1HsMu57m8G+ZSedsBh4iImLDTxEtiwN+ikMCGtA6XdTQU+XA8NX4xy20feQ2
80mfQy0MtVLcBnqzNdQ78RIH2GeZWk1svhzML+i108XLII+0l6plKsS6H8mmVrQF
v1izZQrY3XxlVcitbS/ARDoam4xqIZKWC770hXVqMpdnNln2EW1pXYmeTUWYRhbX
RW3sGFMt9XhxwsrNz6j0kjyCbFtf6KmF7KRewLxYCebezRUnLPTeL57Gb2nP6bAa
73tFyDHam8yImdlwVszko7ojQKBjISI0zBC8LTDGMvnPyIp9uuRTYQiO/Yu6hCHK
K3tGjvLp7LhpvNZ6ooQBlpz4C2vEti7MGQqHdYszDoGrMJ8lzl0vcbk+HSEki4Bu
LUb40mK+gFwDp15E5XmuHZQafaDuLfAAN2w3aDJ+TuykrYQIGsmKtnlZK43g5mt1
60EboQuAuREePX0DEgmPEFFmX419DAY2ODxX+uoxokygCYrXym/whpsYDpn8nViS
JOKIySR6QHvFILpjSPSBkB8hIzBEC256NmaRKrUZVk7marRkPtXUE4OpvqS2rnmN
IogAdZ2vB1FfjU8p/KvBAAQcQSBzziKD5bCpnZUtqh7Bq+BL24NushzyW+B5fyzU
UNr5Elh933pAMpEz5t3rVIg+DHmgTXDxxS8BLe+Cep9mcilzaMUPKil1SbztGRjs
cV3mGsFWgss32+HmEPPLmpje671hihA//6QvXHQkuO0cpNDbJ1CK8dF+EIAj0Ouz
iEfT2e26oxSHjS0dTH5S6hB1fwknCfEF4bQFs5OEDtJZDt4AKCQNK+hLD8K/agCj
9Kbvm+gA/R6aQjm4D9+5uSMUpwCSze1xBcyPDyuuMqghoY2PyYxgg56FX0HAo6v5
kWN6Nye3wXp6P/QPJ908wtAxx6zAxgHj7JOkO8KcHDDoV28LOOAmuLdCPcKZqZh6
f7t6++kg65o1mfFuRCRyCq7nNn97NcMGHcGyKPK49rt5pOfK39/Cq9FIVBRiB54b
J8ZjZTv/trxGL+zuI8wRByFb2gKD0IRyUuEDObhFPIF+ABPhiLWDakCHJVOIhjSU
dw2nWOq0L5KHZXLyKbjX0IqfjoEZbsSQRQRU1+1ZaK0tPoHrXkVgSogL5VL+Zm3s
sk9oTdtZqyaf6SmxeDrnxAGAoT6+h9fDu25+FbUSHKua9eeeq/sCu4FiLDyXYpQB
Liq3xScRrV5dvqieV+6zuE4dM8mPO90O+yIjdPw9ZRWVGyN1Im1FjvL6YCS0VxAY
C0uWRKFNNArFdpGu/JUuDN+Xk16GkN99Bddhr6zGES/gyRjYSnsnSGS24zpC7KY6
AF+W9s+RDqNYAPNK16RaxkAU3LNw9qTHUgjIeFNoP1dj65dpQv2yv3j7shn55rtk
hrRCA1wiOhVq8CUiGGjI/VgJjxp9/yIqgHHp0mh/Y+75pCBy0vNFsfw6ptEiebYN
+bka1MNYWvxQWMAXGe/0TGLp43wwH8N7d3SJtHu8Ct1WvHWOxozBKgHe5rZFfqus
vZuD7vXxGabW7O4SBrXs18YYbkHhtfA+PvNXmeBfDUWPgavvFEPYkQ82M0onrmw/
5z7xpp1bn2X6RGDK5Gnw+SsCYObIZ4tCwX/bNmTfXMcBORfowH4QVFRJ3Ohu3va0
ba+32jYTn1IAXRdiCHlP4yCjy7OdRSueDWklwuWdoDY4owxgoTMn8yARVNgI54kV
FUesP4fg7Us1gGvxTmLXtURFhGy55zYI5HEUeqMZ92XvcIkChhYhgppt1aoduXS/
h+zCXkmPMIRNSkU83yu4dn+2hRuq6Fen+5Dpu+XYTBEpT0wVdsXDrCEGkp59k54D
beZpHfswP5bUJIIgklnXnHZroPfgHnkqXduL2KI8GfzdLf1igGk0U8PLxSKpptQb
OCy+JWB6STEFAPE+OiyoultYs74MEy+g2SUw92p5bmKQ/MbjW/KlVs56Xa7A6AG3
tahHYxyvBjFlvrysME6BHMhpOBpGJiR2fx9ylAy/dEFPSDdfy5CVGrEJN/eRH5uo
T0rFBkVD8ZLJWNVTv1bRFnyBCyjoJe2YfAlITxPDnk1zw/QmiGFtm4Vrb4GX7eOb
tbDP5EuLJbqBKHQHeh2wwxltMS6lrACSQy/4e2yFem45Og/MmvwYi+oPOruk9PGz
3LwHczn0KN7Aka4xhgN83jeTOjHsDimuWCpkENopC+T7rSDIZ2b+DJfdZwkS7Koz
EGxOtHUhUHDrUoP8KqcYv/OCVjJ3bTnSVyR2ogYwHLmG48Jfj4w5+QCnfk+wqjNT
VX1T5omPXCZ23y/oR9t3nr66unp5MuCEGFPmf8rZsDYocKwFZifZ5LOhb83i8EEN
ZU5Fgv94/A0WYXanT+hTCija1t8AEWzteWp92BWiivXZVv9X7mZn/ruqh5JfvsiW
6V7oM4luZT4WL3gNzh3WpXLXQf4Axi69VRNotuPx2r340TeQ4ii5oCNLX9B3rAfo
WrXUQ1S+1TeWzBmB6fw09aGnG7/0wweNacrUYfHPT3C8LFTQife0TJJ6YTyrcu/9
QpgxPNgD/P53ZRTSB5P7E38GcdnZtF7jnnsi4cZjf17PP+s0z04E2Yi8YPyJk+cW
3c+Nio6hAx2cDQ6U0Q6SJWt/2t+tmnOmEjEx25oZoHYnTUXt6YoT4KFiZ5Mgek8x
naEB9RzFMIgDYaeJHL5EszTv6VQVw58DljmadvNK1LYjA/48s9+YCSSttM1nyuZL
nZsDBmZD73WF+Elu6eQOU5EhiLqN+n/I+3rj9M0M3bEx+FYnDfUfX6h1tyI4eHIA
oYNGnC3xIs2j5+8kBEcpJ6GORnJP6YHixJMDDcrsyDHp/x4riv/+SkGcPZyJsGLn
Ju7+O0jnsyLAcqeThrvxJqV32t1nfWdUg53RwlL2q1klsoS425BeCFeUrUES0Y9d
qZbaSlZHO+3VNqSwHEgkvE+hvQr7/sSFhOLN1lv97KqH6D1U+DCZ0kduz0HyFB0j
ov72D5YDmvPHz/u5Ts2EKNXYTlygFNDylwF9x87cAuksbO3QzAo+lj1JHvSV/ONz
IKDmnDx3E8jkDpsR/FhK35C2KK5b4DgK9WoPdnDL5/u3F0u41Fh+mME71eiY7WT9
50q2LiCu6nItZHuEQIocDtiCfM1uLQV+a5MZr8rK0tVeQYamqLFcrEOAwW/pteuO
6zpuIdNI8bzrvXB3Jii9EN5on8TepF9ZNG0oICHA3Pxok5O9SoViQvmbBM6I7Iwn
xWaoALODx2mKxjuUEuEvariMLwW9mfAgLfZorzwDkkT350Q9z8hMeqcrw7NncYuk
TNeTBeuIPo2pAinNB5Gnn/xeVWC0e4UsWDnit8n0poO0vKmzs/YflrVQzH4fYfJh
ykyziUPnvvCr5R1dw79a1pIO3JWXZMiGuLUU0SMJX11gOOk9WBLQQwgpgsZbSaCD
Puc9AU38IqRnpNtundNWcA1UsavX/ROrPpygEVlJDmCJw3GdzZKwEFi9rzrhaupK
0mZ0hXwI5CsPw2v2IeytL48EDBjjHvsMEhnDT+F6UmJ3aYI6+m0fEFT996vGfsi3
3D2NSnufvIcTEHI9COmWzUKLtfopOZWd6Y8wHB5Daf4fAmAgAoLxFtErl++2g8iD
LrjhQFQ76k82bs3qetdEeURCyWi0mRSnTE9+F0jvbL0NDEU78fJwUqit4lJt+D89
ewitBYjtHgxaFkA3xKPW3t2knnC4PY3/x2+2eOXJg7BCZeqZAecVrzWMHpZWKSgX
JCo+1TVeo59ojKovyF5HTlQRt7Cru2ONA8+aYBuZMoQ3baZi+XKlWCxtxJwmWTWA
QZln6/e3CQjBrDNqBnPDEV867+n5TdEQcr0xdMUZQThALjprQzlnctuhwuu9PtYo
U3geaLqgE4bVomlxnE/+euHqi7WC4EipQqmgThCPjDoJV/gDfN+rXfynydDfdPa8
Ifw8hMlb1EWcPC247Np/hMJNMzBa1hkY2SF3TyTktluBC7L9aMrQv4H9XOy+Oaxg
6z4TwpjP24zH6N0fSUTxjEVtx61G4CTBAVpTaNZMNuPIui1EVLkOHNN8u2r4BUHs
ImNpMwgKcwp/oXiSzUnh10fkgForrYHq7MPwcZ9ro05Ju01LmH7P/cFrxVL43xlR
9zJHe/QGnG33eiHSEdkFXRKWY0qRvUa5kgK1ZjuJ5iDRzRX5vxJo6Gr9cjVrfQip
fK+9Txfl/8Rex+Jysj1CGRa4blzTMZTu3mnK3RTydX01MkJqb9R6RVAAKg1J1SJf
mIaXG3IhIT3x1umF07aDAXlnjwpqJjhDy3W8UPqWCvbFg531YM1fvRuagKWzow2u
13L6S3MT0npLbvzjkHb1X/UTUk2Pnr2rY40XC6OnKSpcWbgoTJMS6UU4UK9DEldM
hEWNudf+WNoqegpS+IGcSr9JkH/ZM9hPYKZ+WtDUA+8+4Wj28pjgwlk/+YkmvjkB
z1MzhBhJxPa/PlRkA+fsmfbiJvkjGDv+JtM9LJJSZTB32fvvywu5U/KIf4Me6fFG
EjXPwLJhtKy4g2Iejl1HVc2TdS+ICj0N8kKC/Pu0GYiqK1AHJk3wMr+/6fRIThJJ
vdv+R969XYGD7Qj3mStFKnEckiRJLaWgiWNLTt0yT+IQVZwO41PrgtaOhRwRr5lm
Sk24e0MLQRxQAF9Q5i/5zuYosDEHTYPVDo3J9Pc/c09y3aB1L8cZt9aBxz5CV0mg
CvKYtv1jDEfrcqhzHzjeuQNNkqhD46g/vqxFJE/RFIZZmS49VYiQfMOb2NOmb56R
i/Jv58Mswc+GzMxr1KB7/On/DMsVop5qKXzrVPCh9yqBwvkksA1UXQsp1R6FYEJ5
+JPtmg4EIIZ2ahbMTtceWObVGRgwRB+45ITvxcSjQQN3BygxZVgm2fI6MOFvuWsO
uTvkQ9IqPYG2vOAHgeQR/wYVlxwTJmrA7MnYGpiOfUW/eXEhJzhIv9E6SFAj6ljL
AiFe8gAXbMSi7THZO/WE663EN25wsW7KIou3DstPh6PxGtT6LjfpDiB8SNHaDTBL
cyClGU5aJiLb+sePu9EosgykUb0lQbwjEYsilY76CMk6RwzysWVhHXNgj+iuinTU
pEtnpCfhrYFjL91CG+HDYLkSIS8Rx97uxPo895vy8jz7w/M5X+kA2IeelZeGQv/H
/Kco6+fawwNb74RQAKY+j2CnCmbVEB7rULXEdFaqKUpGfb6Xta/4XmNHeTuG4Jvz
7UavekdkD2e5XcKBThLARyO+Va530yJATmXOMJCcAL6rFwH8kIJjsWO4bmzNKJY/
hOhuejqCy8PgkfiC7oujLkkw2gvai5SuSbK7nlmaVhst2acxAsA+ocAUcuyEAdoD
uhddTnszTIQnkLFeMfZsgao+QP87qUhXup/Rf3dpWa/ci85FQur6kueXpGqaE1KQ
mgBLPXJHakeZmbyCl2FIE1RdGO3CLNGF8tP0d+2vsGkdECdiSv6gYw5LDhXXqfpv
oaDkom5nEBT9tFhniL0wLalXglSa1By6tztHzFiLdUsYvFOZIxxAbo3zbshmMnH4
N23c6FWg1dFprXBZMNrmkLtFKBn+6T+rY805LYNFJFd6VwERfnmu3eDql5gT6ME4
CVFwbhGENd/S3+XbzlLZDmlS8I3Fm8HtigV9LSUnENbhw3lq4oHtIsjycngF+3kD
iXMZgKCp7J/wmE8X2Gf1W/32gqcEZ2tRuRfm4kZnICQABHAjBSLMQxxujb17pVMR
EbALDyr3p4YoZJBgiYSl8nQ6lugTa91rxRrdQO/jsRZz7bdy+rIKL5tVbeuO16Or
CUhMUzuGtzygVtPwV7JWzyn9ON9ixQh/tLlaiyWcNx435sIcAslPebokipAeTqyU
hXqPIdT0MzOxFZ7xrxjlMehXi+OCCy5s4GxFB6ocrS73ojRxybV4y4HMCbwR4Hte
uQH9EJxNirQv9VsOqUf4xiEtoaTC0glS1n3PSccbB2Gt7fb632w95MFxC1l99nPo
6OO6/u0Yo+3P9d9hNFG9tJ93TRbUV505A8D1f9kX0BzyLC7yHT9iw+7zl3EwBgZY
RVP9V01wCEPgDck8BZ+5HWNo1x27DV/JyNofEJ3zH65cmbkVWuzin2BiONFBw+c2
7tHdgDXablEj9BJkOBuHLA1L5SHC+Ou2To2Aj/NioVqOiMuqQkEi70kE0L2bexwg
FoTeZIMPfAdk6zvCP3TqiZax18sXcxcw87YDecWqGMLobVBU7sXJCAz+eQ4kmPGf
xX1v2QLH5T+oaM+vawXHXVCXor8AqORLkKBejkonYw/0PER+TU7Pxx0QMc2gu3vI
Ef4Z5hXVoiIPRHa0ITApwLQ6zay1zRBNXJzRr3OzjFpf69Q6MjLorzqVxl2W33bT
r4nTocXUyvnWAmEsga1Y0mO5AmiAZtgZ3f9n87098T/aiqk1oFLh0pJDjHTV7R3g
B18OZ/q3klxhJ/P0KsRF+AOr3yXUJy1mqMvaVH4HnXypZdJcrf0o9SSOteIGfIJc
JYlhjQW6JwIYNsoJbXdilI7FY86sMA75NU9Zxro9ErcUgumAvxd8Qr+0EK1ZmdJa
NhzmhXT4++NMiJl/UtZODW6/8B5YtnEBmRrOzRwt4iJVWHB2m71BjkEfkMT9Qh7m
OLtfrWe34w54oxE5piU2dgwixzzRcz8uFvhoL0xehlxDpMbo/TjdwlOSkS2LfG+U
duFrmFAQuW7LYtL4Vq9fstSzNCNbglbPYhcn81916JepxAlBQyfyDOB6Ty3ZOMKp
9FTBaNl73uKs328TAMrPCC5f7EXoMC2DdfjJl+JICaDpRtT8WfT7kIDTFhWrDDj6
8QnzAM/Bg9J78G5FMxv0/93Gl376pA4WwdDxwCAEXkq53znIxRbv/XC1LaahuOt2
E3uJHll5T70DZ7PCTgfhf94pjxNc9zmfm1FVXLuzAv91+uu8b3zxtjG5wmRGdvwg
UiU/JwAPWtO57qmbe29XZcsqCAEeACoyw/V3fBYYxXYpT+dReKF517DYhhGJDR8/
01yqq/CwwId+fenE4JgZduEmGui07vFUcP8HnMlpDsRpgnrSUXhdMytaLAI76TuA
t4lCwHO1uZNtR3F3Ax+k/7eZsV00/EMY4bMSoVkS3qbFYn7i61OzTZ094AtVYH69
ugHM9qYttPdcjIvN9J0E+iB2PERLNn4arX7Ysx6Ytn4meqclaMHErm+5QUodiNwk
P5YbkPfA1hXBmdJXEBLogUIk0Pm/NZKHVgy3jKOeoLSeU7diJIdsMTv95JdWxEc1
Q5dqtJiSqWgaN4kXgt6yTEmDoXHjMS3nlT+2MyGifjjmPFI+PWch0AaHAZIgRNH6
6I1FqSnDaEHSSs2WIQAran82qUKKxTYlZ8vrniPFozgp26igStB3PVEL6HPIw/nw
`pragma protect end_protected
