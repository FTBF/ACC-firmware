// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:41 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NBZW7wAbOpdv+V4Eyu0oAQJ2GEK/NN0tiW2UTyOliCca08V5dRHmzk+6+TdjClZ4
MZIs3xe5coH+GHBN/oIskNW5CF25s38Tx9jT12VJ2wZryjUG0WplYeNRc9rG5lnH
WwZ0M6a9c5BRqz9AyHH44pcQux9SYPwAd7auRkw4KXU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22608)
UjxSJtepoHFNEY5TNACLTiPk/DJF/Agmd1KHZ5c34KDLH2iVVttwiaz97m54VHkQ
5m7bGtPcatNj5d7O/e0ZND2JTjdu7KafDA9Ejecx0LkKiR5bJwTos0l8wSOLhlAR
ExSyIrZpYaqME7m1Rgo+sWk3we9w9EBBvQ9wKqWKHFQIHLtDJwsYrENrLyS/nSIc
HZub2fYSv+HspBFvojhhJs0cSPrU6z18bYyt71AQf1ApjhrXIGtoxx3WG80mqLxp
KPq98I+mndBAgF5vO7AMVKmqDBgv0rT6jujLd6bJp5NJHtHWFU/zog4kxKzB5JD7
5cnPmQ/pf51L89AWkWrNs2fKTKiy9fAuPfjZC/N8/fs5tt5Red2iP27BCp8in9ZV
GSvLPJR7sh3bLRbqwEaMXAWWhLFWtCDiOWpgndALm3XhXHiOCKvCsZvfZ7aSVjm1
XYLXstPDx8/50gMK2dPws2rWG2yfWRMIywof6g719eUsahZpS1XQJDz5phvJACrw
q2zWjBLoZmtWN0anHDUKi2Z+x0R/r1nAw5r2N/iJ/qcPDxmoer2nDjaBTOyRYu/q
w3NNVBIE36zqI3scKnd9tUPEAPV4k1PuyoUVCnf64Wt3YYWEiu9MKhRa1Lmuz94D
rYvdaqPQY5VA/dlCcztC/9qBji8wbP8I5spw8p8aUrs0Ma+bcJ9v9eFylKz/LIL6
3S+GQ83W3Zsph6qLlSdZ2IBIrr3NhkbpXhS8Gv0LOlgba03CtR7ax59vUZbsqKzG
cUe2fFNBp2i0OIBVXUMvIUKOWxrp+9PfDt6EC7eN7l2xnganUu2XVywsU4zmNqne
CH2xPtHZd4rEdXKOlO3FDht4PWXTzMz4IyRaEgeQI7fbG88lwoHhpxNl8n4FN6SL
xCHS7sH2GwOwUvsHYT0KJRq9UUWAbLzSlZ/hEpY+hLhPBiA+RHiXVsJyW9L+BpXp
0BVH3NzeAAD9WDVokrqIcnhGNJy8qEr7M/D/zaBkAKHN7EDnDiKXLt/eLpZfwLsU
X/pqrcZZh7kx6u4opCGFsb3/HgR6ZfGX8BUkTkCaQ9QM29HS/STdraMbD/0aZxke
rElDGcHuFePkLDm0tjy0EBaXkkCENhRAJ6jyvRuowmVBePcvrbmaqZtJfSnx5w+6
hop0ZiWgik3XC8JjAGzjYC8tdOzU6DvEqj7XjlPWCqb5v9WRGSEvHXL/kTDCA327
fG9tf89gg0Uv1yBsu98FRzijeMO8/FfcQ4/Ffz7Vtr96+nHBnrUTXgwxYPx0Q2B9
xRYooueHSInyaU48YVOcnyJ9qFqisEQLNX/ch3SZT08zlfFQFLQNdcmsz7yjG1Et
aCsOBjbqn8zfd80NW+kz1CIsQcFvvac6kyz26MqWYCe7EK5He0Zxjrf5w8fdjXgn
eKRlkiHgq96I7wz7YQT+eNWCbT70tbgOodDJHwobvvmKQGRiWBm5V5neeyzdcRKP
Xg3Sd/NATICnlEQ+0w6l7Ds0P9I1tyZwxuAyexUxaib4JsVjAYUGvx9BOEH/lZ+z
S5CsLVNwdIDsOyVhPzpXpZN/DWN8tjVeqGa8zGTo7OPifLQnRc8rZv74lVCsjPU4
cIYC/oxqLi429LFczDoAvKOLBIc68akpMiO5+HdZOLyCr/eK5QzZKNvF4exY7/GF
LY3p3k7Zhopjx+rUSAsVEuXE8GJNU6vbnBvOE0B9ZJwMWCG1nbRuKWC6/1MFsgUj
01T27r9MJozaOqjpoB4auGAHWQMCNU3N3DepDRS7XwTnJbzPGLQ/r8TOtAMiK/q1
OH9t347kagk+lswvijfF89rr/nzATUWzazoiWdR3sK6+LV77rZrghPN5vPn4XonP
cxcty9epEG2+dRsXMJBC3/cYrPXm/gGJXHsWrbqj1huex2KBoa66wmWBv0fdE57s
tN7D8SESsYoylq/CveAXlI0X66yx/8E1fbasmfPVUB95IC5FLKwQll/jZBw9/cRX
cJCXUjeefWoRI1LybA4qA7hoWtlcTkRzK5hX9Jn6KloRZMp1SD947FWbJmuDml0v
iQVGzzGrw3NJgGeEbFs0rdBy99ZD503RJ51p1wr7ipwbgbFM2iLkS9V26B0TnJZt
xNjoXNpHIXW9mbL1AAGQPpWXH/b7ySppeUNK4Xr5MKdvA91b3iWPYo4DuEZBecX0
y2s7h+pLEGa+BtvHsiFOWoua3DsHLjAig56iFxDBnzelc0V8P3c2w81xkLn7hR3c
f2w5ZhyDDGvydxNq4t+exyYJ8RLukt+JTHjf3EgyLvSzhLj/kB2eNxYfuNVeZYJp
JM5qoRUIHUN2EBDvTKjJpUbSI0ahIGS4eWmL7DiBrYpQUxklDTMTpSyL5lkKUJ8U
fo+f5O6HAzfQvkoUUSM68jL2m0UmaUj2o3b7lyBbEHin9Z+feQ9w7uQVhTDlPFvj
ZROq/VV1jMWKZUpY0TGBSZVffc79791u3ZcQwV19yHdDBeLRwBMru09hlQEGrUVi
VB1JlpmUN6EZfSVh7iAiqiJmLSBUnJ4SmLyfRaFH2lPF69SRPFN6EJEuFSMdMR1B
+hEii8X/mgoEHXsTEHHagT4z9Lr4RD3VsiOrGwMNMhzGZDFOhJfkz3mkjiwH5NXD
b10nxwdAmcXjlFcjKB6RTnU25032jR2XTh6cKwtGE9QivzsP0HqxNhb2MvH3laOc
G2I+BYsimvb72LcsmeEYB60XGa9Jn6KyJjOvc+svqG30BmiB5uShk+g6Srixs1B9
NMJDp9e7Idp43ZL1wIJw/YFiL9sF3J3NuvvD22bt/eUMIGb+VXk3j+raOrUp/WEA
bvW8GJpJTdzTFl2jS7M06yihWUuNjjXgHkSDYZbQFE7czTbomg6L13CgddRdSH3J
AXMB3yMf51VB6Ve/dcQ9JNpc5JALq1+3KruzYagXxiWbUxSQ33qcPw6inw9msoSa
FZsiwLQloh1sWX8XBRKqYuBZyCkoKE3yxKBO4JRSs3BEnxwW4LGGQdIEj13iVkGH
uSCC7RxuWzi8Goeex/xVU8admtg1xvnTRwEdqCpoARsKkmLg6NQtqkBzWvfmCDRA
PmX9pgM8/acxbUZ5khzhtyveXAan4SBGrMdDrDrWS9tTBlpu4ABgo89qmoz8uSkD
MQ9ibhc3+Rhv0LDNYcit2uR17ttdBDW8lqyAS9Pcnn7i0z9EeKj9zOF5P/u6FZsu
soKcE5SViPrDY0QyRAIAOR/uP3iPabeQURPBwC3o6/MyuyasKjX5fQscyBBSnabz
cKhjivwy3E/17AWJFWQrK4a6qYA2V6bcnBBqj7Ml081u/v5klxG6FQMakXxidRyf
Y0dVmuAhLzi3eJd5FTSr4r9SkGqDQzZXO6IwiBbxfSu9zaTmyrzGzhlb0ny/u18p
V6Cyf/RbvU+u2M+0W6sxpagNP9npqgyTzW79eoR+PONJCY8C7pJD1Frpdj048N6A
04N/Ey64ohTekuNTfL6+OMa1Ie6da8sodn4EF4VEb0NGcHgHiAIgL2JeuGq/pfMV
olJD0rUz6LgUqGbEVyrm9RP4TO5b5RKqnnufkrbeoW2yan3sLMX5pRm3lOKcb7+A
P0/Ny5qkYXIK8rpeDlE6qZMyf57fn9X2gyv1Mi5/PHPvaYOl3CIhILNt0Tc1Pmkw
LRI/OKsKZmAFvWI6uT6qX+evEYpydXWubWlVyxFEkFRrm+LMqUgOKTkf+fWsuq2S
Ol8owW63Ej31va4tTqkDQO7qmwy5WqSIuRgLNP0jRmPUTgK5nEwXxKvIJAheQegD
lJqyJSAfG6WMQairVI1FI+slKa+XFM9+CYDAOWu2V3w8DS5wBxylcAByBYCOT9pY
NjhR3ClfKBuYjakdVLpq00fGwFtvgdc+RXqY4Ua3IMS/soEbyG1obkc3w8+Hv8KW
NuqI4XS+jNhaR9uzIaYxFlC28wIFNsAfRCJJdr0c3uA55511Vl7F2gGHp8RY2oAu
7BUR6R9PP48b2u+XNarDSdKc7og+Bgw/3eV8YwM/CrSbdGMwFblZMOmSAMIAjb5H
ysUjtb49kGEpsZJLJn7PLAWNru3bH/xYaNoTw6eJD0AYndQGkNArhxMxiBY2Ijlr
V+VuKssmeFT+q9t6MGi9Kom6qkzOKu/27gfllUGwOi1WTZtQvDebr2Hmz19dHp5H
Ai2lcpRWzFQdeofTwMwe2p4nBQ6KSBeFfxYSWyIhlCb6jh8We7xhJp3lDmJtwjKw
AxkLd+detKzOyq+LcI0XAM82MP8YVLa1rlAKBgEMy0Q0vXuAjyQCEgI/5F/+XsSB
CAkWORrbft8cUt730BivTnG61CZNBZ+2nbZv4+kzW+gcQEIouWX8lYNBZ+IpiKOo
hCodkjJ5s91TLT7O/5WVMDuBrZH+dpCwe/a2aSFinscPDQmCKw8abRXRTa4C61ER
Yiyjs8KzTg4yNTzM0ceppg4AbJm3CPuaGiFAkVK+HZ0oT2T0nVWj0poT6i5qSCmm
zUP5FB/jPiOuqw9Pi//He/9na3wjtum4K0jBFONjKiweT7gbxQNN2d3Sqd5792W/
DdH54z/Oh+NxrfeeD/OfUBi1+fBfbHBOPPD0cdn3YWGF++gbTO0RumxVTjvi8iPd
IiEjhSCFUP7II2KXhK7HBvr9kBOKWbu9GHwDMc6bAdENJk0SdMDx6KcpRR3JDU8g
sNQQv/IskAxr8iURibb3X1fczyZdqqA865alWP+6xX+kCSilLiJpmwf2bEURPgOc
CSfOo51RCVH7TxbgWw1liywBkgRUkqf69c0Xx0ciulGu0jar3/HmdHFTjlFulBE3
eOTUAmto2li81ccd8DuuzbFLDwwuLKqbT/NbN3xXVK/WEmXakKn4GnTSUawGx1jW
NeSN8s91k6jrCdL3tKM2p2NnsLJPEGlS1hSrZq+NlIddciOTiEoiplH2apK13kiw
i2FmZy4qt2r92DTL/dECNqi8bf3NBf9R8CWTVs9HGlG/tw55WZlYCimM3oSI6SMg
tu/RJRdyk6enBj+3qDbwzYxzJXr3FhDQqAlXUj9b6ksuLqNv/07T2EiURJr6sUXH
UuE2kguxhNvVAdHWKQS61/sQbqeOzpP7PKZaOlsbnZxpPQxl1c9k+uHzHrvb7ymq
R8F2jTxT0868PoTOD+IaXhrr2MUcK7iY0c7w2PO7SK8jIbt/ntVImZi9bythsDCj
psxyTi4tf1ICNWEs9h0radbDIhtrj0NyN8ELpDfY+ixJLN8KvFrawsJOElYn0AGn
IodNKUnyhBKgfllABuHhLlSt6wumXYhkSNMAopSFf66Z9zCyCIF8ZQKroYrobHFh
TxgXIJdfGG8Zx3NzJXWmGmVeDennNWCFKN4dwtvjoWQ8frvymuevhRzQ91SbUIur
vJQhkN/LlXxvypWvfigr1Om7wQs7BK3CaDwunV7ILfdSlbHwkZOKcCDpqwJPDit/
MvJx7wWjLNX1GHZvaS77hlPlhvPcNwWgInC8ZslOXZX3FbWwC4NSzCIXbHeFS3AJ
+RXPnbI8bdsee4vgD//bOWPWhd78MuOlpROFSkQWu48xuoMOQ/wb+7jd/p00Pu0u
eddnXuXjclf49v6hVp37LmioXfy1xLTTDsIF9sGtf3GEzlSgLP6xaEJfmHl6zrVC
14ONZ4BXVRJFclO6YBWBdjIKIc9guHSJ51rwCS6sApS3L4P8l8Ac4H7bFiEQT9FP
TRWr74HLbQmljFDFOwPT4LOBe6b6rTnGOcLQ3jnW/Y+YZhwMCOy+d0O8P/WdJinW
wqkrpAlm+hvjntHi0iaj5HKMLQEZ0R7NQW7GOuuTUf93uBUzxcl23+dfMOmvGBFc
3FOPdCO5lvOVmGUX6o3vrv77Y5fYo1+F4ZBAkBqJG3C36fhndUvwiD1DpPowWxaH
tdbIN/Y4hvaJmFAH0L/e0RkQpUlx708S2sSzOu9Rt5R4Osberoj63pLo7DqW40dM
QP393Ti82mjwFmOKHFMmNJy3giCKkTagn0uOQ5Tb2mly9SMoKFa7U4jKyFqyAIUo
QCXAhr0rDXEfnrz57umQrcXP/hazOCrfzBw+mbg9/1ZSWd5Qfr4XXPJxoxnXHdim
qsog+GwQeO3U558LLfrAsQXyyDBPDjqpJyx/h9ZZQSo2mALc5sGP35b30Nk24QAo
8eN1z9dXLExI56FZZNv3EZhnVZu/Giv4LzvbBWFRj1sAQNPdR9hwu+nmUJt6P07p
HuKUA/UcFku9iaw3kqcINWHoX1LheiCsXV5dq0tLZBkDNpqHrO1UWEdBeEaW04JT
Bf3eO/pXlAB2vH/A4Ypxp435KZt4n3y8bQjUCdnDEf+NpOajZ9gAVJxdbAgRO9Bb
fU+Y/OflTMTj3qZbwlF5eXzZMHi6xnarxbV+sgt4W07cp8knsuQ6Kie4jNnEwWUV
OAPlJ3Te5Tl71hnHYervShWkqa7sppIiuszqctFnzlp4umqppZg24RxeHmlOSo7/
TaDVMaOXwGNO+sdJlLqqa3Q2fmX/tktSI6jkhJB4Wvu6H/ZaZI984caqUsh/iJsc
NYSp+j5NYYI5vSb2uyuehnHbVn6G0pn6YbGInfsXBjukEEpenDANPW4X8kYqZzgV
+lZCU6KyiKxagrdlGiD/N7sPBgCWvT1ZbYwQpOnCgLLki+GU28wjrbcOHPuPa4s1
fTw8pWHDUnJREjRNDkfdpHikdDga4FvU8HFcVDAVVXy3j03lnSUbV0qsoQXmiqJm
UAnF9rKkzDBcllSv86SRq8Z1xlHRRo5fqyqMSrLTl9Eo9H6/Aq3keJBeBElbdZZP
yUBHCoycd5/YpHaUp/QU1zPGfB1CJXKJeqUD5gcf3L+I+vykdRuYRsZzIMjadiWS
zq+CtReebGwuO/HCzZQvtPT/hEl61meFjXAMCKHd4G4yNa9m3I8RRKdUnRg4gLNe
UFy+OvKPzPkXZ3ZsvG6VwF06YdEW9xX0/l545EeMIXdpqj+ixu9CoDXFAIKJtbsC
NUFbrzv9DHcLde1gN4nxICXUj9Pm4spBNO9v9LFyhmzgesb78UiHeOFzZF6CcrpO
Ch3glvZqrTnoe8ZtvdxuzLGLfzwRqUqw3egv7CSLYaT02JzR8fLlp7kEjGxNfoW/
OdO1cDIBdoblP6LLBbTJdgM6ngssw8kMuchji4AiG1E8IS+qhAH0cN73eFzt4J29
WluVtS/wvOyCrsUHHx0QwFzpxz7RpM1hJ1XTaYFnkJ8Q8cS0xNX2Y/zONWBIf7Vt
L2KjoWJ/5xHEsK8x87X0/oFuLWCp68eh9tkm5epeNumyByh0+9tRkhMK9nv0/Ahy
m8dGarBldpWIVJlb6lmx3eVyyfuMJRDKP4XLjwU4D6gWcjhQydPH9VgAz58DBjvQ
0u6lphJObPVXCwLLLaXIEBZv6WZx57LtX1TCy6Ocy523nU1VI8NQxKkY0y2Syj3C
v8stOTqphwrIDaa3rD9Aooe6BSshHOVj/lJptWvPWanITih97MguxXj8UrJjukTW
AJfH3kK8K3Y6+7xX81HsX733NE/tDFDTVOFoOtXapl+1KxYJQHZrS5WOAAmwA4OR
6EtwctQt+EQLDYqPJt1OfpQ1NnQ3tpNi+D5q80Mre3dlXc0JpVTv1WnmXpu7rgQI
5thDgBjFLGEh9PWFGQF5jyZ977ThxmELNKiYkR33W5AkuoaosiAAvD7Qo3ovkUEF
KyO8/pmwwwWU5a17G1GF6neaBwSkUW9KfPWTN4Wto1s+/LBTQCNaqUwHqBHzeJ4c
WO8/7F+KY+WlpS/Pm05jOuQkcsRKzo90ohUSEBt+wm2gu9VACYJYHYzQ2e6Zlv/M
A7kx5CwM5c2qK8e+ZT2VFjPWP6Dx8KG8xQD0NuKBxIC+KaX0GOg68sQyew8R+mxr
AyOoQ4P6IDIMayJrrHr4D+hT8cWcx/SJcLFI4brUX5SSqeyNQTvxqObprQQMm7Ez
7JkZNbaIqTggP1kd6ILFl4KwTVo/ozxcn9/3nFtHqYuT3PZUvZQbIqMo7KORXvQT
/SIcU14lW77fipXhZs9wBAOzdBNGSc2VaCtnyXgWvrb3ap6CeohpHJ4L5QA7Kvf8
6SPXnH65jgzYLmG9VAvcbB8vbfW6OmdODj1B7zvZ9tLZStmRf/623BeQ52yDpEYb
PpRxJl9UPK/RoBn/i+dh8b9/UZPf18cbiv92JBs41WB+4amm7pK0DvNIH6/4UpdF
m5wT8IzxqAzgLxgxw7yHgtVyYyjRrYbwKB2cppi2CvkZ0Wri7xtsd4jrRsYy1iEs
EdH1Ln3vtbLMsPUuumfBoDP6sw3IWIUl0A7ZfhWe3mUU0l13PhTKapNmy4AaPb8e
LXfmey8WoC0VfOOFe6MSoZM5pUsy0r7LAGLlKcMjjyBev1rXDCtFFnDZQjRejknZ
443eB4zjNckgeWzNHa1u6TvmNAInX8PvapHuDRS7JxEIppJKlDvWkwP6KYQHshOg
YpgutIqMvFRvXVU60CzReJi+eZRaNlmwRBVkR9AWS9bCdgXiXoehIqP/WMssf5m4
V7vNsM5Akq/o331lZq2UpXtfHc+uEwVtVXHwVctUg5RfainSAV77lRmFAeiEOeYh
xcNs4QszrTFmx9fv7Q/Gylju2UT4y0Binc5x3uPz1QnCRcvuBebUCCnEi0JdfhUP
ZV64C4RG6BvdEKPEypAASXZ65WEoP3hziwJTXz1BPz5QVSsDkIoRC3R7rHSWD7kL
vERP3eJpa+P6vxYNK6SqmWyUYdz8pZIxGv742NuQY0PPZHOfIi11tzIJ/pm1663y
jYsAXSG7zbxnJ1/rzI6uHBGN6rsOehicRtL43niQPQzbWCZuXqGlP9JJWoGChKFv
3Nnwkan8J9a/NTA1+aM7uX5Lds7VkMWJxHoC0yNWF7kEG3IRJHxANR2AZjMVAHgD
D9HPaSrNNyGm1zDK3LlurXZHi7R/IIcZEnbasn15os1NCAYdyaeFCLGjTnKKS42t
7+tCQWvjd8dD3OUvJTmqKO2SUL0xx7QMBBbnQkKoueVcGffxD5Rrc6c84bDF42ON
C6nM2T0apNmPDqmPWb5rKRhsWdDEzxFD1TMLrZrXNqcml9wXMduB1Nm1FD4XaSJo
dZpjTFTJKgJq1S1U1O/A4497U4dS6+nVTeaQ62LvVH8kIpptiP2nPcup2PEa3bGh
5GlIUUvka8XS6CE+HCmj7Pm4+ZqWNcQwlg+wZkVn4zSCoTqPMMKAVtVPqz7ErSnS
wTBJi4CJcBXk7j62ni2EfdzX2/zjVrUDwDiF3qdhWE8Dlx9LfWZH4pYXqyXs+OHA
Uf0KZ4FQVnTws+IuGJHu4Ai3nca+l0s5rXRPiohn0mZgESMnaPKH4ox4HWv2hopY
Slgp9O3BsWgV1hOgs957ZSc2S+nUlegtKE44nmyCk0dCUmE13h7UEYzxNPo8SP5F
31iLN2DBgCvObthqr4TGrw03JFfQSIM6PNxr7MJ32teXqYGtCk2EZ9TGhySnPy1r
cZ67vu8Wc74B5vnTj2lEKnamwNRXkMaZEgBPSfsIVKHHWpiCY+HeIMIYWRUyoWzr
kqwliAnNT9WhraYyZlVKmOwfOERvNDlR3TwP7PAD0VO7fM2lyqK6DQ4+rWRf5Ty4
sGqeovuK1o/28EC0AemIV8CgCYvGGfF7pXYh/Gv4jjA3A488kpQJPSggMp7wo2Xj
n4NlfqEpkBN9yaNPIFE4jORMiRHVxDiQd/24cN2vMXSLGGOlAsrIh/W9AYq7OLpW
RtO6/gB0WXnO0nfnw4ahoTSQtxZbFhd9E5QM+YwsybI3X8jAfhwSJ+tkyz0o5L39
b9LvvsG6LcSKkJ5U+qjGMFMCVdv4AFOhjZ2PikLlobN61/Y1ByhkxYdZVsHiKJRK
o3kiLEN96IrC9E4Kcyr6pMwxc+kc7Yyi9fECharia2HSJJehGGamGtiRDHTgqRzg
8Ks1wtlaOVE3Zt9Q+3nOYdqTliCnsuKA7cmuQEL6b302IWkGmEfYSAgyYDM1x0es
Y9w20kzc5WSY8wQxV3oHPyskXMIF4G8BCb2fzj+s1gBE+uJ0z1FuuKF49y0STVIb
BCXzB5lUXifXe/gGz8VA6v5fSplcP+XTEyluJGkeGJGf3Af7pYGnc1qUd50vUgiQ
BHDPGlUZyRp2nMxBe20s5okEfpq1K4WIho0vV0kDIaCHmsoD3lIpVSMSsYZJ0VHS
UrRb5WDtDM9tapY3oRbbtLOmF4Rsd9r1izQtOq44gLZNj1FYxMeGO3NkIx/N7cyM
YL7ylhmcVT9tRBCa06YxHG/3ev9Vlxbg4dxLiEQzGONSpScfAV7dpWiwWt7LPJ+M
7+SXNpXoDDzPsznrU0MJDKry/ogTdbzF38RgGb9iRli7zkAkUCbWIPSqQ0oAkb0+
l/lERPrgMSQug/P4cwPay9EZneN36Wxdh8Et/NIawYJYhIh7TLa/GwTtpxNpIMm6
OJo++te+7mNNuj6phC8FYOE9KRkU4Db1wI055TJN/OyrpIJWfXL6UD0CSckh1SpQ
3DQ2xR0JGm/JX7IfF5oIBgdJ3vrhJebMTlXHUIlBt472TDAvsrAND2vJgfLBntz1
lLFNDbQ2bqTspmWa3argI/KYmfTL3SIMsXGcMAOptl8T3EU+GCq133A0ex0S+Dwr
ng35btdGmqRZmLCsbOBHrhnjcvuvOz0hCoKhxc+LRbGctWM3MCSlqFMqJ2daN04w
Om9BJ0SSDicczpD4OdgcJcslVdCVaRHH0CAgWOY/VQY1wVejMbhxTff++Zp0tVzK
gHcPtOL8VjN/6ctVWa1GZCXwO2n9JMYGxt9kssUld6YGnn8aAoGWy0AHmn/0BSAE
bfqkYKcWGTC3pEt/X8mgxpRE0Xg67HCSWfllomPJe9t0xApkG7rHOu7XRm+FEX1G
ZjEUwJI8neKfuxGjr2gYgPSmZxAX71kwxbuAsGkuAQznzhoasWucr1lABxe9RNde
5Fky3SNIYHnkYOVBtDwoAVIYVOXa9xANxCJHQxdugCfIds8xoP0X4DWS5d4RCSGT
aQ+QMxO4L7I49OwaQekUfRKvhYY2imlRfM072MIgGn0dc4JHNO7e7QL30M6OnCVQ
7C29nuOxygMvjkd992SX0fx9h+4ur2Wvb/4ktJNqZWLczFDY5B4DmV6uM6260OH/
lBI3YrkVWdKLNMHCTv6XcnP2RuWEE8IEG7P9fpHz1yDeiYKuaaLSB7mcv35wrb1G
js8/9M/bdji7u9Ae9/Cw+Vx2q8SF4KrlsMJ3U6K5bZQDSsWDZtbgIW1ZtWvSgEjh
8TK033dp/m63ukDCZ9XqA32R6huFWD8oP2coUTnya9LTIKv0lb6M8FzWqhpTwcka
jWoDbt98E1sqPF+w+eBPeP0Bqr3/GB20axYHboo/0Xfh2rXpprxmsgEbQm82wDAV
5w87UhbaThlFbahIrK48yvG6+xXNnclDZI2kETUQEiAzUq4a4sGLQQVhuCnRjVNI
gqU6/wCWWjgRCDzZtpFotAuu3KN7lYyze5afsUCH62g07wi5AUXtiBcSdqJB61AR
S85KwATk9AbiGZXffC1bLqUiyVYaTv/7QlSo+98vrtNhn9slwsb5oEfY1a7E0ZRt
1Ed+2igqV4wK2Le0vxp2ewEvC1g0mOmQIZkU3GQgutXEqdOFQcefxgfB9urvZRPz
pvztXiYp+yQY+E8ztkAnEFFfc1XcDe7sTzIdbgubz5X9O/hFYY7lGMtJSnmujd9q
jwGmxNx7U9CGmZMZqMeB0lFIsyh1BmJH2KKWWkYtx1mA9ThE/1or6YSb21UEPEpF
fD3y6LzuGmR7Mz8hr3jr8VBsdsgfPjUvda8ZyL2vH39Ycr/CuMiQ9sxryr9EbNds
raULDyUEDzw6NxHDHZ83DOUQeicKKYKpqEHw9FVnlAGVBGqeMmTgl1WdkL3rJ3En
zR3XQlvE+5ByeFQYmhXfwxoBRjNSaF3GYC0gk2BRz41arZHN3iDjuN4ss2IY8eS4
72sDbEnJbFvfPUXUMzRukJV3RUUsJwBi5E/5gW328q8LlHvukeDZY0t+oX3ebgHY
6KoMyRD00tBMP8M5BDXxpmQGEVMeh62+ff6Q+jglfcKxtYGhUij7x04eBldXPKee
Yh2Fxq34uU2uxBm/6QX7ADayII1fUVWFfodT6lM7hakdsxhwePLMhJnIqJMjc1Q8
vnqWSqljVE2Pb06wJo8WQsBaM4rqNE8RpJ+25IDLoqiSQCGtISR0PJ49JKWyCAYB
7dmkTtMzgHWVhoYjWxV1RenidmAiWB/xiG2tgmVSenPkjoHlG1V7Oj97dWkN8Ba7
Kh+YQKs1AoP2w+8t20gO/UKBPytGowrABairOI/GJjYh8KIkN/Yry9E/7s/yGT30
7pNWXk940kg0jPzVzRQFUaiMtPG7qIm/mA8hb92IpNStsvV2u/oQYNpWp8O1sMJ3
9+Ez9EsjuKwyvcAIhf/JQllg3t2IpfW62hAEjGdHz95+YhHgVNVmI2Ce426uT4b5
CKRSg+g3LKf6BsXfk3YJ5PajuPGrXrgFSy74EASRY5dT8MaAKfiMbRUR5g873Q6H
HSk4J5sjC7WE2QaxD2nZy2xf+DHf5Jq2Opkb7Xi92IdBVvDcslc7iClNjHmrfqWH
QQ+vMCeDp/X6Dh4RZoWTp3UEhnPzis8/bP8OTKM5HG6OWTw9BVruIq2c20E5iknz
+sRjH5spQvKVGj4EPEYcgzUUO7IPgmi1Wgmlsr8itahgzsrufyntljD9pWFCMoVr
UzAHQxjbYDsSewu1WQcAtI8vkfFqA89CGAL3UCSMTFSTkL/m9QDg/4w881CicrJb
iKeZ6t9EAaTqyySJa+cqHnqo/fZUlU6MnwxayEDQKnIvWeyA5R+wgt2KQ7zU4GeV
YRtPXFc/R3zginx1s0HqDpPDksJm0ROTeTwnk+pLnp0c2+ZZpr577UzBr0leAQ8Q
GXJLYtFBp0wv1J3LRwKGMKIofSoYnay6OjLt0KUQlmTiWJ7cW0T5dagYZ7E5Ub+e
StYgMQIAQdU4HdQohhq0BEDQ8qbZE1hB4OSabKEg39hiEgIqhbmTNkBtdpNUA0ZG
AFNLaNie6IxDSQOinRwtNCnBjmzFkyi25mt50CoDETZdQcs7aP2jwCDMsEHrnkGo
2EQR2beoDURd41xtTrbYjvZJIvli3Txv4XsFXvkRsyunQx4koyZZ8x54Tj1pdiIy
GuBD1TK1YrNeuKEpdIuGFYIB2YDbvIf4Azn0bH9jpgOBhkvkfKmLZR4sAyXklEDK
9wu/GLA65jezgRqFF8bdOkl7J1r8YjCyRqkDXI2zt9KzgDZ9AaV6bA3CVfQF+uSM
9MmI8JLsEUKrAdWmTQg1Ry9YA/iE34RLZ2uWOswmgwfeYwOCvKW8AY3VF8wK3jM9
XMEdb+hnrcxRfO1Yi4fzRjkaqH5yh71WD3FjUI/Po3T43QZsq2WSbisrpvS0ovv3
CW7s8sqHeNBReprEjwEz/hboqZAIVgioPypADWEdKra3p1j9K2/9xpbaNDefkU1A
7JhLwhhdOhTvWnuR58L9wXadDtnTKbxJqBt43AYUFYDDHZWk6tNHdtLEUdePHtn0
8hbXrfQ+UnPDxslwAplL5qKFr6GtRYfPJqvwvtZG8CHt0hzvYrxw4CP5oJbChh8/
vCYi0xl06jJKpq8YZUZbcYgjBW3trapboO3YGVpJooiyMBreXaBbTL1suSW8c5De
C+BzATFKoAZE3dRAEWm/m2iJyU78UfZRN8qTZyl8VqVdx2pJm2/cg5YMy80iu2g3
2Wi4rQXLzAaKNkcUPFWWhZqiN0/dYb+G/+2/2FUi1SogvEu7rjoJfphCsE/3YTJv
9yRrsuyA7vfJJRDPwHfXleCc+o9dingsK/1ZL3YV9XRrOwwfQU0CMCxOBd2MS+So
2BI/Pn6T1i7Uouiu7PpS4OO/AvAVaNPxH/jAlruK4f1djA88gN/GHY2n2GjX3STI
d2pUvyJ8xYQD/Y73FaZ55kq29C/iL8n+zw0PXV6HPi1nzjVtAlfyyd2ie9JkQuZP
pyxygJCRumD+MojbPzIe8vlyW4O5aPrWB/KO3CWLEICMq1lJuVD1VzcdFpKb8cRr
xHCD7kgaSC1S2pEwmVovox+JZIYhzys910fu+pLIFX8u/ghMoTwXdy6ZA5V9xNpL
+a9nrh4TqCcfE+IwcG+ff5afDpt4VymS5tPts4S/30FWqueHyv3OjeYoEvP3d4EU
ln7uhqQnohvCbfR0SB4FPPpxDljYYBwDGnjwyIn2ozyWHVfOK6miECovGGXmB91O
wNWUIVDWqPBGQfoBABQQul+S97qmixQUzalXx0nSBZbfz24H/oAPR71g1G38+yQM
GxUB7SompIPKhpz5QE7W9q9nkxE5uvWrFZbHrvpXWD9Y99G8F+wJIe+rGOc2E9Bp
yS3rt5CAd3mmYIBL7cux5ibITW1cBbdT+Qmd8/slQPA6PlyMIJpE8P9ZQEzIVLv6
nsjN3BB5sGbXCMlc7zscV2Vqf6aRGVRSTcKIRS57PldPKZO1DMsEpuizxDhMMmUz
ww/fD1rkAXj+MLb1DxC2nsq7SVoPwZq2Hr8tdkV/BSCC7XSjhlhCyegJ4aQYZiZ/
2/2hW0qayHTAjOuyOcG5bUxic9a7jbyTazV9YUze+C8v3ydLTUO7gnwDMTxb+QsQ
GcTOi1DUHh6JMJgXlJkoRhTWyGMTUC0dpN5MbjJeoP9gguKRBE+gkeCw0qEVd6Fo
CtZw1wtHqvVbiit8X3dodogX8BfCBoq1WyzvUYkic2v0gxsZlswbU7mavV1OCv86
q07KZncEXJIGa6Kj2ocKRCr4xfKy8c1bNf+6ut5t914Lht92QrlIdMgqGeE00ytp
MCJlXLCt+ZLMipr5jkB49vZlkfgi6VCrUuhk5f4ARY7bEVY2zWli1nyIJ17qHh3C
vd9ZjoAUK/w6uPeU5lLAZLRyX9IXqqRtFMOwvTz9oBw9Um09BCSXD2TO7vAfE2ij
jy6mqnYocyqUok5Du227AnyJPioXUkDyWq5DCnjTxqrknCtHj3N8CwJlAOcesmte
Yc7Hm8puHFjEBMZtj6qWJ7HJ0tqxr5CuGzVhF89DTAuEEqvSRT/1H10B5970R1Ww
kiCfPW0fb80qe9vIvAZCJXylC5Lk1hjvDCAh8u6Yy02kSStQfn3j0eHsOhDZ/k8w
UUSnI4H9UYkneOZ9CVrFaRFLcca3upaOZgGjruZ/qCZQV+VgKzXPmxH4gRkd3DSr
7HMy88YZjCqyiBYn/b9MTJCtBZ362K8VNJdPwGWp+b+4k0wb5XtkE5aukqRLv4zD
GklD+cvjsot0crAMOn5nOTJmEuGf0RyTPDh2l8uXfwu7uieqsMTGvjp/NmrM10I3
vF7oJR42FWe3UsqbB7SL6cRezgAYZPFxNLV2MEbX6Dn0B2gycQr8zxM7regmyNm8
Sy/pbyLavYTm/GpoueLzOpCepNNKZ56QxImcHsBa6WO6816/RR5UZ+EgpYWXes3y
ZCr5KWHfJk1Kdtl7ecZR9zdf3c6rnUl/sQdN9fuuV5GK6TjSgfhp2MeaXN7SXmAu
q2hz/c88xgNhrkIm/6Ge1EFDA+JqPcR3dYyMp7uKzFK2DlKgZBCdc80q9wPYkJ+t
F9aJA526K6qw7ZRviD8SWBZ3fmiYubLZf3OoWfft/9qvjZbpC6uOj3k1FbkWUc7h
Std948UPo10TfNWRgMyUvdVb7tgxazITJC9ePuLK2KXLEgvq6QGHA3+Ya7Er2+j7
HKpdlkeHSCgYUYmR1WKGSF5HXcg7cGDF4MCPYuoxgQHczdiyBnGEVwQ8WwjnRUpj
NulxyA2bllg207L0nXzCiUxmyY/lAoX3lnEf0PaGZDcWaQtMIGQhlMEI25TaPpbk
M6Ds/NBE3xMZARHLG7Qxjl5ZxVuHtOze2kqXUfpan7Z19UXokUkj4dcSZKmhoo99
nwxtO9m+CjslN++LvIuWoxwjsqxJG8fxEng3YDukkHM6lMonnb/tAPvfTDIdjmh6
R4D/7rrsymecsOT7oBED+y5/OIzQTlE0Auvf1DYFzza+K/UoChRQecqSkeNXPbN9
OlKVDBVtHuF7M2Tv/PxzbZubHPKqMWVlIxTupZEn+1xeSoAVNW2038c2BOLHuXwJ
B6kYpCIt4PdRG0E5Si0lDTm6KA7S6nikWXUCz6mp/TPmWLoPZjkHTwi5QnQwPA86
RnTFplBDwOjUeh9HV+QBXFdFwfoIp/WpKBTY2fL+QN9Hk5udfURUwtyVUuDcinAI
e5KEG6kMRuk0JDvJUP4xpg5sp5axP4ieyGyrQvD5rbTqLq0ZunDlLuvpCJvQOZGJ
tQqK36RiYJMsB7rUge1Dr1K1k1CfecE/TrQtcaLGP7yOfagx5RNIoYFyXedTTrVn
FBdTINgHGzYTDAfKpXZY2H/ujx18iZjvcNhIBZV5aySxZA4iIR9SLoOlc4DP6W49
5VDnHIaXVbdgAKm+ljVoqZf+cqM644qLn7GQUP2fe7QvkoCxterRZbHoXJVxy0Or
cMq+lOh/c3SXXv/J+C/2FHQDntfUEzjjqu3Ce/UVOT/Q523zuoEUCxcItaAGCi5+
SLFFWVtlW48uwGNdC7pnrM/0fhIvNuHdZo3Brw7YDzL1q3/xC46TSllvBKjaa3Pu
ZQJeknFH1+cu2HbDi1a9SBifQxtbUAQ13hP+UBiA+0gMevjjpDu9x7tdv/x/xJ+y
MtPYmeQFxNSz2M4Q8v8heOfdIZAVpTE5I2P/4UrgO9SQ77FYQQrnPx3nuNnMlgI3
103yYaE4yiSdrrCnIKhSANjxkAGYrp4rG0YUhdj2WbSyMK7bbxqnG1Eh7UCNthvJ
hyVL1+rMtfY+9g8DN+L4so7m5gZYCh2Tv+FFAPVorrHFV4dX5J2JCzsNi0ux/yHY
/75hjokqgERYAxth3t2IyJWKaXuybfx/EXGyw0ShfM6icHgfm2KAUEjadDhS2FGF
PJqmPeKXfekt4WzE6rr3VKGSN+k+y/GVRLYbb6n0YD3nC8PKsGH5Bu09yA6+oOwA
1SlVF1MmcVnGrOVu4tNS1k+GjWS1SyEA9H/cL0Ee7WGfylvBpinxRg9Ugr19tGSk
ZppdUdyOPRBojfRDsBzzb3GDtm/enN1o0v09N+iLlGqvuhGUiZhigwuGuKm5EvlZ
vLjIsUnW8jfZ2QCMCDXaYEHKQm7e/HB3kyR5fxaDkbXYsyiADsjVv9mkMAKANbXE
+mCeLFxtaU0qlQ4G0zPWr+z0pBKNLCK18leFK7lVctQqBV+7dghvYtJmY0dXIkhv
oGCH+4lf7H11D3oFvEmhM4oGu+xP2eOd5yYC2Z/ABtx+nR2qgq1q+QppKiIEzfIY
8LYvJst9gZfR61NXYt+CgleYM0KOSB5lh2cJkaAmGx9w3Xohwp2tcWK1zNjzOzD9
MUOmyEEELz/htDfUvJN49T728taAsIxyxQZbt7c+0jHg+Xp1hvyouOUTl4BbtRRX
PExs7I8XdMK++fxu0HFKsNkPawonowZGqnJlT9oVmLsR+yYSNY+XeeItGptOWfjx
+gJ0UHxo4qa867QeKjTDVQzhfKHHGJ0JD/6UsAAHieL9Oo5tb4ZKai4HuvB2vrzb
cgBJuH20dhxN6/JN0BooplDpMwRFitUSo4X+m8CTAqb+kTPmYBxnnTwqQWICS3lG
fFKXX1OZAbyYLHbTOosZ+Jh3lAEOqsE6vkQYq1FBtmpm+Qs7yvcW3LoQkGLCWkN6
fZfp1lQpSjvaRdJv4uf62zA5/ZnrJX7MH8iDNQ8oJAoBEo8JrZfBzfzkpZ2EwgMF
iAm0u36sxFCZ3I0edZGGFJ7h0agrfA9zSQxkcCGsZFhySmRqugbOYdK+Mr7+vV0M
JaCIyxkefb+k21Epyf5zBZ0QrakE+PaM4+CZ6JcYyymvUlIfjNfYG2G31IqIPfUi
YX4YA88x4Gwg5uXkXUvzdpS/H9BSuxDNEsI9Aj1iqhZSs3XgeFPms8j+IQH4JA5W
x3mVjYRlNV6MoGToG1jIbqWS6TFj4qBc2vQjJyaIBVFl+hDJBHtER9V1O/fkickH
kl0uJ4Fmx0HNqT5gS7S8fucTo52SFksMbPnEpoO1jlSAePwZI4RuhQAK31E2dOZI
Qo83efO2AdSoInQq6pawiJY7+gBm90gho1VjjPXIIKya3VbOSA9idYd4975+PCX0
DKj7AKvnHMOBc0Apo42B98TRY9jN+3fvCJeWMJ/YEab4uFjhWmVGRUeBncdQ0zXZ
Ioliltx8II9rtzqDvnfqzvJRaB0V5qAxocIXiqCs22K+NjqZ5U0W4JNHRsSPbndd
7LSYIMxNhTjdceNXlmD3dU0KLwRBRuPuHFfHl3IgtT6Bth3Gb90tc7JZOqxD8PP0
HIf35uTZOhOA6M6ROkYpqcnfDl4l2w8qJGOFNbLIgJWZhHKXLde35J9Gyggn9t8M
IGqxbRLUNx/V2aqDSAunGWkvhVLlYj3mvz780WeNXSxEGz/UH+c9P8d1FwgQQEC1
nZWbYPoAum0RC7QCgxqqatDcJF3VwlbcS+wYJT+A2vjfvOoYWUdTE1bcOn+iVfL+
Uk+HcjyltAwUVxRQZ+E9Gf0hMdRD4C6KfKKzNOt6Bkg+ujfyjfu3e6ltEbehG0Gl
juF43fswM/j9ysXrl/FgUfMlt/JPI3f1yMT/BDWx87ZoQI8HMTrfRo0OqDpM309w
BHC70o8TeXtgL4jRtgFEu6inmHPMdsO3waFWgb3D1X+PsJ+NZXL7NNb8DqnPIBbK
Re+Aat7zITZRdT9MaDireCtdMdI/xh8cYjOLGPHT0sQIVDtJTKNgM5y93gRDm7aI
8Gr4a88LekZQQg2MZl7dWJDbdlKiUvCrj7lt+zhRrmVm0QX8AbdXUbrWo1brIeLs
frFOUvwwZT6x0z0yyO6wdDC1qfjFZBalh0+s1IIDQL6rlG6C4FgoFtJ0POLbvgtM
HjBv+lEahBhQgdp5gCvIPX8IArdO7lUZXAENYJJ3mlfdXISzu6HJyo9lbGsSnHmh
MsM0UG/YOh8zEW1g9hN8pUVxqzGM5VHvaEtuFGPfeYpQJWJh0IbwOp/5OjbpHzZS
WgoMBdiIKd0zQwVHqSyS92PGb9hvkgBFMVkrtQjwgB6aD/yTn3+SwNlRKCV5p8ru
jO68+NE85Xudo3Lrym/DVu11eu/o0HL3gBqLTBCUTsqG9vwoGXGaDrmH0Jk7qm3w
py8S2AYi54qCCYAKeG4HoY++I6XNPAzf0G/ZBQMcWFgxJMlfMf46pxG5OtpzjurT
mVeGmSeIsHNi1KuXXRVpCqU/q9Gmc1T3qPkKwfMMGuYIbxLfT3abtALnMA677UNc
R7HepOglFN8reAyJFlETq+oQPaA5BKbB7tfA+yvYZnhnq7eoSBD8YZy3cOdoA1gg
MbXTIlF+fcGrgBANtHCMRlMWzykiHbrvBtqSlIPOCNJYaW69/vdbb1od24f4aAS0
FDG7etisD3z1ZLe9T+JtNFm1bPnAYrqDrwRgUqYbW4sY2p0rt7U4sSYbD7hjwboa
g2VUqDhxo6Kn7L9M4yv+jcqw57agucFeZ4cyY1mphof9OvzygP0Mgvs+lD/IgywY
/D5vlU9NDELer7Lsq9GGr7i5tY4LzTiGnNntH6/GNoAEJc/R7UPCGdH/nfSUaN5q
ehjcRZXaqlk9m7JgMi6aAfYxJOVfmVsKJ8pOjZpbImS5kRg4WeZOFQPVsh1rkk0k
It+nG37qDk/WoqEvaH+nWBYCxWILFVO3upbM5YrWhbjeqAACKS119IjbyaHA+RyM
rI9Tp0xKxrAyOIY6Z84lcdUmpTX3y+J33hBQDXiknILka+/Hk/IvFgl6O1CYRCpx
VduhYbQ/Fahg8zqcQEvhlLX08fuh/XYtYPBzc7n5DFQ3fB5Nakirqcq2wDlLusmr
3x354u9TrrrG27TEDc2hBNIhM2mx/uQ/Ker7oq6zE2/Oy7giJ66GpHVImPSnfIy2
O1+WsKQr2vW+fnCba7k/HAN9zqiu5a7/ZvgGzchJtCNlLYhNdA4Kneevs+w8GvKn
0FgzfJZYYFojclmhVFLO3wngXbkAZJcZUuszQ8xdAQnk+ZZZqggZ0sJ/+Y58dv07
r5KImzZLDvjSJl9FNW/ytclXf9tCFbJgUFONwd75DkMY8yodSvp0eWXK2o8Fss/t
4+Kv8DCm4g4xPTLplkenyym0CpZEUpfvmK/OYp2sqBOiNjQG+j0o9doxEyczm+nY
bWgHgthsC4ReT0CIPhqWkUXqzRxmt9Ud94OZwcFi4MewrTNhi+CGfmC7HK3ZuJh3
HzpGz89A5VIdWunwieEbgvRN17GRDyMFHAIzufCwsqiXwcEmiDgc828JaHiPSLfn
hEdni7swshy/epJGC21iolJkEPWlC3qbeLgOJT8dvlk24s0TDAw7YK60yUaOZ7zf
lKVDkoqsdkvjUPRlJ4VLekGvoFywRXmWhsnqwx8i4ME8Txbv2afng/N8qdw7WzhO
hbi/6ZQhYbq3vpvgKkDPWCPUwgxkCmOfhJWIvdfHuu6iRkJCYxCJK7IIjvZDWLbV
j6helBU/DS2r2k093Gu21IashyDWlGVso+P0VKWWA73HureRg0iGK1nuKxovtm+y
dlbS3loDR4/DUK9Y+rbLhNWu7WL380RmBcpuH9KoSeQn4x6Ywkhkojgm5n9B/Q6K
9XYcKDzevWkvyCTWIOVs9oGtdE3gHllu03srxMlKwQqy4403HP3RgkLYDi8J23Rj
5atGxRdn8xQr/4X+tx+70DxM6Egw37fCdqXb9MTDgZvm2kANonFvs6Z/ZusKzgag
aSst2kgqFLyHfnbd+vowprbRPo8hofkosE6ToUFv0c44rg3ts7RX4hVs/DBwBmw+
WYdXsAlN4tIrghRq2AxH51nXoeva3Onbf9qM/Q0OC9FDXRtuo7YPjhArIPXTOxcE
6OsNh8Ya87PKfm8PHnjDPJwuP5s3pmO7ix6xr3c4DGad4IqB3JA0djytXTd37JWn
TcvLwq06bqkNdTpFd6Zp0BmyH1P39u+K/6md759ffOf+FitQHkwy6Nc7nktFbbpY
30jvBg6u5e9on4M/K90qk0ypNvAIP7tR14WDXezVpVn3x3KlK3n0T+IJjR/JDYpt
2r6hYXD91Z+shupbRI4pSt0ygVmEpw1/T3ebMPlTMx3bB2C7esUi4PKn9kS8G0VW
k/Ec79NmBPdqAtLONK8CszwV9ISE5Nz+iinvJK8zZMCc/1QfvTka/3QXuwTbUFQE
nQCRR8wpsczdDXLdMs5l6RN/RyNCgWIlfjW/cvzdeValqxaWkVG4q/mzPwujlHhF
ywDTzxzMQnuU0lBhFz6MxSWlpOnLhSEBTb1//3F6y3HxZZTLc+HwLdFLUC/tdlVr
C3+sm9CVawR5jcuriQb7f+D52avfSv1EVQiTBsriP024L/j5Dv09z+R+AuUiSzAY
cwkmA6AvCHC287u4tHBvfre9fXogHGdqNShJXgeDL5JGM5RUMz2fBy0uCvbiAj3T
G+z0l/HwPM4vqmYE7fSU78/V5FjOyaxSo3GpROFeBBNLBe3aCKybPC5LVWRTSLOt
g8/Lezn2a4RDJ9mZjjTASN5AUS4ctPYqZOS21kwUwB0O9AS4BYJj//bwT0eZgQL1
12saZC/LGUrToLswSfsVuOukacRdXeMTScEVQFNrTZvOUU7nbxgmYHPmSYNabrsQ
rtMFobvBrjeZX7uK5pxQu9DBb6lJsXK4pjovtcJFGC14P4JOBT0kie13vXvEnTuz
+RbfkjmeiHRH7q6WfBj8HU5fPwG6iKahMy7MypYPwBGo+cwc7JlyFg3gcUwZWHKK
lXtmXEQYUQrLVlbYXo5cCGA/Qx6E+/TObHhkMy/oYOOOT9r2iQN9V1vQ1yWlAaxi
8VBPQ0JzRzNkBgnODl12sX9AbuiJPbcmkWB5hrkTFEzKnPgeMFpzHPXXfQ081KXE
5Jat8V7uw0sqPouGv1iLuwdRJEo3F84/Md0k3voOHbWIZ7U5lQfSAOKADDqNUwik
bpE/YAMwTsumOVjfb2efXol0/Z5BMC1xWG0o9X4e7TnfoHdRSdORDltgvLY+QFlB
WxU4uBlwFNYyCTCN88MW4H1t92oGogEvoQUhckZTKif4WlOcqXVaRW68M0GAm9Di
hpvQr07VQj0f2vOvWa/9G/kevxlloCd36NDlPTp1xZsOs6d5sDvV4x7Ow9UyMRFd
7eqG/sGm9pKV0BFWFSG0QB2x4d35nuXp6wa1/38vGi150hgCUUQTxiWIc9bZlhyj
ZK2SdfnEYE+zniH+pbyd1bZYr9A3aYYabME/MREkdxzwwARUleJWVN6+FDapaJK8
wnSsaVD8kwvwrteJVfa9fN3e2AkKdaehCbHEHnToIlqOTMnuRLgqAJPPgAT224bU
eDtHSUSP+a41YF6XhrothgjF5mCmQJnZsn8G0+uBXmzGukHg30oyTLVrZ1IKO3mI
rKmH4cPvtQQVZR4ehBu44Vf2xMWCVeCQxXPQHnaJkkrmoP6W3EdH2zw0EuT6x3TU
fn6+lRAtJcwo5Uv25J3SCJ19DFf/R9qDmWL0IK2dcnFhoGv2BUSed5y1SFPB61ZN
1LDG4j6CjBRbp2MYxJPXGM/Qbhd+0eMj6zImqNQSwYiPK82dH1pdfXDyd1ym6l6V
VuyLWBesUu8RCm2xWNqYfpdjvTEu9Nhc/VCjU6oTAEdL+94OA9z5L9vdlwqml9eu
XOuyKZV5ZGYR3TGTVdv1VGqTAGbDaoLdUoAwl4oRsmpd3TOU7W5GkgesmLe3C1Zp
8Ta5fkBKgowAMLPjx+cQBkKrS7U22+yX4/NhEUHNIkHrT7t+/8qFeAs0PBcrXzUr
ClXyk8bl6cfVp26Ref1G9ZmZpvYSQb8IAswueAxFYqYZ1ogwKjOL+36ULcukndfq
gkrt2HLf571BOUtaHgXYgp42yXOTRw6gaCHpV7hg8ssv40cNVpjvD9Y6XY9zxFRu
Y0VCyVJbjyV0EpBL6NuYGaCBNC1f1kKnNBbdnujZs6YB5ux+wTJl2cqPkuEaZyox
X6pzv7jG21ldNfLleyqit0BNCalzgP+9uTJvdWOcGzgx95uMlZgA6GoJeoRamJEp
yGPODwG4btWRNidU0sk3KrQ7WMRxhbi9lfx63Zn83ZoBzr/xEer3xdDVg0zfoFeW
B+hR6qa9mZ9vksl+e4OxeR54UH2VIgLlMWDuXp7FGD3rhJtsJneVWSav5mU+pLM8
xaRRn0/8QDFHvvUJ+KZcTbXpDQMp6YwxhMPNtDPXALecvitGsU0QCcPjOsK2VEAp
rL9/ZAl25QjbWeDuxNFhLMPglZE5eeVmVfrrMyr0knt8N+RFz4HAiEnsZtG+JlL7
M4MCDwl4EQZ13fwLY37C0xFetnEc/v8UVPCp5pn1Kt5TvIvuRqRP+p5Ns4IgjZDH
74pS+aBArOevBA4mIWChEn/86zFULa5fK82oD/gRYgibhYU8id8FTDa+w3XZF8HU
5cPgvXHEfXfv9M7w0uyJR0GnWynio5gOCYn4IuDhdDci9NXsrQMfTuY7P+HlJXH1
/vueo68ALpih2kPK/FfynKJcdSsAk4up9D5x1QqUat+xyqJYED/tcJPVoFt3e0EI
LehfdBOge3oFD3NIBQOUi8j5KBV1lxnCEX7xmWvr+uOFddLTBAAyzAFrPMX3T1Hz
fKio2MTup2M5hNKZwd4g9oBThfP0TJfHNTnFu6wyEBLl61YZcgGsEKo+hL24n/HP
dSxxdZ5v7UQX4MF5VKr0P+a5Sn4DUTUsx5wUm4RVHsBj/c4N+qVKAjZkYDzDRR6P
M8Wjtb6mKlvA4jtleNGg+2a8dG2Gu0whd4QeICaxiJwikLYndRGcLkBhEyNwbB8v
8SeROepDa7APCGWnsQIJlfkq6nZzZvnKMqOgrVniwMd8vuLdQzWOq88pPtdbVugT
C3Y9QhyQorSQeBjRTAl30ApRJeHumwqtwO4qU2T4ygglGzvPVQU6HhLHwpnkRJ4h
bxOkUuQqmI2ElLuE2UHLHiuGXAnZDxoc/PHH0N4CxwK4LqAqA9wcVhPLwKy5RV4k
jSiqw9PDoywnoKFsezhSTAWEr7Wj+DyQqlLoAKkqmT9F1G8ZjFYiIA6uAbk/BXuk
76UzoOMyA5GNtXy4vlWb7+F+VsxoJXTslZWmktHvMnOM+bEaPk/pNOYkQZbTg9I9
agJfQIvJLcKAxkDVdtMZstr+DtI1tldHVtTw1HbHVb+uN3D02ShuZM278kiz9FWe
EJg9+gl0TmzfKzPpBeYZGG0Pb7UB3nNnt5eDUI5xs67woaQrBu66m62nQGBB6dbU
0Bvuyyb0wk8X4XIPRfsVj3SbGjwj/Mkr4s5coQ74e53dIaA3opjLZLug9tuLrJav
2R4MONxgCwt7kM1hzgYdaZ3Cttdie/HVLbLOB8vwVtfVW1uZchBhNdOOMFT65Usd
b5HLXt6H1dkyr8xA7yTu1qBkCg5HPzcQzOHgn2s5j94HQtrj4SlJO3MGTzu/ZMFw
1rsXAW5S/aeEHNfPPGnlP+KVr3JVLHGWPFcXhxVKcytptMei3vFRAb0N4kOyv6Z7
QO7cAsusPaKn7ILDrbLDav7YmCwIzMlMFB67FPavCnCt6V1C8r4WVTB+R4WzxniB
GTh14AlRcrfa7H6hiixNrcvdZcAE48RwvZZFF5Vl3D55HL4De1S1SCzrKCrDf+vH
XYP/ZTRuJCmQCGsKWOyEW/kMAAk0yYPkpseDYTrbAjxu+QnqbJgyAzafvK3owcO/
28lhMDzJLiZbOWAhSBQOQUXYxuoAbzyebp8WCweA/9vQMNawl9W05Dcu3dpaYqir
mNgUcn0aYOSSltZCAIv2awBk4PYfjs413Ol8y9NEzlSCBSiFS8rZsn2r/xx4AQZq
+NiGTh/b91V/LThOmJ7YqjynKYLm3ayDEjNznCtdYMq/biYcScywpWhEY9Ub/Fwm
3r5qOQZJxj+qbEnAEtOXWd5NFFbyVX2LmxnigKG6X2usLgsFS82lC9+/SqngpaGg
si9tbjnFRbErFgkkRGnKrZS7Htf8OCAuw0oyfY/hNVNZ6FTt1JBqF6tZieY4mLFH
FI6pgQLAaI8L5H57huA0rXp2y6pczXwIAEZxfV1PbhF80AU+41/L0UgJ0gmaL1dr
e+rfOmtKh7+gw/2jNs06cmMDrq6hI6Mf/I7oF6g/8uSVMjyWXRW+3a+AXPuGOAtb
vuGI0GxrvDzOqWMFk/DMLSc3BiQ4siKpU9FZWUCsJ+f3ty9dkdLlR0qPIoV0Gp9D
IkZFe4/llqrBe2p+pgdmIfGmlCj7U228Xvbj/s/Ri1+THmZkzyOnaIsd5qT43iIn
Z8m5xLA8VbHYsXZqEfCkG9dB5Ezo1u09bNLlXCCshbwGyNlS7Xoke+/eOqBhFyGq
38I35Nd3I76pHT0OYGKbd/ranoIU6JRJL46EdldOJawnTWOFCX+B1SjtxLm9DFMV
QqdhnsOem4hY3+VWnG6o0A9aitzId8thpznjvvvFLnyObaZ3vvx9u8poRNlgGwTE
v6Mdjsmu4YLBooX6bjFbx6CeAiBhYjnmQXuEkRP5ETp4+zpsyJUuJfRGTv2mzEy8
nKk7WXo+l9IoUq3KcMdwkISNrPHz8v9fmL3Nz5COyHcSaus1QP0k5dbho3v81L5X
Z5uJwlHNl8LQ0xX5s17Cp0w/1C7zRDKDO3gKfbhKgC+VFpMo+2WmTguSCkJ9YO5d
CVv8QzRVyRjIFnHYXI/EhcKRRH3CIWMy7jyGelYoAjLoO5ksN5fz1tr8L08Ync9Y
QhYixPpo3Olp8XhDfuE+01X4/YvSaF37HLQB4gcSwUG+N/EcozKSh53Vn3sNZjnE
0kk2NY+Jc4WXTmdbeoovc7qGrIBgrVbCd9e9munFgCw1Tqa+Yv+4bqXAA3rlzxpd
itCufmnCBCqIOIUiteK8IczLOGi7+R4VoBwoP5sOlPyBpW/cj//4wt5t9MJd17CB
6AeRAD02seS2rZYcgyghwYzFEZn0dcooHJnJVZXTkQYP64iXnpGPehdnMZI2oHeW
0mBbKRLmeW3cj3A2e2pnoCdxMyGW8DBYJwOly5/F4WBeRdLwFMBzZpA9+a9GYGTs
1xpnem750U3r2w+sgVyAErq32wa3ORvXfT7OAWjpYuCc3CVBQzMpNtd/UndXZU1a
7mA8DWGo7zABSQy8QV3sBqFEVekzuBqIStS+CrYsDiwq/ZDrxj4nKd0v8h8OesoK
f/73aER543hDYLQN+d8uOiM6Y6ZGqf+bl3YCz81B8HCrTV9/WHTcJdYv05XvkWxw
r95MwaYtvqbcQAVz/ewijp2nz+RdgDyw20PBgz8yfhsa2piGseT/BzrWX8iSTEAt
BvhrHo82snvwq5thRSU8uqUUK2G4G14T4kBsylLLF81glVWeIgYu24ByC84B/ZKd
nUYfrFKZpEIAaOtliqYImeNh6y8fCdtRmVPRE4LQ2mp8io/2emTr/3j3ngyi5rsP
6B+NiDdt1rbnc0vcUGunokqEckkb5t8YZIo4F6n5MweTwzWtfIIuAcLHq3aFAioc
xh9toeS6PummvnDmeGBdMNnMiuK0aVHl4kF4K8X/rQOZVOK2mpeqft4pmHQAGONW
JZYzvbzgicub4gkaOZeR+i88dQHOShKu6yplFvphkBBqKcywCXt4iAsQNZPRcEn9
htBr/uvSi7zHF0MwOF9pQ+c4dPqpFza/rJEPtAE6GQuxc5lNW3ujIm05ZEVD5flP
2vU1MW6OKVe4n264WLoN5obNB6cRZ6E4/6UCG/iZInN0EFOJ7QQZZe3Bg2pY+7L9
j7+0nGJ+LbkouucX1KOlTkB9m1rYNkrh46LHcH0rSDq6AI3i2pOFw6EpWPL+1VmS
FYsBwgR//ngsU4qSjyZSfqqot6XeHR15E7ObfJR5t8vEXqDWp9U7qYbit2v5eh2k
LLondHOcj/ZwoGyQSyL6fW1izBpNNIM0UMgR4tiojHW0uYXrXtlCbHXt8998nBZ7
Zi/v1BJFr649wGj7nijsXPAHPLa9gl/Ea0Ag1bwtwlUXygpkG/EgMYNMFe1/gq1t
hfNvNP+7aSHv/OzYFaSNS/yQUjGWOvCWTBava7Wj2YnFEmGYn4csqHp2vcjdIbRg
KPLDBfJZyme9pAz2rjECxjui0llS2SUEt6mm2HWFEDQTgq+k/uWDMu3W5NuAk+Wg
FFXJ8XVLzTvjyCkMmYhyIlSqXB9/A4753NjWcIN6ozKdYypILFRcvv/QfxNbFyEG
pCg1qYqkNjZrvwooNp0v40Ukc2J91HnGAz/J1QHrZdsTE68oMxZfMG4gSH2jiK73
Zen6Ngqkw41PE/OKG4p7C04TuD0lqa/tWJ5u/SyuSdbIXGOI4w4SOg4JJHyGcOvS
MY/yoOZt/LTUariGwtp+bzt6ErXhLMTttS/exgHciFx2IK46uvBzh99lXNa6HQkR
Hu5qm9f04cZDYA4Fn1PHTAbbpoL3WT98jpZmdtv0wcDWfUX9GzSDlRvkq8VVBqh9
9jSJz2CYvxMQBE3G+zrgD4t4tyGZRLWPF8wAk8HHb7jIrooLze4GLNqkPVdKwjn8
q50K6LAPU746NCLP4yMm+7lH0TJ1blukAsLoGp/H22JWZK/HckBGHfm+W6mKl/tJ
W4t7Gcn0bj6NGHUj1fOYLqjOhygqD5Ztk2soaUKOwo+lkNqrpevwdg/KQvfpxVrX
ZLdVWOD25xZE+XVKwBhu8olvaI56n0ShXhWoS0z9vg2NUnAdbCAsmWzLFuTOdhb5
O023gwHMsc4oQm8rkmngCk8ycAYFcyP4azulAq1FVpQrY0jG0Vp7fRGZeRYCOxHW
2AK1XH7CtK6LQHNjJ/l2Wi/3ivIAoFjKuLpcecW6TK/tcXo0sXf2eGNkTZzSOmVK
A6eybHOTAvRiMV8kgsrlsaSjqQVBNaAPXdnE0IdhVkVqViswjlrD0YPQfdVn3Htx
Ld1oQJrDchM+C+hwJAgBoYBMDLvqONDfOENBkDrqi1v16y9Ete1dUlfqSxTYiDy6
zZ+QWjlxBFgtouaqf8AydU/7XmsfCKZ/UN8T7h8VYEPCXDE1iiO5WOejnIhz7k+q
gU3+SCeX3JEB2S9FR5FaCLf8TF+qFNE4Lk914FgGMTwXjwoQeYxJ+ohpDPwKGhn6
5SxdgpWkh8rwt5DKS3hZjhBIaRLxexMZ0PusCo8PP13nkZHr6WKNEb0qEqKtjQzF
5psbQiN7GaHP/YKZfX3iF0QiY5fKPiiCT5aHS9GMbJXKayfJuTnd+8SwLRcAIOth
+36aTwa3i7vnoE2CLEluugkD2lSQk0CKxTvV/X+FgL4m/ktnTyMNmrWd6ZNHbJcO
55Qtg33y8HgstbhYbsoaQPzoHAOz29dXIrLf2YeNz9Fxexbl9emjauhWSD5Ho4Ua
2AJg9zqBpTC9GdztDjEnFBt//PGUJKhu8lY7C0BWPhfEHn87InZWuM4e4e6KJ4EC
Fu4ZbwdhHDVzhzVZwMgPseVTRdCoYvZlL8zfqF4nbufzntjvohqG9u4Fg7uCu3qe
P1qume/eT3cIUXUthQoXcDpXarKKks/ImQhakoZp6ZeSHNMoJHB7WUug+/9nmiku
ZZkoyN2m0fD2rfRIW7KgQBtooStalyg9n9HocThPY+805R7zs/UFAm9n+PlYbQqr
riCFBATgVNFeu+sq2fgx4wNM22OyXZ5Ti/crfp/ObJ24wqlaqiOmOnVHbWvN8v+/
s9Doqr3ZJruCrgQJJRulsYyYWlQNxHlkAIPWRQcIL3zaKIoKWHVwyPr8bJXdUQxa
kaa28ZiU7PHd16ApI7ZB250Gs6DROtucSu3PKAw/IBvEvxqMn6KV74oQVIAOrT88
zJGpLlbT5kdM/FGoTdbmvGgesDswUrP7yk6GzZlXWGLV23r4zlhuSubI19pLBGDJ
lSt2x9wowobf2ASioDSs43fMVnXEZRCn11FaRMwuILGPv6Jo44VYVB1I7lPZV3Cb
63ow2fzXFSWSQdjDRyBeIoAq4IAMl07fhimeppJnXS3f7r3mmQ+vxW/VhsfAg60J
X/hpBrNSGJbK/DTVACX8tNHTTUUyCGhoFMQF+zNNNg0Q29CVxoT6kWcbo+LMlMJ5
AopbdgpuozUDucKzNha/GDxbP44eC5mmFr2g5UcjRxgRKTCPGLdwtMkVI37g+jwU
1PIKTnB/QPZbpsNR12meOx3q+iU/idTpCTvmdXlTiuos4oUIYG8eN9nF2kblemY6
PZAnaeb+rVRTF7IHKC/u9+SvCg6K8/MqYBMbNJEH9Bw15PiGWWlLup1R63V29HdG
oRHa8HvUAppIVb+Lr32DEXRSnoeGZz6jkotv25wBbl5ERSs3FZ5oo0jBb/wFzquy
Xw2bpBfuXWisTQPA/x3dLR+a+K0r+cjV3PCowWtu81Ofq7TmPGM8miCPZHrypwlW
MuDdL8nKh2FDZzzrMMZst2tyVsx/BsihZ1uXrZ0Ej0a36j9TvezniOTElzVh2Vcm
nXkeO4TEznW2Aqzj5qQNP/gTUXl7OyvW2IWIkUdF/To/5zCqONemed+s2K0RJ/UM
LU/xn+9zSvTFR/dUpQFdjeAKjrnvRbM9tnYtvZm9Y0UxL/1jO1d2sutE7R1q21Uq
OJSCjyE+IjSvXEqagpzg970E97fe3ZHVzCgpNZS0Xxjm//9fhcR1GNCS4lohwLl1
X5XPy1f+Fy/NSjCHeqTjbMb1t6z7Mec1XfNkYakIXZMs+6ZC25GjZwkaD7dYdOyz
tcPqZk7DkgU0suwtfDb/LRHS/yA1QmBIknK71X4RrHeEzGX+vb7ysfUsKiZ3kr6H
jDIF16xM+8OYkr4Ta0JPIQ/jb1uAJAFI/AfYzySy1PlUjPgEdyEo1Tn3i69JSDRD
BXNOohltXwcjDOne5FC/RYzF/qHhPHvGySScRXwon5g/ixQt1GtsdMDs6Jj8n7S0
RzORaPZy/5rkYOLxLwPjkVTWNmJ4zcM3BwbDS3fAj1Tg201tnVZvIn98BmJzGrht
jwaQOhV8wVsyHfaerD66Q6uin08RcpgTXnBChWv2Sgv0lhwLmrTflQ01oqNMrEFq
1QgaXJFzrlVmsy5pQo+3P5xtXY5fQqoKwPeM/iTdAa4VF1uF0KfWTXfr+U5wHxyd
`pragma protect end_protected
