// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:07:04 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JuJmDtTOmOMheLFpmlnaNRiTXy/3oNllxTTzEQ9+YN4SL/Yggk8lQkBpeh31lCeL
/tYUQ+Ycdd90RvHk94qKfxO/DXEkMQEekVHiAiaHPvdowD16tfrn4csSeYurWWmn
iXc7a7yO0+BTqWiL3tJpYskp+tVMwpuVdihmadlcbp4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22448)
T1jIl3gzIvghDdkTyKiCLbsjCHUnrXKZczqPsy9dcyvuRvrT4CgXEHWV81cnmIs6
aJH+oyVjd/90BHKhWfvoA5Vc0JmU/O/whsZOCKpYQs60wkqkcRzsrHJfCgD2Uf8Y
c5rjYhV8YToyNPMO9Bo81tTLcGEtPuTQyfNEDZ5x5nME9QaTidRLBdADwUO96ES9
y1nZmeyFZZP4Vf+a1CMUtgOqYQTAfECfZpBpboTAj1rPgT3GHPHITgYreufn+qIO
29GFmrvvgup+PGJbhKALggqhbnjkTvXTRaFlltJqP9gIKf0BlHOPzaNr9wqyNxGr
elqvzFj2G+38fO82ER4HllgUSbmXiXiMSg1tN7A2507MNd7J4JscD65yPtJVQMJU
C2b3L+oe7yj/vhem0QFDicPr58o8ygngoeU//8Aq8eoaw2nnMdzR/JMY4tT5xyT3
3kRGPcd6CTNWI+S7WhqxMZxGnnFPEtubjva80P/DCy3aWsN8kgG+fYwqka15xobl
tnfYDBLS8PTIegbXI52UdzGN4pktAtbweNTvkNhW2ZC1kLCI1d5VKD1fnw46xyzA
dpAwVgZjRrEtK1dWylELBkG/ZHBZAo0Pi7deHWNQraTSGO+FgvvyVSgQoQhgejmm
L6TB/b1OWM+A5cY/vhtAu7Pqbszw5u94JfVg/LkOWOteohSevJrARahe0GpSkNPY
XoF5GCgLYVhNsGZnB5QgzRpIiytiKCnb8mmVQbciP6ZjFI/e+f/nvR9/58PPZtJE
Mb7pYUvK9q0/dTOTg28enjfV8mFHTJhK3BSuvzWuEkveLia0VRs4JWOgMFBePiQD
ajDAFPnoDFtARS/poxakQGmSGmuSSpPFL9rhd0r61JEAyACiIImKWIN03gR/Dunv
p6CIFZQeYoR5zfs5koJxCeqktlC6u150aSEbun0BuuTjrNoCDkGtalNCxZ6bCdfI
vEdtXEk06HheEU9wk4nY2tNLumU5cmN+YnDNYKTrfISaMD7XFoXTMUvodEfOZxhE
HFiTAFlaPnMpiwfoIdALTYUWxkM4Q8rarawTf+FSFwzZXveICMDNcq0BRUyrJsM/
vGKU8+zQTCwQP6ZhO3Dw8NfLoxwmRAUhVoYp/ZW/aJYa8nNOyrC1NBTfQxaDRQV2
AJXDf8Wx8r2PEh/D2Ud2+HeMdW0kY3zQTTGgNFHjfh2gbyWP8UTSIu8W+MTQxuBQ
NHRij16HBBm8z1DnZZd/8pNpDJ5f1bd5PLpf20X7mumWbDdu0AXStFjfV4bmaGIQ
ZJO3jrlwTS9P+S/XB+OdxeedeXJThTmF3zXVwoNLYyovSMc1uPhUXiREJhZYaOJp
os1aiecAolHaBNYnXrYV7UdQx9xb7l0Te65kRJTotgCmanCqWvNZ/WQQl98JAoYY
cbkStmoUv6+x9MZ4Bxfp9pb4IC2+eduzqeL5FJ26lC8dyBmuIwDzRPQtuTZyabFc
kKcHKUijbI+iSXn/j85nFwTeUpCkv9OA0JNMibvnxF9YdxVUqQdkYOexhr831pF3
OO9qmdlK98fydTf2gC+N9kxuRI2QNXevTo0GDhfeXJThIMX9qYmrHnuIpN4fKLOQ
wU6dbRr6oOKzXcE4VyJ+7XEbS8WRoQp3WeBY9UpsXgn3KP63wRQCdCpWJvB/vNPW
KOJWhiZjwL1y+Mik3mvLFKIxpnHJpp9P9chjVUS0ZEnuFoo4ZlNDbJUf4pqj62Dq
5Qv6qj/X2XjYKc4PjxpDmDV8JXvmQl3CAuCjAG+n6hVGVqQ1+lq/SUXyTBYNkLVM
x5z13AuPQmiZnLBBe//RIzqacbnYnuwN3bqanyAJhXj7YKKKd6uB6bBM6RwScPVJ
4Ds8ATQ4o2qiCf126EyXSFsT38ooCw5RkA34He+ooewlMI5Tr7m4JdfJP435ZQnu
St4P8up8kqPj9H8MarpuMEDrxOf+lMWy6RudR95Boso2kiKGCmbhOP3MRGO4aE+k
q/V9F00PI6qAzcADX7cw8+CrC8k3O4yQqtMhUTT9yiRNxIuBwk92pohfc2t6kAyf
Ia5Bp184TkRBQgoFmBEocvdo+ltVnbXoe3X3eCbjtCO3IV1JklG3dUPQxZYZ6ra3
Lfgr+cGkPpAozWmgmebH1k7hXqQijx+kbEsL9TaADi/PuLtoLD1bGrvemO3YExdM
BdCfy3hWe2PPZ1MOQPXkScgEVZsMTxeAsNBXwLh9GlD/PPQ6whrmeFaf9IyUGxxW
EgkU4zfv9Mp9Vs8vEVmxn0URkbrjuZobuanZn0zAowboouABEZiw4264MTchmVqS
GukwaBwUH2WM9SH8agZUrBjxt3539pqxZCodOusPTKy/CdqrzfsQXCuVJfBloel6
YtZ+MYoaP9J2JUAWx5UH2t1eb80p236qDxJQjk7JUh/8Jjo8cHgvSau9hCJup3r3
3RMfr5eu9SCqBK4iL9Uu3HrbfQ5bpQB4NuGRSUlpQpSMFkkeQEPFJtyGHXdyX7gp
FAxcyvnSnI2B2sB82oTZg3rsQUUsqyanMLmNBhgp5n6QpcirSf8RpfL/EHoXNxEl
wlp2gKfpqGOwzzOPffWnNQVsQWWMqrzXPvbteRFGtuJH0R5i0M8M3o3GI9uEBRKX
kjdQFgIidgBk+Sx5ePs3JhHNVBsTZ/586ufLvIT6geYVM8BmFLitPlXdlVo8acl4
JioBj2ZmeANSy18prLg+otyOTZWmmA6PemT4kNoK3vRY3/TQC3BIjM7KSy5FXQaD
t8hZa4Ct9XHhkN5B0ZXJDwh0SAyTXqMPo1jOAgncLFkNhWbkCk26EjkIeSFFYsGb
RNUCEvYWOjS2FEkY/fnIisprLkJyJ4NGibnlz9uSRkj3sb63sLHl8PTgA2qumkq3
JwzrXGvyS5/z6c2kQfswbnBH3rSUbGHC8MMq4pbarHIHwKC7NUbrvLI2Ryk4WtFE
cfmqej913j8ixvpmQ3nCDWF1J9BrE9SWYWrmsRhiRWYCfF3ceOB0o935F7Kc+fLj
BRFwnFd2XoqxeMLQjALMIzmgvshdx8ya2mQtnN3vsUEbZpVyMd2LbpJLKkciPM/V
/8OdOH/v3XD/feoKdzih4PbxPrVMIT9vc8nDKKyqtmSHngzBM+dMOBTEOljB5II4
ma5fw5z1LA/b9omV88/odb4RIHrrI8Jp3NpVy1byF/gUXsuo2Tt3d21WNlotDywM
Zmj7cnu7fOqAFbwZ/lMF3Fh/LsI1CxvIJUa7dBlFGvIRHDEFLEYtsDjzl7tBMX+I
aKJ8mCFx1nJ4E2KjeiG41ID3InYWEkWJFI7O4guhgEaaF998Eb9BGSEEy0kUsG/Z
fxVixTJRVPd31x5UyBLwlNnAaG/8MTNKxNkcjoG2jv4hk3Qkgqj4Os3aXujBc6Kl
v3RWw4SexDRPAl1/C4jHAWWFGrscnNkuzzBG9VyHBTjyIGlbb99wwbRJL02wSY6i
+5Aj1irteARWI1fH2lh6gCZyrx56mH1YzbFYKM8HT7fivc4/7n92sLE3F+DAIkI8
ySYqoXnac3EIlLCqM9vTlIXTT0g/b7eYzPW4R2cnailtmMIwP+F76j07CSo+PgzY
9Fb7rPbJZO+ld18h8NtBOawgdUlxKaYqgwph5zHjwhuOE1+P5F2K0IFl5+1OdFeU
iKURYIJtZdWZAy5ryEOnhXiRSg/nfnEckE6o4ki0Xh9AfvkG21jP6cBlwBbFSwT2
tRWQIT8GB42ktJ6r051ILSNK2YS1LO2dZqBUeZhkmSYy2d9RqGWEBPxLEpKzraiM
41sD3vZitxB6zBgemU26xhZwR8LWz7NP/iMsgCQy9qJ6F9Lmlj4ET9ANj3k3Z8ge
Gog9s6Qf8VQfPLRc1HsaG/6LApDKROKXX2/Tv68CQpO8lBIPEWf3FZGW4dm82S+7
dMBHqEytQlQ/jeoUQVcrIdFA87FExCD/PPLhbn7oKuz2upk7yYQMRwhqBL0Bq1HM
istIVQ+PuaQGs8H98kbqfjT64foChk9DwV4bvw6YkwJ4egdoDozgDpb2COAs+xEN
U7dTFIl60v7DJ+5LyE7TI1XqwOWZzwC6HaHIt1Pa98e9SUPfhP/kNqEV/x1Ey4WS
SbDhNwhOvwAyzpYmX2BTOfnpsNg9z9lYyWNDBnxkZNCrR9DvyeuGtaL8s9lx7lpA
f1XYQX9rYMoN4cRjBTGXTSk1DIe7XCD6vTG1pUjyRqoyv2HQof1Uflc22hHzXLso
tkut1bODhS8AfLKcJL6bn7pP2CjiTDV+iJwVhMM9vmYku+zTC3F3Z1LPNo7xDabv
l9mSPk0yZqj63Ht26FuhkQRuaMVFp7M6PyoddTUIiqzhOmsb6r5e4NLrBQxq8eq1
t2vOTTx4zDDSE75vV3rFrkatS69rZ/zZ4T+uNd7kVDPbSaoYSm1yIBoLdsrbQXrN
g/kTvr2bYd6cm2rOK6TvR0TojNC/W/yKPU7RRP5UPxKFik+lQTk0mXcHZS6I4qz6
IMy3rBPh4OG9SPzsRUBdVBszCdqtf8whzLenAP/1PNC/Czs4cXMefGXgkUsYYEd9
d6yGBgYem0E9b7A+l792XDHYXeGz2BbbrNnIds4x2fixpMNqG0M1qYKr8YrBzV8C
TD+QAt32bjZrD/i6kiAc8XvVnogflU8yG1/0JHpNONVXBhJPbHaiZbN4WasE5qy1
z2FLiwws66lV9cF8wMutHZ2mLO6tNJVjAKlMntYIFQmRgsUUW93ef8/pQbt0pnKh
jSVVB6RJQVqh1vA0kBWGBX25d2EcraMIIZQdVFg+shV7k68GhOVOM6IC0TwbaAbc
GWpHKKpAxrdDBUGWiVYrhlVWUSD5PW0DU5yTieBr9GkF4F4m+RpMBbGFHNLAYyJN
vXCLmLaPUWDuGQoQhmJ725E9wR4L+veGGsFksaxsYvsIfPEXCvNZYa7M4+d9E9ic
0cOH3V9XA/K6OXot8ZIp2h0Ti2D6z1arC1d/pmspa/vhfYLS0JI6WHLYLf01pM4S
ZJkAxC9pp1NK6E/m8SDFlyLUAwhN16VLvy6I55ZcQeAHg76hbMFYyoaZs9RTFk1p
QcTZZDAM5GrQ5jzYZ3E1iA4SSMYQpm/BWSEB7Fzssn79UqSmZrrCKqsOx413ATJu
qM1S4FPapR3GHnA9rI1+i0jPISzLhhbGwXuYb1+0jcy9Xsk2CVHlj+Hz5W9vJ1C4
7XEO0YG5OhkpeguUGqdMJUZ2jkGLcCQAsRXI7gGtRO1u0VOWT/IGbmbkI2r94EB4
Ey2kn6NlA2xDL8LHwb4OmI1GNXnlc+uVWNjAM0MQVQgFHrv1Zvcb2GyUeo+nhfWo
lze5u2/SO0+kKQVhxLzgCLRDclYI3cfj+3BGCtGlFpBpBk+xPxWhig1VKB4Uks+m
B95Z+iC4M5aGoIqswInGT7NWdp4XASfTMHO6tl68YolCFJ3gCj2+8FrkUnU5mEiR
0Qf+5pI5wiax3zPuJCHiNBoIQ5Fpx9EbZB7VncyLI5ZE9hrZUPLQd5AhHRmWF/oW
IT+QZZHU8qEsV6dVkXoJiZwmWbb1TD69NDLeaXqIEZNBcZVJXRcGBMM5vSU5RUBG
ZIJ/MYQS70B8kPk0aG/W96T2PV8raS6danSddTTN/yYqL2920gF+LVnJl2fQqnk9
JaX8xn1MEF4gHsV+KcRvsqGXMLkygpNxNEl4D5J5PP4RPjBoxb2nt1vo/x10Ik7G
m00Jv0yunUGSX2/w1LI4+mcuxjZdh52bAD6o/ypYHrPl61uOTUirBnqE6fN0vBVc
RD8JznF/6CFW86UVCucJL5Y9GeBkeT/WtgpL9qphyO/b8L61/ahUEMAFRjxHNgCP
H5P3y1Vr+/LcvTghtpe82hJaBFp06Hs0Smx/71ZJjWMqu+fgZiw8fXZLvt6izlre
+gVRDfljFmdPzXlZ/BcXL1jUx4/icmRket+H8h+oBWw5VskMCmNcEY7hn9gkfz+W
zEjZNBm9S2+eYXnu5evhchItwHdJJ4d8Hh/8d6lAArpnTZTUjQPjO0gly8OI8/Cw
Dpv3PTOnWCc/5FuasfZEdA26bvBIJZlPuK4ghNxbsrg/JogZ3fnRYauLyZKz/qdr
gnxrTkzsdC4hFKvJJOdeig1+UtjFRlW7jPiEhRkaYyNzWdggHcQY6hi3JqxJZNcm
afKPDofFXbdbO7iZ4vrT70xeAcg9Z9wq4H8FA6qD6AgsyyY6W4pErOtyV+y51GTL
Eec7cz0UkeDiWhgaE0Gg/ENNbAwOTih0gE8+JndIYhszx0IM9ao3HTWvi8hsGhNK
R2QyFhoYW2Sh+EGyLNVL7t5IMxb3vZZ/f7eOqkhLAXCh9u6+/26LOBLFbzjyWeQg
IHj7CQrkcEtw0SDg6isgM0Y7Sczw6eoKfi2K5OVKuuER+dyOxzTT6XJuA4iTcGdf
Luww5MuH/NyWNOcvRk+r1CTOfNSD1VVeOxeii4qzqYwTEzq40SPOzMLP6G6n0UBO
z068FgP+O+Icb/oVOK/YxAOL+myyNEPokCYkf47TwkJYUqIs4hrZZsj7SHW1KevB
yTUdjT3+kOTRwyKIPJTEGX6zralqk8gG1C+S2sXlFZgpzjo7mCPGL97i7fX6/I7c
I4dp+nM4w7Gl5VMcdht4Ha5Z4auAyem37I/bGDnOp+CUQI8tXxjClg9f4/V3pSDn
CEQCJYOpjT/l/cHlULq7LzYsRmSTiNUXFwvhvlnkjuys/Opctha4QR6XPxMxACQQ
YHMBlZtjzD7RBJ2IZdRLi3szvxG8k6RvFR+gu/bquVkfgMzDMoabl4cwpnWcmxxn
M9TSKAX1IFs8ei4t+WqjaA5hvaZqifzLu2yqGPNSq6mzpPF97BAsSJnEyzIAjU4e
K115mPBIeTWe9c6gkcZKiLqDv7C45fMNR0gd1s9a0wOy3EoZ7m03Ha6TH5Bviesi
Ik2FCDpxjxP+ZTyEjb2mUMoAvzFsIibiEmQuzXgxT9DoLQpANhU/lbjew/MgAa+o
+aTBjnlMAeuDRBAMYxtdYziwwAC/xRaAb51JABeNPG0q3WxmI1mwvFNdbep3xVY8
Khda4GFenodGVPbA+syCri2LRka9BN7LQIVXCPAlkHM3T4Bcqx/Ei9mCtyf4XlL2
NVdIKB8gxSmA/WtJKZnM2hgAVIOzd3ZUaTXOlAxjJaMhm8o24/Jdidq4ADStMg6r
9ndCo4FE8KN1suexKG6eHmBZCHMQMI27nagBl28E67qQDmgD/oE/naa4onBDBSiy
KU6UiucCF0OByGgMiO+DVxYwh2BVYiW08xr/LWQA2gq/agkiQn3/gk+OnbGN+nVp
3cRzyM51PoDHM+jMX66yNOVjMZE+2GmAyGVb6Gx73r2csyCi7qJIrjEhd44ysg+R
/vxEZbtkwJDSc4yozsxKyb9GvVY8NJdxa8BW00gzYgEmgPU1M35fZm0SeS7Fwhfu
bsdaOvzxaKgsx/tmo2wz/+8NIp6YTPI+z+0fxdWiAN28LhCAnch6kuFGE8GSU4ja
kx3W6X1zf5PzL8k+RGguxWnIISAtLJsxfrlIchBNjv+mVmB1jaovqRde0aqO0IUS
Dyezhb5BgIlFXeVGq+fU4NSPBoHRw+2Exre3arCjf/2w39zQ5Tr6xOPSNqPasx9B
ZS4E0RDxZZF38l7TSTU6mf7520WGhCJLOPfvFWrQ0GXl/gzuB4E3vbFgOeDyKFJE
W0VKyEwNAtH+XOSGbWalEqKrOLJugAXJGtAP8IZLLArMi5481fqbI2mKoGew1t5n
KvP9Mdnq2BR424dEpkLj2egukPkswLVSyg+fGoPwjuXWJYSNx6vxJD+ohXrFm4Qi
4prdqL4RESLum/+ZN+LMaUnv4oziQ2RC3Eo1g6crbI4YQ577u7bR4jQunqWEBlyI
33ZQ/7IYQRInpVG4VPSetvX3LSjvPno+LIHiJYF5UESBqZRFgVX+JDAnRmOCGXy9
M8MvcrvMLPJZI+THaRgXQEtOZBmGyHWq5Vr/tTnyIsNzsZRJWeEPJzobAxUQoPaE
jhHhR1VFdnjIGkAarGn3J8b5L+7AjSlKCx+kW1KN1UuIGmE5Gq2aJXyx5n9CdqEg
jlngfBR+SOxxBlI7DVdG4CsO1vqyLVD4kQDRZln/8ngohq5NR2wGGLLgPEcdNZkX
UG/592a06f1jFaIjx2TyTJszWz/9cj4uKwelD5kYHdkHMDRJVVFI+wPI8A0yfGMB
7io1luS0G+TR5F2onYHwda7D+Yqn+LOFVcEPf+8sXYj4tMg6xK7hbxRhp28EzSL3
/F8Wqf9mKdQbVcw3ZqxjKD5KrJ8OHu2vErE96tExKTjuoOSqJzUBF+vLej+X0M/1
LJGwf0RQADzXl/b74q9SPq/VfcUou4Z9Ugov3MeCMBzOZhy/rfg8J9cXtsxqDwL8
2ctvNkv2N+YRVN/QqkiNPZuj9Liv5JZRpPwFNK3u4v4GoSdeJKSxo3ZaFkVufOHq
IAxOVXLFHAE8x+XyFDxdDOooLKpcr8oN0QCugm35EiFu3nifO87dcqqkBwRY5ROt
2R0HOb7jJNOo66FIx1cE/xjIOSTfFAza7m63fJv76vZiDDk0De6VVt1xD3LrX2ob
D7Mkvof01fxR4tZiTlbPjBL6Jvkvy7dRuNRvnK0bn5HD4JxP5lL5ICv+KHcQy31h
64qQpdqyYB3/FXab3VTEii076CVNiCc4JMfHt+2ACmZ8j2hGWtg6pXm6oq9LYI0r
KetFMEOMm7RXZOmJvJaqEmbvUNxyU5MO6OhODBU9+RLSljERrSirHOuY0I6Hsbzx
PlrgSXFqe04/F0hY8YtGmvjNXF7UBh7bnCDMV9tqegFV/deAwaB+IkdjTdMtA+hY
er90zipGAX6p9i1xUJC3dOOsdUeHDWjYay6jlfni/EtcLTTqrqUZ9KQZTYHawSdY
eYJKh9aC0HpQIlA07A/+2XsJqj+x4GrldXYJdAcC1aQE/7ljkAKmp9Joco+6pwaZ
B7SI1BToxcNzKVuCVn0wNqDuIbvVNG4HTpGnigiFW9XJMmGCvEfuZ7DAx4GeJ0X7
iUtBSgLNgIw3OOUSO3BN1MA7MPoaUt8aycl8d7WkrwDD4KsZJ9MCPqAJ78g0RVwH
1Alynf2yMz5tx3HPqmU8aaZrBtcb7iBZWCEcO+evN+6ciC+DBNR6A+VIZN8vJGc0
6B3OOFDLA+RSAJa0W4xJQgClCsrms9NFNLOzoHOtY+B/i3su9lPHzkXWBRHpWPvV
StB/vbse7xx4xdLV3gqnvgw/bIzNPxBA9ax+GgyeLIcBLussbh1KemxUBoYcK8ke
C+/PypTWpZodi7/Zy0fCBO+C5LuNM7KxkuO+kV4nfSYUvk5JyYJUXnYV3OAXcx5O
mfkwiJQ1/LHXn8q13QVx6Z+2Wq2Pcr7NM2RZ0Bh9vli8pE5iIQqyiIepWpPeaX5V
sPAF3Ip5QKulZTSK1R7xzTtjbs4PQ9HuJH0/Zul6zpGtAuFCERhuTdn6KMvHDaEg
f2QpU521vZHvyIqdCld+xRNyyJWvhuJJVHE9h9VuZdkfkNpa6u/+d3txAC4Ij3II
66JWH1ouKhvIrO9IQy1l57G980jziJXoyyfjfkZrRnBpZuZJHqQDAR3hcBb1pOkE
oI26y+y8DB21D4Ob0Nxu/gyIIWA/M9sro7OKDvhVpmpYyp02zG1xID3lr1GMz9Tq
75vHRg+Cf+29U+bwfZdZeIydnM6tztXWrL+ETlTfQUc8uOPVKzA09295YjS/SpSi
dWv5UUl8l1FkNCB91KVAqI7IjuPU+Llja3Irz0hULGOEdqMSPuVO+7OSMBbu2F2E
vbX2KjnMem+Td0slBT0Ce4jEst3ttvnR34N9E8IQldMQvHvRrvcCaOBsNughTKrF
9zOsv5cOGEmbEihdb7MCJLLzkAoxMIFr4xlQisqWsJgNlavAHC0pYohVsIFTzyMn
j8uCbH0oznEmGpFABzLxiye5bP6ZCs1OwaFnwuCNO81fAb4sYLi/vSh+VlnRIJYD
lLtUc83OFe9QmvyALAEnn1T5ntNOUKoCya6ny+IXKCyBe43a8d58pl8G5LuOjF+C
gUQu6IfHMry84tomZFwL5ikC72EYVSLL+/O/HORxd+lloNfiAetmZ1wYkxRZPF8Q
+8iBaqEGGvHYbC8l4K501OhY6AN2fJfrSJ6ey2rX8OMblyUnAr+qALpl62JuLYeS
6Qck87vwUMrgtCtgPfJnMognxb9upzsWLUSUN5pJIkBr0S6vzLGfkc6BJC6YL17Q
tl3Obb87cl6m7fwj8mQp0hcggdzZ+LggLK7pyCQOL0moERaY8+5JqPAZMppDyGU4
HkTXHk9/n0Szs4WhdyeV43T2NAKO7aetS/zwftuCyRe7Le/FEdo3gbfzFsEVCH/H
+N9x5IKO9pBRd10sK+RHUA8I1pzYDvoPnra2RwTCtTyxTQWDDSsqjHuFMc5vHOhj
ku1dgMEOGfAaCQMoWfO3AAk2ymfcRzZ6uG0xn4QKD4D+Sfy5XM71djPgLerXa8RX
IWB2pUeGnDrONGHOIUFRmkuB3oBvJSJckVDN2+2CtC85CZLxF9GwfMIEs/h73ZUS
fjLS5OfmykJJ5QUt9uQb/p5RJCYg2ghg+qmT95GCrQI5ptMLlYquTKv+UPGoHqqC
a/45NsfIFlxG/TE5XlIQTvH0KpaLJ6leXhODGNl7p3dDVa3f+R0tqCrKjlVG1EN+
fWd4zM0zbeptcj+FycpoCwaK9Cq0sSyMhzHAexL7spxCnWVzR6JNr9r2X/KrPrVi
A6kCnhcFAvH/E6ojki4Th5/33eyoBjpocARDHqZ+r1n7XwUcrSxCSnTe3ajlKwvq
juStXMBa4Vqk8gDp77BXe3+WCu2fBDFwR84w4fBVDA+pRQ+bw5L3agmcRQCaiM/k
MXmB1Ewax2SMd0RLw/iFmZF3A1PXe0UfePaozITs+hXdfH7TcDcItWoM9Oy9zjg4
Cc4okORfbMarW4JqbYYYJ9bnEGRCkzd2VgbulSEQoZTBD0pCysLwEOxrDY0zMJ6P
Y2HjPDZ+5/qt5ZBAq8xqoWBIycyvAWuguA1BwLjDxyclDYFWsbtc/u8ahuY7uaNR
HMQcOyYOVDsHr8CiDEA+wD+eiYzTw2uu8GfuLwzIREbnA9xvW0P+U35Sui3JipFr
l7LxqO+8nhPl0HLtBxfsu/7RRci59uefFMYrTQmCA7iWsojM7xlKgiDmAHz7uyos
+on6Cu0MQO4t+Jnm+SDXkUeXIschy5/cq2kU0KLXG4BDTLiHx2+cQoi2g37A+/zN
HUZ+NQQDLmJ53AudoYRhQVGm3l64Ns6ZJVQ5uCl1Mu7DJScduy1l+fHCRS+qr9rf
lqvFWooP3n6GXANBCZqNZVxFhQ6wEZCR5ZPh8AnTQZKXXX1lqHlyaWz13S2Omnmp
FcV8jvmXkhAV+oVCgNlZIxvOdDA0I45GNE+scnwjCGM4RUqOI22kxCotmn0s+eb3
lptFLzt4mIubWCmi1wwJketh/6ugfv8NIbmkJpAykxoTJ8RL4AI06Gk6e+SzK2UD
t4uN7k1Y8l69qen5Y1lOzWBFrGGvOGV2MAcWaWq1ebgYp80EMM76B6uWCJXaJhCJ
dBjd6MKc5/GYmZtgMitfMrW/aS7IKRIYARkViGcw1Vg2tpIPgP9yga4DKciDhPbr
O3cfyQz2N/8Gs8L8K/LAxLPwVFFUeVvtuBZ5dcCPc09Np4ZWHSXuYJ0gNyQixp8b
8u9npEYVRgLvjwHXedxN5mM9pY56j/Ep0FQu/+1DEALVWwtdUWjAxgzsStcLYu/D
+gnADNUOgMZUYw8WPFawDbsD/xCbrtbPCWD7U8vk7CB10533T2ClzmRuiSwLS47f
i+0VELUHz2gFlCv4amnjLCPn/6Dof5j7Rm+YbOd4dIYiS1OTZZ26rqcubiLHhJwg
DO71441k9SGM01omp/i9IHdKtQJXL7J/dXyZJtPsmj7fhZNUDtdMYesD3/UaKqUm
zEIZzCNg+/UIcTyMJYZGvel7lUoHd7gWr6Xkfr7Q26sEDqNpYUJbmIXRgFQDE1L6
zxnUChoA1St1hY5wxhl50htsbLEfhxwT/0eOkaygweBAio9pL689EwLK6iM6F35H
5IS38gv8kfdxhszK2Ig7U7RMmOyH6kmPXrdN1FbuCQEU0fcuIEpoj87jsX4O+p2W
K2UNxessn4S6954riVIQlI5W0YVxlsPwmHz4prbOZPzOf53Xah8XP8UTaxzvzaAe
mX3vnLuQ5zKK/mEe3uLML0qlQAC7WLd4B+MjojHXdPBfCjTViBgqanbwBXR0A1YA
/9x5HGc1Q3WBZQS10FxhiEpepmDvULZXHHW0YUWqLW1mWfmQYEIXYSCaZjlat5Bo
wGvYwtBfmYl3pWb7CB0cEZeNikxv4U6mEvYMNA4K1DdTjoCqfiHya6Ff9srxPRo6
wwHPFMXO6KOhgmS5e2feaGkOdycIuS5QT1ze9au1dS8hGPw+WgQkZeQmDWnkz5ib
Twa8ry8madSQZ767LKvyG5jEe8PRL2EplBANoFaGCNCSdnBK+B5fwSr2GKZae/jt
KtB7uZvuQmjMB0vhCKaO6PwnfUXKwda8F62Apl4e7cKvQsEoq4MKCYIOibUwz+To
mQzv2Ie743crG8Bt+W6yB+5zCGcGFWfduPe+ULI44AaF2t1RjnDCSfOcMJ7wH8E4
HVYrGVaEEpVlLeBwmpgJmAFCB9SxZCHG+ySy/L1rdNLDGSjlRLGirwJEMOUUP9v4
FGQxK67HSZherRo5IqEvdfBu/UKNrtbjh4mmGVRzFOPxaIJvRtnJ8m4Cmj5hggjO
JbiIJMWEKLdtSgm/oyprp8/T/wO2bFGIZmSWmT76SfsDZutf2wrnZ1rKnoFH+Csk
jmhM+8swxJWEmyxHRBsIHRhw8+to3DqOFEoRw1KmPsxnZDHrb5bVr55nxsNfx/Vm
gtJrK9ThYBbzKYUFXUnTDLEC1rLyIB0dAT/NsetVqJ6xt7DohTgLIuN3g+QIPqNZ
DiCZbRBbD8uQJtP+IriEwbP9vAV01ZPkgJ1sqZzB9sP9h5u7avH2TLvNOcGty1ZU
gFIpRbbtCS6Ipqe1L0I09W0OAID8u2V3yuS43yjAfdQrMynsHvHGCKw7vfddu1r0
hjCt6E7D7jEovqVGfxtr+zcvIPYJY4dQQC68gewKNvI08nRtfxlZK23we9NjLX5u
ZMf4cMP3tC6LGOCiY0ATXBAZqBAJAjB9fHYWTcfn0DSvlp0XHBBH4FUR/w0Rv/5N
wIg8xQKJJhhz/mnA6rLEpKL8EA+Iqy3z8BnRE4gTCqenlHA0ijMw9yKicexvgnxa
otYxJR8QOe9iYlNQj9wGbBSLzpnEoM/1bYXVUOayOpVZZMSsguOGflsSDeUjugNp
d4Xgyu+RlEVsSFzvSV/5+gnowOz0hWi0Bmh/K+gViSzlOCl0TKqjhYu6GBmb/Bvb
RXcnN6bMgsnd4jLqF9bjWQa4vtO4BmGyeYfakkNik9JW8855p069wW0yC3Nw7Qa1
2fpATm6tATi1kS8UOPRU3tUw7Hj+YtbcFNV2iX478PsrxRWJLgrN2dr3HF0QksvV
KxYw4i/Y+KN/26iVnG/exql0U05aJad0ywP4MWsCcgcuyaEPvyqjNo/EEfkIKlXf
owfNTq0u7JI+o0VvsNetGs+TdcxP47IPpe0/mCWG6TIe1iAZdBSoWRga4jjIwuNy
epl8FnZa2DoZiAhaphnYnKcPDq4WIMdXggV/L3V1zOvIgXQdf9yVXAj4qNRSI3Fe
wgzBEz6r5wqltsh2DB7M7N5a30Z72I2i3C4hnZHY5EGxrn2XdyUpcEV8xLnRC9Bj
dEDEi7oA2EtwwweDQglWkYXmziHyopUCId14MdvxxUWTe8AcHakdcwDoXnpi21ES
gJ61I6mp+hkTaBp29wUgPJxklDGijewiSNhHL1F0enx9/Mw0s/2arkl82lLkOA+I
uP98+00aBPsdJCimQBfXAie8Z7R2ufOeGSRafDCI71zkGx/UqVbr3htPaBC2GLP3
Nl7GR5a6br5oumfmOYfhxB539dLmhXisrnQQZFDlwr95pf0msqHPBXJhnMZM7pg8
6DCSDDyixOSZmgmRLGMfqCSAx56yRazeQfg1orVomYC5XJbSpz6sPDmdGHx+wMSi
lIvx/RGcU7FatByMMIOZWxTwTd0kT8NNOAqokTfGAwx9Cym5hIXvWzbOlVQcdH2G
6FDsIkd/gc/If6NdGwFY/S6OY9Hz77PcG6hVp9w/fbs323Slmvt/D5oJxYFaXc/6
7vi90G+V0P+9kVdgJvSsTsi2px/yDtkXUiLTJ8D5KmYPbN9m/7wFceZiAt4AmH7s
374c+N+75MhKPPCKsnKcnMF5a7ke1dQ92B7UlxZZD1198I9TYnlH5O3VV/tAqLaR
TJ8FTIQQdtNa6LXPq23swE1591QfGpAqTYifeLJjVGX4thfq4m0YKy7Mm5nrGI4I
d82UeisyRsp4GqGOmVtH94smCHNgFo0QgtSTya8M++iabU5uzh49WV5/RM4Vsqcc
tesMsSPxwIH1hZ+0wYuaAUCKqRgpomSrT9N23N1pFwhZRc4wql68VuVRl8qEOUu6
nzCgDg/1pAbEEPO2QmFRqyUlpWyTrgIXHouVOY9hHj87ZydDzIvNG7dV6/2er+ye
urqLEeH+ud8TqWcBPsqNsRgqnz6HKwZbf8VozkyXQ1p7WSmcv2qaX5JiaOPnQpx5
7MV2ge5tAbTtHsdPxnlelzf+EyQSNhitdAMVpt6jfQ3/H0qtcUl/WteKQotxFjZZ
3piywXQQgG127Zcj5P1aidMX7QbuqAmdLVd72JVIyf7ZAqukYrEau/qfcoaM/Fca
DPZf5NK3aXv1GB2QkeGoCFM5Q453EITAtLi6tjpTIodbCSayamHMSMy1UpE7pVsg
cmf7C5XvEZF9GjnnRKu3RH729S7n8uElf5suIuX7kV65C77/zfohZRqTBfKMEpuO
+li7ChxEQKkZZK/46GOEGzMx22tEWsp0oCpVQfOmXtGaB5MYIgPrQRjqc3DTIAEO
W9CbpIxVVvZFajNMzlxEvEbnFXacwrf6rRcKXrwu05DvqVE/pb9SmmHKHlcLKTeE
rCDqKj3CZXC8f5nOfnXsoYHuo9KVZTgNnZgLIj32D4jRrTnC/WMyMGqqzMesdeH7
sr9B7x4WKdk6QcTIlSlIHlwjjBSLYdt3TUSmAHu+q6hdq16Ge7KAkdPd9aEav8PN
4JF+yqR30ydumTVBM+cpltO4rU0Y8nqKoSEURtNgvpeZ71OtQ9qYhSzD7ZE7KcYJ
bHuID0lp7/47FAdBEI3aFoe49bIeBcx66dPS1no0p+AFiVZfZcq2fWoLOCRRdAvL
ZuEbuBuI6FyAxQXpx+Nq8fREC3/jS97t3zsxt/vqlvU4yQUMYjcl8axXk+u9xQt9
huo7JOTwJ7jIQlIuag0EP7dfNGt0fK091ixSe+276eZhs7NS3X8K9u8d7xf2cpyc
/PzL5tl6cKO8NPzpBMOpaCHLm5U9lbvRu3PcHlnt26fefgxePqp8LhUfksitJTZJ
AL+IHbVaC3Iss5eW9+ICq2iegX1mFYJEBGJ7s8nA3fDLKZbohWIXdzyeUEt290pL
RtYAJ29YOP4Re39X9cvPmAo+2iSnJAR19CZQDuut+6Cvmep27Lt1yQIF/U7o8FPh
yiZU3PY8k0UQp1u61Uw9bsSmga1eZuvHCW2k5YyXUFRk/gRS6ZuvaBQr7RrxzWs8
4A8a7KDeiKX7owRzCCHcdYIqfWuin85FtQiZw9YUF/fVZYcx0JcOhAkVoxNpFndY
uy6iKpI06lVbE7CF37v+6rStJpNuWOBrYVX3OsYBpir2SNUngzWKC0E3z29Z7rhE
sj3MTv3Pq8XdsOjEV4XP7B39Tev07HS9JqorbUp7QF44ZRgDhm6TtDH+pxrzqYAW
ywbNEkoUCtvGtKAzsYSD740i+4MKiU3rN5DuER+oEfXMlLglseqSBEwWW1r6XfaR
SJw0gkmkOkyVEfZ2d1S2KVDBqoyOl6dDGOYOMpNWvuDxHy0a4bjmzMJocCvXG8jG
m2mPYQUR5RSIn8rt8dbrQ5olzf9t2V4c8wsptZshTtcylSM4Tw5wrI1FQ0ER4xUQ
yQNAUjWVoi76sivyRKxXuM9xeP6R0+wxPjrK+nyZHuKFhh0zGV2yA8fPdXI7crkS
RLy5yZmYzVFzIY/s1u64PFtWvtrdiZ2NAp9VAv/wpc8uTCzrPW6MbstWPHgwGDs1
6i3+hN+G4j0TPDDJbKpq22xBVbpAv5s430+9ubX7NMv/cLIFB2dwEFYKBQz37MEU
QN69S6CScqShREkWCcb4cX8BkETC/ftb+LCzOrV/tGqbr1gbMNYthOUA9sYjXmFd
g2g4LeYur/k3nC8fPO7JhUoe7isSQrI4bGw0P+Mkns76iNoVOBuwohH5kcMbtM1E
TJ8eV77gsJ+5XbVUqxG1mf4IuGaqAr8Z2oWOwzjKfbndIanJxqluiVUaf+Fne5zh
sAcgl5WN3vCIR5bDUB2Tyxfe6bPCm3BO1n/8CvwiWi4WREzEqZcsrE0NL0juVWKy
KiRjCAQlzQdrKnJ3y7qd+JxuU82J4UrlSyvbU+/4pFZGUYjSppEy/E7twJwLmuWu
a605Oly8J3gWIPDWW3Zdm0OL85T2YWZfYEqp3obk8pJPzZU1TUEnDM025jcVbKhZ
A5bfLM1p4/BK9B13/SzmZTgkLVKoQFaaQtgOOz5mc1b0v1tpoHK2LVrbIVpO/xng
dLXIqhBqkyhO5OqvkaBpsquW7g9Yq2eGSoUIyUjWxEMINIWmln/HHMFObSV4qYot
Rok2leknj1t/3L9J31TTb1mwyaNTSIlCozKuVd9bCQMUZpAyw4YRGHxZPiMn+BO8
rzLIpTGaXblEmv+/sC//FwDXTF/MUKtjhcxZaDoHapv7/OsbPMfMOif4klEE9AQz
7jn74HpsCajgzjUPuuDWiJnWazQGfSWG6ulSBkygw7Mw641WbfIIB35ryQMHhc4n
daVxweuzcjUVUi6RblD4QJ1oLCY0X4i2oA4sxC7X2YJ+c0/8rXXPbUKogf+gvvRP
VXv9bzugOirg+Q6wE8lMXvT0SJaCRzTlrgT8HDFPz/f8CNaiLgl2MzSCfNXFc484
goyM673t6xAnTCG+hpKzH1mL09JbLKt1nFshQjy1cyAPyAgijRh094nmnz+DqwuH
yzd9kQwbmLBanO45mYhMhsrG7qsyYl6xi9KIAm4I/I7w5LjNccxzEgYVX7GkK4oy
yojX2TvH5hR0d9hC/hhnkfoqwzpy8DH/qpl891bMRlh3pILEuReVKRKydy/vayVz
8bw9C1CJbj7DpQwAZ+QsJwnskzW6+BDDWOqaQADvEa9BMqzvxHL2MZ7fJx1bKMGc
RPLIK5SlXpstbcv9JIc1fxnKPXn30xsLqkcbuH4XfC56eI5egqEhrrCh5Yogqq+t
p0NChwerdpvZys6h2zjGJNs9+Wc5GT9PE8j0qiFk+IXIsCiPeUGG40u9p+ITbJr0
lTAX1FXewG/4MHjiZyqGo+mtaB+mLXNNPyFtHCcGlIL73U1oPmP48eXv1xwgEacP
Iua5f5ahyrZuW5EHmXi8D+Ui14VX1LAlj/g5B7nMmtmKRgCyt/OCz7CJHUS9Ow9O
yhcjwJsa5aadkBbmCUmwDo9xZ3yiqAfSi1izbPMqpC3tOGar8YHt9vGGWajtemOu
EWylhZnDCUX/pszEsxRYJCXf918I5es7CI/Y/8PdpmZ/dUawKT08EmIWhKPRZdx7
8U7YBFssU6S+ggTJQ36iU9HlI9vC/q+B3CJlmbUSgIslkCh9vOWLYl3TUxmgRkIT
q2Vtuaau1e8g+XQ/XgcexQp4Sljxy98n47VfrXh37Su6VJN/OkweGsHbVl/Uj7rz
FrJCHoVycoYnAzP1P4076IQco5uB8RZ4F0EV2fD24gZXApHjGy5VHMY+9BZjVblE
jQ+KaZaw5qwCbAe/iByJWGWqKOWmncbIj7Jr9j+zRGqnjyY5I+T2x7+MQiZdG7cy
ObtD84VdhIa8EjhFSlM1sFEWNMMgYNzHTfcBXwFPucYfYvNfF7y+IuKjTSRHjqoF
jsE/iLbetiiHadhGcnZcZE0051XsuwCIr1FcGElQPJ5LkNmT8OHj8pAr7DHpMEjb
4EXd58eBri/2gqY2kPYwc5yUxzrLFHShohz9dCeqeNX+jjYoXLL6FglffDt/U+kQ
4SgH3cLWQrc0s6sZGoZdD41nATxYIqM/Pyw4kxvnfUfcnvYfwa3YcRuLKD74YWO0
JXD2P5s4xMNvh1ztEGMDkE89+ADKqR5QKmgnteLHhTkUeIs3R1O+6ccSw6DYUCZN
8kleX/YB3+JFY82sbIVd8kIXXunZeQWjptyxmItJ5g5gAqTZtge80OxS4U2KU/0A
xPDflWZfVKn5B2rlJ1s6WrJlHwfFdyynlfWbJXLXfdoi4NgMUCFpiyHsJxd8Tpgz
R8BJMeq1AJlwuIYg5hG/SesoHPBVnayrQ+acmZFEKAVLoYBoSN2j/C3v3qcCGe5y
Za+wwWlMvuwvewRtDhzNIWTn5T2quOhUyd4UPfQguiHuQGqJBhYgWbNLA0ajrW9J
nVKLBMXERNbnpoTNQbkicCfUdIT/S5fy8CSqpSweYcDsR1HC9qMzu07Iz5dxg+Vf
b9X4UGZuKeoabR7veejHXv6PN+tYlgjcHMVd1lOxbS3EMjTLrsqpQqce7/qkOy3P
lLtEtII0hyS5UQkq8kIYYQ8ubE+G1i3ozDVIIctwAC59Ht/qA+62aNsx42VsvHYN
ulywSI/ePYOqVBeEWpZSxWCIz5mOZ6iwAGWMTFySzcq05MYu5uEjXknvNMfzGtcz
UxHmRJB/Krf5ZfUrZNFDEel9jITFQLBty5TG9pAFJDE4xH0w8KbwFv8xar5k0l5N
6zH5vyBVlhg4Vn1pTTtQ4z+7cJWOu/ZnyAXd8d6hnAt5V9Qw9FMMYNVHnBLjLbAh
UqJNu05comySOFpsFDLLzjQMIbRWboVRU/mK4hVihafokZZeJIBNGUZv4D9YbiGA
kXMX+CLIMs7EP61O1D4y8hRfY1QGDl9fg/iHNp5enAblz/MF2XoB4zkA61hRaDIG
uGFD07EJgasccdT3NJ5xNoVbR4DIMzR89d/6bB/70KNzSkOQ6fsHuEydic9gK1yO
nO8tVppIXj8xn93V5lL1ekd4jZ7yUsgOGPnZZ3jp92sV3R2+mip7TptymvBAj6bP
pKvQdWH7uq9Ys/EwtKYDmaGR77r2tOaPPoV8BrvSYYvYIxEIZTJnFJAEhEqcfYZO
mobxrEmprstqqj4+s5KK1Fm8VdctK4n4sFTb88qSm/rtaAuF7Rc6RuXwmkSCmJsL
1CyvXtL5JFbjvtKKMsaAL6Z5Zl5haLr5EsvKPQ4KFwtgNoeNWSH+VyN1gcYRjeqd
2IG3ILaWVmlG9ESRe+wZDz9ZJKQmP6+dfHrkEY3cU9Br/K246+dReQ4jkhnODDJD
3p30E9yL3KZQkmvaxggWugxyMr7OxpjPDnKFNdjg783a0t5jEpDnVP5+901RCYxI
vPwGkaY07KV7p8MVxSamYrBOeTogqnWHA0rlvRqe2L1byPBNXr6JnrOcBA2aTQCW
UfYXUI4UYGGWN6yuapJ3FRMMD9jbbbkl6PYPVLo3vmYC+/vJmF+cinwawBKkBkGY
EHmmoyzRHap3jWAeDIjyC234qBORRaezlwe7XJngms93pOeNc1SGD9N226ioeIxs
GA8snfKXLD5HBIhdd4P3A145NKDFkCJSmtAtr6khEgnzW/PSnu4dTLRI9frlYimp
i2oM5+l0/ifBgilCgj+wPzV7l+fRZVVkt0oe/AdZUu/lYiszyQF04g0hp9vjwXZt
h/klVYm+x2aIkq53aLA2ep5tPB7TV/3JAJCcKfsRnAtnPtT7RTVbyyRH04tFzldE
/pAbKcD8GN9Kx5EaeA94VCrsScZDGN3Y5fYafi3uYjkyRnedUxtTTQR7GLwkR9Vr
uiYa61oN9f7s3KA9WjLKBoE/2FBTSJ/+Qv+ECklr4v1ItMDDOEUi/q4qIEeSvaS5
YIr7WGKcTtABYpS8lhdIXfGD42wWg7FIC9it3JIPr5rVqHkjg5QOMRiwhpDUmUzh
NAkpSZo6NsjA72eGXVm5uvb1dekyfgjh1yL3v4zoeCxnuDkQihlWYqRrxCsjwZJC
jLgQPySMwqmHQ7qyS+fedAbpTDnuTXtLupfZ8DuPzH01TQKWOLom+OZ7l4xhpcSW
VThu6kF1yHP+vqMwQbz9c0WrSnVGdkd1xhHJ9W30sdLClfiobIl6nFW9nE3reYrA
br9YDe6BJZSJk5/3/IptROrpGME0tGX/0780uotohAun26CQQ0uMgvubrTh7COPt
spS/FLsXKr4M1bnH5gq7wc88Yn/bWRt5f/PpIwE9gBj4FCqcjzeOTlUKTAXyvfM3
/CAVOFvYb+piiSY7WUk3dAtaQvRryvtJ1ItYy2fcEfolIOgcG2DQGeCQlGHcCCkF
rziDMzJUKSjwjSb8PwNO4fqygfzm1DRuLIp8dj6mjMHTQqveXfpS+PIGyCyApIxk
CdpzZ0pjBzv05hS16rbcIY6Lnw5a4Ehnz9a1AOCfGQJRnbr7IhZqNZlDZub/RU4R
jBeEDhlYnHiJQAPLiPXi0JX77r2kzVQLgPByZG/dtTUkcbfiVkvMH2NgxR700Ir8
0WLfF5guryn0tP23bNh6S0zibZIkTFNrHAf2xWNp1yzq+u035LHy9+Pjcz4xtJzo
1sYAGoPGDFkQgPwCzU12WzMmEmxl3hiGeHHG0yR43kEDHqEdtljKghvX1cRKnAUd
MTXh2VwP0wTyHQiLildhXv2u5qFpvDy/kfbU65S5MTpnHOQHOE7Sbs2HUvvb1OZf
Bp9ns/u2xAgMWvXyVvnSXCsAKUD9kRaFf5Vt+4pv7FLV6IoE6c/XGpYbFb/Pel3e
MZHpJ49wpY73tbCuzCZSXfjD+oVAEx1bD1iWWyDF1SQjic2E9U336OiZ8k5rb8xd
4f89Yym249mzoh6k/fpk3w5tv/k9wnsCyucRn3RSxT5IJB5PjvADiPZ2NbHKyxnI
pCmAgCCU9cgGiswqaZLLawj9lQBRAul9IYfT0VKs8ht9jmDKw3Af9zfWTyrQA9Vj
b05FeHwRk72XiLs7IibI3uofD+Pyfd28z9/4qHHgBXZMicBCqAoEboEiVNdC7D9Z
ykyAqOKzzwxTf3RxcyJDlZsvxwPS9874Quyu/RtilGtMYLxXe+laQk2aSgQLEpvF
adQ6MIQC9OxHyp7qrhr4ucZRPlSGb+LDbJgs/m6QU5BhvRBAV9qtKHmqHjiqogaB
SavTUk8bd9xTYYCoPyhbrkYxpIQb5xV+Xougtp+TKrb5nQ7ZQHPDt7z0f0IqqByd
UhqlyKuNg707g5PGFNU3moxEjr2afj1/THBg8Icb3JPKgEXLrYhVANzA8JYGd6P/
t8PAcTtnywEAmcrvb51tbZm356egOI+6RIiaOdbxMLYRG7qDCiCe9G78Ym9bYBYC
guio03t+Ea2Bil7umuB3/lMgrZ9kRkb6EL8auD4ES63spGd1exAr0mnhS0Yf35JL
LQkAKDINUJHYbattiG6IG22WUnsKZpUi0Rqh2TMH1TBVGFEDbHZTwgpK4hWXSiL1
phJvq2U+WYy2SW4CirJvZy3pEtW6qoSjjQd0nrSbT7p/Fy+J16wNHzwPSpBKdQgb
2dznl0hXraKWFlis8wXj93+90lhV7dx7/C/Cm2cXxKndPpGr/gq/VBPxX+J3/S4o
dEVIT86atjTd/yLZH3+2cqKW4cCsScxk8r4m4sWhS2W2QtOztO2atmD5z/RJUNJr
V4Es/s7DJ9ilxKvc5KteQRsPI94wzY3yRlBYWu+Vxtu/qaeNpLeuxeTg/wdB/681
3F2iNNRfy3sg4cKGuKL3EXZbpiH/xZTwBbIv7/eJSEXXyLYxBCfBeK5R6r+qlh0s
brDcmhWFBA3qP9GtaDrvHB1Ft/mZNVA1And64kIsxOLYPb5e9dTmk6/JO+by/Ifj
Zrfs6IyaKwmAA+mrjlUpvK5rcPmSugctp1AVw6Z/D0KAjLXnCTlB3t38lr77Ilra
75D9aILC0eaaXZXw3ecjU633PmHGIwiCX7/pkvCYGismN9QMZaqQWEZYqPedKoxY
hVOKIhiria5dfZXTfQgJV0zO3r6mr1+USGmGnqnUq5w8PSrS6+BlkQpDldxmVX4B
J1wtf23HSc6aRQGIK2BJ4TR70XQQp2PvAfDG7lpIyp1+HcP1yNgEsaxnFFfwdQFU
KofN6D5I40XUtBKCCGoa2iKeFpfo8swJ5Yy3lEQXpsfU8Z/PMgWxvYK21eJowZgh
WwNp49+BaTipgvBLzUEIFjT9FaqdH3yuB2o9fc5ZRUKw27IA5bDjFW2z0t32R5/X
Of6BJo7Ogq7tyAVSACi44nN/OerCMWKK9TYgoR+jQs0my4gD+ZUQvOwWidYs9bhS
vESjKn58chRDvMAZT/27sUgilhuSvkmrb9xzcsgBAqdkfvJaPtswYhsN0s+9dGmE
sOr6N2h3rlgA+yYLAo5x6ZL1sd5CA8R7OztFizljbZcLQj7Y6iP65g3pD2ySHZMF
YYh6gK4h/8yafPBs21tuw7tgoz7W9UFx7jX+4TJRHwxsrt1Yte1c1J8Lqu/yFEI/
s5dvQC+1UY7rlydlVkRFBRU0BEyTn4+tA0qCX9epJ5krKlzliyrTCi/kVhnXc54/
+07pPfQtcihfr9NQiRi5/zc4TLqp9zMKHkBpYs9wjmkuUAEUX1wSoQsVTzL8/LAS
pD5y1+Umec2H1wK9nZLEtmsoQetHcDQZF1rb3+NnhSp02znuYSAbhdy7a4iDYZtP
K0wUfyNQq8q9wjfhIB3cHtP8SI0TNPyM4zFvORtXcwklUc8r2rINEbTmZCiQTu9o
u39j368wnoX4D/Syjsx+9giWETBs/uJWNnOCTIaErcIJY8s9Bf34vQghSgi3BIqp
Z4VGODEHvQoSjwCI4rEEFRlhjxG/ybkXkLHYzVaGekwGNv8Lh/US+/mlFN9l4jG8
SS+4xfR7Cpz2PaMNy6BQ0pPflg1YtsKrznx1ig6b98Wu9B9mr19NyT75j8QTTvW6
crO8Nh92QCS4kG1+U9Z3AjDJ1FyjsJyjDFh86dkg8VyBit2l2mZ91sq4/LLTIQIT
O0OupnszQPsH7bCxdY/wxqsswnYWdVXbB4OhCUik2kPG2+/TNBiSsdrIkLzAtwv3
QycP167X+54yApgROF3NIA8Edyc5tVojNQzA/8Xa0R4pTdtbRjIzLTVurS/jp/Kt
OJ/BEsb/7PXR/NISZKVIbrYUVcWsCsETpOyeb/5ZMyuFK8bhxUQqj/ZrJu+qgBny
30EAFXf0Lz+UmCaH0hkkRz8YroL0LZ8amQBgmwtWBfLxvPUiq5btx6D6UHBC4h7T
Iakw6fMGSeS70mmGGpDq9rTg0t+9I+5Kt78kr34/v1xKccwXgCtLzl1Zb8peHi5O
HDIzPdowDWqW7tDjkqtef0dORdYteMc9QfNn32MRusKFhBzvq7GLDD+CddG75RDc
1rhAq0/UgWWEak70FwWlZkrbGkaRgm3yW78aOaNzOs6n7pWDxXc8B3kRyOfGAQEd
BwKLe2SwhgBGSLhDtAzjtSIQ82hLRa3JqIPNj7JAz52VUEhD9Famr5qEEp3wfhod
cAjk/Z7OMBQOg9p/ZBxoo8jnTjFFoj4/v+Z+nZrnG+lC4solsTKf1Pd63JcMGqfm
Gfi5Y6ukzCbAa3NbW96EvQiwLjJ1abrrVQiE265POoBNuOLHfgPjRoTc7Nm7G9eV
Z1Ieb1+VTUp4/sNfHMgIFYe0MWDCJaSZAoynK6MaUqaNYd/3fBjzuDIrWi1ltLM1
iYkH1oqDDl90FZzsKD2Z7RBIO3+C1N1w0J6eUxZHw9Orfl/bZBkRSRVBOVROC49l
67HziKB/AirY3SHogVUlV3bodIALxBITrCm6xUxJu46RXg6Qvw+29xsYb6iYH3+Y
e0o3BPofNpMp97JkqReU6WIHyo55tTHIEwIOz5AJiZ1Ga/M/CB4Eh3/fHKlMkktk
9NRPLjsd5Nnlq3DIf4kS04aHxS4gdIJTTGQwdUsMjEfT/HY0axUxfQzqp63ow6tU
f+IYEgpu1+HWJAsgoOIZ6mNSX0CfLjljERDp+pEz1eMXnqRLK/Z5sOHiJZ6o3wuq
HcydjBtm9u91X7gGanD1ki7JYoDP4J8z385bzy+72DTv0WoUZWA0XS3I6ngmMeFs
5sQOIDOgy8i3aKXHVpGcya1ODRQyZ8grejlEmbUhcJzsPbr9aQe8qVmsvemAQcYs
Z2ih2shAuXdM/UZpy3f20M6ZIV6VtC9AVX4LTTrrLGyAYHO4MySE5cJdVodPxdD4
IoFb1iaPlPY2WTQAB62ays1cGJBg7EdXORvgprN6qzVqHBNALD2Xig1sVjsu0WOR
uYIxDIWzbXJUd38Q7WI6KAEknl2kE94DO7PdWfh+QwshCWRJKBGt6MizPkmNDCs6
Ls1ZBeWJjnQ3Solg7Q/e+C114Bu0E9XAO1eSK3r7AekhSk6I41mrU0X/CGGhbt9K
TIIf8AGrIcRF9Y4EIIQjpbxLUeucxieFU4yJr6HFt+cnJ6rRZzU7jHpgjKRoJY1r
dp1Dbr781/87hzRZ8RP9QeLUL6CwgVuDFNfioUH7qydD1e6UIw++fNZ80lFF5yUd
fz89udAdQmseP1e8WJcw0GBqQOkMuXQF+TEiOanFWiMM9Qpq8MbxLGLAVGwL7LZ0
5i8mF410ecn8UzE97KkjN1QgKl4XQeecp7HIk7Kn4MAbBjrucVTwzmKhkLgADwFx
LmFEe6d7lEb94lDUtcnO+ZTIIweXx5BiMPU2nxujBYkOqZrkZvHOhf3XraN/h2mE
ypBJYVtd3V+3wnqZk/9dibMTsLCKU1pp8NLuSl+wcqaQfY5ZnV8Qu/MtComvWIEk
nJKl+OGbFJMmvgpFkHEUkz8JA8WB2RZXN+a2n5RwguW+eRUjOUnCZmKUzwDQHa/I
YD+m1354poGEckULhspn4QPq0W2xWEBppTSPW27HRjeWRhlE0UlnNch5ZND9qJJI
g5OWirKAruzjaDkF57n11DTfIMKqIBKikFEtMvQWUVmgKw0UAXUuD6MrtKO34V7L
qSvCr67951Xir52ZlAnnwFyQ7CnlKdXVWfdrGuL1TXeEY3NKE/cM2eO/k/itUqiq
MVJZLXEsl48fxL5n/w/C1i3wQRWHRRYkXA5tdqzQXN5TYv33pi31fJxy5UN6DnRX
B2PV9n566zmTZ9ZiUZLPQOPZyvqhLWMpL1vEJmuCCO2Oam7mOzmuFaz0dTbXnugy
qqx3F9XwuV4lWn9ZBjrPc4vr0nso2FMVIfrR/VD+6fux+zL8EM1j+gWyq2R5ffCZ
zFLLILx4AKiSj9tZNhuHIjJgVTxDkGna3bdPiCcBmovNbij0cpwmub9AmLecJO96
Axzvj1bRFPRqY6S0pp69C9C7J4m1TY7c5UdXWnRIfmSAv6B+NBln1svlYyHD3oVl
wAPG8c8sfQ3lkH++y1VNcGo7I+oRBdXETpjQSmiJ4fw9Peh0OcRChIjCnzpIJ6uD
3EbRSdASXt5oi7qdq4DosdhT7ae95ppFonX66fqwD6fCH9Z7+FRxw2ekAJa86fjx
BO8+KkCWnBRl4VjguPkQzTwW3/pnpqzbIdim5ciWpf6zay+IIKQdmL3gZJWqP3pr
Pp92+xx8EcZKAG/d2LPE7/ACf66jY57kJOGmtocwDiHoVxuhUV05QO5JUVBzMPu2
ts5WmsZSMSzu7MVEc/P/IVh0xORj771423xjwbOq9YBOLCHf+NTqFZxHUw6GcHZo
ozVgppLI6VlRzoRxcof21ql8gC3pP4/Y1pkEB8qXUNwcrUe11JyOenN/5WC+HSR+
hJaevruiG+l2sIfOB0djMhBA93uHPlz4dwwF9zhHD74QCYyGq7b9BaXyp2YfmMdL
QfJrCobU5HUgvgk6zzSw4fjVDxX8fx0RZoMMop0wiH32MRU+5OFTGgFGbH3nOtjv
uuZP84lcyswop+twuK7YqaRPggqU4h3L7sAjlnlL/o8ZuQcS6rD54hhDR28DAOoR
bikIIEgMf9Dt9kcdBq6OsqWiUVOMfztUIiOP8r3nOyRs9T+URGfjN/vP3OBE70Ru
HY58z7Yde6wssPoeBj9WSOTw+ie4n16QGILkkWWLhYDChV5XP+6xr7Y84zYWBNZP
7V8l8uYIPq8YQrK5gRrb4I97Dbi8bwCznHxYasV+om14zKplsPaqG+mv+2CCklvI
yEv/gbDZNDguzDuaRgk8GE8vz9pfEA8MENvd38H80zP3Gu44+tzOgy8l20L6gFOd
wsuGM+RXkesy0ShPu8OJ1LVzj/focbeJfMa7HP2cFlo6ultobPrZxOBVx1i31hrD
Y8KTXzythL5+jzPKoHynzTsG7i10FyEIEtV7S25ulC7iffHnG529Unq6ekvFLn+C
wiY+XR0XVHzoz69utjVuMs5KW4dU16jF56zdReJJkaTYh2zb8yEDKLk4E0Sre8lK
yynQZdoOkpvRT0S+58Qfg7+V4kfvmA6IucIBrU6kFSiQPVKx83S86YIl4L199NY9
dj9bs16PwuGjckojefBcQxUG7Bf16QjKiDMBXng48PRMynKSGFYiSLSG/rZr6ZzS
eSFrjU0z8/W50kw1MY5RUySgoWK/5pE7Qi8kfCigTbQ2eN1KybU1Vxc02aOGckA9
r3x1YyGCKDgzxjAYm3xHZbTBnSElThm187EnprlQC5+5QLI/bHK7tY1/knuLJWAs
yez8cQfT2x4JpUpOgIlBHZTM+Y/39ljyAH6IEdWgmBijclpS5sVtf11mAIeUOCvB
cNfao18ZJQ7YpGitenDxDcX3TSKuXJlUlQGkT39zCChQ6O5fTjSDi1hQH7m8+oTG
tomH+YX8Xl0OJpExfzoKWR5NtCEubiztkhcHDNVjKJ6H7KQbkrVy14HUAVvQXwQ0
5wp67j/clHVxLne8zzf6cDbJkJeIxdjO3ITk2yzQTYD8kndVlS735tZpxWNXRVT8
nEAk2HLm/Pj9MKE1WozdtovYdOWe/WL/M6Kgm/4OQbTt1xH8DItsn5fRZgGLuqqG
SjJujE+h1YNxkhau21H0ycbAeizCuZq/E7LTkrfO16txOAgSCgna5OAQ/ArCuoLf
ghBbLH0i28yTjsshZkgL6g1VR0jC0tBxeRTM6SALn1WAHKRVXjOgAxEvJc+XYZeA
lk+Hy7Px+IvVO+U1gQczw//IEPml81gazsGs6zv5ypKTtTIbZy/LNB39vjXwbKnL
wQgOeo67heqMh68qbbALRp5VdctaZMeChPXFSIpvGDTVKIQ9CHJBVloKrIFI2xBC
15mYeJxAmDsJByuu6SIUKlpspy8xbseRNUDW0ewRqy6BVG38AsGyQwIiNTlFoOQk
tdTYFboaszw0PEuxv+NHIhJz7z1SqLUAReYMZZLA3D2/ktsfwiHvbLp3+NkdEOux
Zj9gSR2Hf6xQw/53psimPANUP/sR+vwOtOrhiEC/RyBWWX8kRAueuHwpFXUFyYjx
mLs8t1QLoF1pi+4wPANiNTDSi4ONC/Iqdk2W+Mfo+gaz3vg/twnSBsUl3DMbzHNy
vI0Ro3CzCwe0fCNuCeLuFAtIGmsqG5NgE1SB02VyZOaa/JSTu0yAETC4Vdha4PgU
vve83tZ8gZFTYvCNNOIxNHsCfGc4OBQhEYCrv81uCl/MQrj+p/J0ywKxpIkEpAwS
1WutjjcUjjDhB2jtzb5E8+tjIzWdXZrAsEEGvG/PVh3izw8QcbzfHgSPmofmO4Km
6JbzY4qcoveJJdFWJZ6zT5GnkOAqZxjXzeB5zF1E8AaGjIbIJJbFdQtcKDePNtGS
5uIZ984GGKaco8Orgpfao9YwvcJeJlgfzwvg7YNIOiJvokSx3Pf/Qsh3M7fBA7Nh
LJ32hkr76V28FM9lJBZiutBitViXBb8ylUFX9VykrE53a9WmJkSfWAnWriBNoEg5
bugaReyiLuxcObQb664qdAWElUXXevJ/nzCzk7PYAZeWRw8n/2ANkQpcZlYqxmsS
i1c4iuPR2TpLiVk2s/fZz5JBUES76tobNMrNqLA9yP4vG/92UuTK3LS3JJB92sOl
uvzWH2WSxxy62KFa3zCCYdjRTLTVqiHTRcQSOQTEtF9QPXEahWYPOzSYUn4Rf7c/
m3Ow1GK+/ikQmczLXvgTN1nqsCAfc0b6SGnQOf3cVxae09GwPVmv3JO8tyIUF9Oo
i9kw5UZhCyuvClCzxHnWQJImK8RfP6bS0T2w5Il4jDTpOlAkMgzI8NI3BqnSVHaL
/aSaCUPA62oKQb+juMw2CMkLOmdb0OScSMmEbQ9GuEmm0nUtNIB6hJ0SoEzktr0x
Idt66oTm+fGxt4RZldrEA5e0sZqMa7ZC5GAJ9wvlOybY62t98uIhghAymuTTdDv1
xzQOsB/RbG3uug973Dl9s7pZFeQMmKocJsLzukTXi5ofyfumQkQI1Vnx2dkTezUs
Msxyc77fv9qkzzCBS1JlxShXRMiEhYoP49hXyZOJ0aaKBP3pcAaZB8iA+qb81LaL
58JusH6/xFFZBPfjpwpi+jjweMVNe8DzJlHmlIGAnP0MORgniYDiTgUleCcL35tz
/e2XpnBwG1q1TssyY/Rkn/VH8q4DSyR7bEVbuXJP1+RGZ1COtgFLmAUWstALPVCX
1DO84iQDZPftfuIEodEt6OHVd78YVfw9lJL1qElL7kE3ek7xf0eOoLVVgmSbpm4a
Xd3mn2QQ9ZKk8cuGiCVSB6bl0X0H6CiK7ia1KXmvjR59yeip1HzI8nWy4E2ub5+v
7vRWPdLEoZ+I1KAfFsUcF6dC6H+mTDdE+Gz86pOZ9/vWUJKNMwLoQevUCf+KnS47
LkIJtV2kOB7Emk7kcAo6BDqSXkYJhtJnXFyFhmMQpkpmFvzVp1gRkOY7F0/S2BvG
VEtqzJy8OL7+QWm00zBY/MmThFl+RsT4g7FUZv+CV776pUUqu/HFl5UCwbFH+Jow
fslX5I7o/gztHIdmqiavaUL5DV4XAf1LCYyQS9JxwMn+g/Sau6FUtpZz4GmRKaig
zHSeZEg+v06v2/ppiR5sMiOn5wS7Fg//gebZO6pHft4S5tgYdd5T1uzWdQ2lexuT
uV8Bh82VOiWjFawvshZ6+vVsQ9kUQWKGkXlM/bu6NXGmr+FJTZTb3p6ew5erDBMq
teF1xU837T++4XLVPBFOqDJfNcP+/Kr12UBH3cpOv/5NhGqwBFaiI/zn4pOxPL7s
/vPOd8I3XQJoxPrQZzKJ7mIMftZWx5/BclGQkWLZOQv1yRf7SPwjlm+cKdnc9l5H
+847SFB8uVNdOceHnqE1ejMZ4MKxZutFIT9GnpvECowNOXg64OW44ppCtS7xeAOO
hVulJZn2UxZ5Pswe8SpLbzrufgJGpALQcgT/v56/2tfVo13+GHMSv1z5sR3drzMY
UkI1as/K4GGaEpuBxy3zKmRPQu8y54GHOjclkv3BrRo+HzXy6LlXaxTcW16DFIzk
apsPZ5j36c+rBhBXBb8rKBPXeYwyHrNmLNsCYi+G16pDAAlzCXEk7+bYCfylmWQo
3kPEmWj5VwMT//YjFnii78xQP0JGB01FThLUJCbkBLnAkvXVlwdRFte5wf45caXr
IDGrBI+L35KHv04BbVL5P0uwx4w6CoIpQASCiaRi7zu70T1f4rW8PqlAVbjiqnMQ
z8W66yXnz1ty/P7gNXXlWLvcDxmgnS8/i/ytjUSa+rz2guq6GZqLrQ2fqVApS+9v
08n03rtQ53FIGkLhfwYnxYOskrApt6bxQ/HrR6DbVQU=
`pragma protect end_protected
