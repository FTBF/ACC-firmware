// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 03:56:36 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UjkXsqNcj+L5LN4Jlai82kNRjUD3346iGiCpscxe5NCs0Lg8x5OvSPGSqSYHCG65
DNum1Vq+wl1CUBJDK7ySHAAeNk8U9Q7HHarsmliU3rujoO16X93rV2JgL9PonQ2C
bbewLhTQPN/R81kpQ/eDPTh+6AEWM+0UFHuh5fxcVLQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12432)
hYvSUrvltlKE3TsSx1OobsWn448yPnAZXLIKU0Y0zyx290o/WNejjDDECohf8wuq
2vgS0mQeYzYCzBR8hnOEShAC0kPdqIkhC7S2vtkkTWw3GTMCeygILQp5E6YWJ6Lt
xdo6S4gCf3LkWyG/42l6DA5LaArPDjOOSD9TjC6I8E2ik/rSrFI08YsdctNJCe8t
BUErFLPARq5U87hixOHp1SdttfvLa5Ewx/K127smo+DeaE43lj72SzuPoqr1fP2v
FSpajJSxM+1YatF8xqrsemA7gPmGtbWJ69GxDIEDS2rJjhUGgrLhl1vfz7XuO8OK
NRoJcQYxx5+30Zi7souJ1Zw05NJ9OJiRN76RKGuQurtzQf+TohNObQWbIuNQxXvm
apgnTFvWlPmOAo099sqNEQFM71VXPQGrxMrtDyW7ur4nD9GUeCwhfySPBQlarvMe
LR0+hZ6cUBqmEvcGpgECg/25xv51n17dQWBpnPhDpJFwsY6dMOg7GX8kOsqwTQ/Q
XazDKkHMDJ+Bb8zkTuY4Rz07sfHdkppv9iwtG1lNnJ9fYKcjQgkr9D0XdBriEz+y
3hfVc2+2hTiryqGF0aseYq1Bpmn15FBqkeStW4VdxN/fdgjUIbP8l3cEVg1Zew26
GT3+IdDc650e/+im9bPIZUWrTKhKNsIc+6vsSfWv8U4fSmqrXWofb4loACmbVddj
Tzv+D3MWi6I5J9VBOAwiQmkoDnpB6GvYFFDhkQO42wAfUYUdou0QvmvxLvrq7OGX
mdk/uq73XIuPJjoFwtuaWWIhsto1/50dQCxqKyeHUi2B48yjKwVLYoFC0xrBRD7O
+9z6OXs+XF3J2djBOYYCE89uhCa/j51rdOIFFLjNH8tSsGLrNwX4tgXKBI/nT8gi
hFVQp30MTJuSceYq+zNHRQXuF/rrRbvDbIyFbAL3LyQ3xiKOwGF2rEnzq5QHZJNH
gMkqbU0vlfq+Nies/Ud1GiJw+qeva4HK20EiBaUxVsPBnRvqANkmB1OwI4lUAk5E
lqe4NfTWEpDbMOAi2gYhfF5zfA0P5FWzZkRrySIwlLzaPp4o/oOb7CH+W/y3YTyr
VZzKAWUa+17V8sTVeQGFmQ2FUjftgvQcAIzPAiHMG4yFx2jqn4EFcnNmZBqlqsDo
rxTr6VzYdN7ipANz5XOHmxrMfi/tk19Yoqso9eli7mm+6UisA5CkfqSxIVuzny+J
qraIss/Lasm+2knVYw3HtE4mY+MQYfgHMepVQi8mVPYlmhar1mlDvJug1gqeVWRU
AAJ6VLJYvuE9QMlvLcJKXlrJEfokuGPCXaXgt6lZ/7CmRfxVcZUNCZf/tlHQCY9S
jlF56Gk69KTWPASzSnUVYsJdgHOoWegYSyfznowJmxsOF12D0dRZxtfING0i02Gj
EAhfNT7SBvysFaaTiXVd5fKtwuCbISMI3P5hWTclMnom3zaHsXU7OLPQ27f9U2Hb
8Fhz9lg/H7YKYoMTZtPwL2ceDPx6wBBlFhqPYsXwiXhtddNSXtzNbLe3303tXqRT
0E+vLt7jIq7Kpa8uqu1Wnzv31Q1Sbr+QhjrB/HWsPU9e2/GpZ/PBD48XPsVLbDXF
JY5PsoQZynuFiu0bftl8xJN1603A9gAN1gfUIb7CnfzPKafA0CIFwx+vFo8IZLSH
PMygufTf2E4Nml9W7+Nf+90+QbJ74lireplqL/LgF7/N9vlrM9cKkGj1F/9PNNLo
jnInVuzL6iw6sBlmtr2+Ysq3rT7WS0Rfpi6AIYSrESG8DJK8aorVDFT5BYVvQaNP
S9vc+5gubrCKFuFO15E+yFXE/N7RMs1CosbbJ9FXJ4ldJgdAB51jLNnIS1kLlOWi
NrNwt2GX51nywoqNYjrfb8uu3iuMEFPO+K5b7WjJLHFQQ8UGtAY0kFXIhd+zzMIg
rbOVoRFUnI413oI5/u2Ov7DziUUKNkVwXxtGpV4M+E8AKuepoTBhqIjZcJNoiUlv
E2L4lj3tioaSQURrJ93YIgYnrkoxacR7c2lhMEpzE22vcPxsBg4IrAGzenBCJRH6
PooL3ewokN/xfUYT0QmIKo4Klk6vWpgBuhv1RX3mpIqNxkSrRNS+lSAnHPVXvopS
i5Ck1YBhZFcj4lU+RnPeQ3Cni1IB7TCati12iL/eEAxmj4Q43f28Nwv8TkflzVvG
6t4CJRAg8X0Kjt/OOIoaBpPggvENNcGS+CLF3CfQmVmpEjl6Tk9sto7fH68vMWeW
/5fhDN5K7nrwB94f1zqJU1O6gEj9xI10BtryAlH0sxGlBvFssAuhtpTXLR0RJFH5
fBq6EPrUat4nwpfSqN98F9RTR5QccWWsGYLS5gQfrwlZ6RW8ofQYvvQ9oUPhsnT7
otFtpSU+DdmCi1MqH88XzrAZh/gv7CNfFCdha0NnP442DyS886GQ3KKED7WGDpL7
tgJzQob0uBy+yApdLhh4cvbMQ6SxTQppmtFrRa/KyXDneq9D6rq71KXTUf7kw2xv
UI0If7tdm0A8mPZVhQLEslN8EWTFxULolrjHxvQqUfulUHPyNFs2zjIBRCn+4vvQ
zGMzS6tWzwj6uNCXRr8k3h0CoJSw7TQvSv4ZyIEzpcMgT+8stqpozDtk3AXT+A5l
4LmP5r45DcwmbPGkos6ZAGhGLxKmvwOWIdIKKwiydt5dySV9NsOePKApmHfizgH9
uFsX4+URluCwUmifZ5t8Ssg6yd6BwDM6/26cqTzD4qD64wpFmfmCpNKWfgGeE+7H
9SC7Pu/T+sOQwx381xFMXBOJwzsfHqhlZ3c6/9v666bn/NR/Xh6nO3g/0ik+Idrc
buMA9zOLIfOVyP/kBKKYgC7dVW0Wwa0raFpc844dyIXlusCw0s7mGw19xk7BqjWs
hHTuvINarXKzhMJANHycKYqItuq/iG10rP4GaPNvflf8iIADslFOB9zWQ5qnxhG2
70Xk6CkaRVbUrLjgWpmh4MlPAXAwOGztSegAxZyi2gbe4ILaf1qSAKtHAHVBiNVo
L0yPpGODDRukFH8Kfnq7ZN3f1dlOUysu2LFgtI+BZEM/wf5F+kDACLIBsN+os4l6
oorhvKssgwJx8BAHoAuIMOdBkXoxe4AfUkr0+1cJpztutM/RXUWWnDSmvwvjZjvq
C/xmYCbCOGdqnW6xs0efllFz0Tqyy34r/9p4X+idkbi/ne9FMYMEttqUdNx3/Ug6
AaKhOgyFWbGBEUSeKeM1X5Koerqp+BXpiGMJF0/t6VlsfZcPO92DqJkMacrjG8oe
58B7eLXe/Kjob/4D0MfSEEzD/tQ/8dkKeZbVlei053OhneBALQOPtp8YIeTbGhEv
5BPOUHCmwLh1UECy0KmeZadOjY+KqjO4e9+GLV9nM1s3/MX8YM20JxzS4zV9oPF3
9UxrgjuQo8vPxeppi/VXFX5EnohXD6pkU4ZdDYrlBJBeBIp7kehcORzF0siLWTWj
QSlv/h/LTKZ3JUQbPSncrtdzMAguB5UHTYRSEgkGtVjQy2KAqQjU2So+6vmGCPP5
IwFkcpzN/Q5WnlhnVqcIWuFaoYLvhUh64Yy/WVClBiUpvVshddyb1E9Ll29PTSX4
S8W2fB473RF9RR+VWQwAZLzuzMYOaS65F93YplouT62w/BTsvilXwjvX7NhrOiYf
Sg0w+Gc+MqxcKbx9hl7LXJ3rgzOy0fRLIK4zCxFiIt0lOXTl5kPdfA85kGpoAD+9
nahoccz0jlyFs1krze2D6w7N62kNodAS6j5n1xmhgHe4YLrZZVwemxgCwUzZQr8p
T55SnF2elnYY/eRSGH+z4/ox6cwYdikr46FDmaWkTrVlZTn4fxTVCu3wU31QRPCm
zZBMpMqvsakWno5PgYMBrFqTljq5JsUV0vGe3ZleLjb0HZnXawlLVFaJAYZvXgMa
Fccr+xHxB61az/ehnIwJmW8TsA2TnOtQTUMpnJutrrZveDHkG4lrZuPeglK6GYPa
0XR/i/uzDCzN+tEHaerWSDGZcQgVtse48ax3Px9FeaDUyjPQM0ZL9/FkE24A80p6
Uc2IeHkCBr7n4yanE3acwDi5kMXB+nUZnW3IFlpp7m6sbtUVutHpGUuLWqC97irY
F8wuIL9xbd+bWstxiEcVqJnCw5YK+47jVdZZEvMO/SfYItgvG6ylIlYWPBZQZ9eI
eQabInbsEvgifTHbCT7vaCQyGPFKSbQs0UqIOcH85orjMSfjVanEUGLGsofIQvw/
9aH/gdRtN7+rLsysL2bVaacNVW6P+jCeq13OgZRKWVpAuzRzkqVGyy4Usk9kLjyl
Wf6zr3Cm6NSLUHrxo8TTvO17QNJnV9irG1+Kn/dtMHrsnWzWpa2AbjCrRX2VVgbc
zoHZXVMJusa8GSaXgDOYrq9NeTO7xJme47ErNnjuQRQG6VehlTXL7iQC/Cy21ULl
Y4sZrdFD9wrUoht6kNiOnVQcXkzUyW2sHO+epnAZkAIczJ6TscU6uB+xrPZ/ut3W
HyMimwD7gdT5Wycp1LUGj33aLFzjLrr+nKxtUWejfcAxbYihvDMoy3bt21Q3Ih35
WAcUidXnHx+UK+clYFxWdqNz0zZqaVKZDnswpaiN4PuFMqaHyS6LbXvodPzzeiBP
ASuv5wAVHOPZKH1qt3gyyMhqjkxFy4COcpxNtYgAOs+4a9cOmYs5gfQDsh0Hije4
RvDBdqCQgDvXJ8s46y9Hm1KSX+aP8H/v1UJHzxe2DdTXOvN7hqnAPYxt37oDRFv2
jSDMB04ilIccc4E17OAaPz8r2lHvJMuPI2cYVw7frFVP/Uv1vV0zo8zBA2u7QbSr
gum1t2eBmHunxbyCMA7gwA8n+V2qqsjoti/gflFKjC9utqGJQ3fIjF79rqMDCzUP
WX9PK9iL1hpso6XL5lv0QiaqRlLGQZfjUi2Ek7T7chI0OtYRUfZPAsXvOZqFTOf/
TBiXKCIRINTb90T5AkRxNMwX8xzcASkmCQhM27lJq8McetPw9FAHK45iUB3b9kbb
CnQhkTcjpY3sO2e3iu2vE3Pm9v29xBj29W3K532qYa1Wru8HTEQ3kgEgrDMp/cC+
BJmi1SniqHrq1HcRVwcBK8s2mcCGqmKdkxhlWk3+hLHMy+nk0LvtC+y4On62du4+
2eMIiOAj8qoGkaq6Rgio0YwDodeylDfZZ/ai0c+C213hgq+xAI3XJF8oEhPRPXut
Hk3ntTEvDKd28EMmQz8r1F5FDDoa4unLdhV6zgCPK3wiC/oSmNQvAkqQhxdyI7dK
O5I+TjoRZiChcvzCRITCRquTYopVJiIZSnQB2b+5yeu6cbEX9LwqgQ7yiyWYWBDu
ze7os8ixmrgn4NmHpMDv+kJj/8doyfMu/lpGvKMZX5ZO+Pgmp6cSIefmWAQOK7yM
c4CYU0By1EuQT6GswEAh9sLwegEkFmgi41O5du4541dab1QuPtG3zAxhszLM9rek
gyjEOCyTZSjibiKT8sSkFdnYtW043FmcqZV4zKiVC5TZsajtDToLb7pRm7UBmQdz
0ca2IKgLc34C3wXXE8IFhTpxTctn+Ew15jNmX1fb6jrt6Se/i1tZ9B0gHENLwXyu
JEul2yhmI9+ZE9RkTb7TJtKVr59k2E4qTeIgdFYUECyMDcD2vdn7YtWwUJQd2DZR
9wm6DIeCxP28m+zQ29PnTvBqWLGaUr674kKAFrncNojOy2JrEIKjpnCvS47wIYQD
kKiF7AC/EXyk3BpfO2+JG+QkjHjACekjUUzerIEuYLsifmjsSghUZTZRPWUD02Dk
S77eREHxr5O9/YiUlr2S8NWkPVULoM7tzrxurjMoDUQHrvF2T4PAdRtcMVIoem9L
nTxrGwAlpRq9wbD0BmmHNWS3VyWkctTZMvHPldQSJdFBO7v+ndouhKpc8AX9Xarf
ebfSOPLlIOtRPHyPQiRzy14USSUNGxn5ECAuHVkc1Sm7OJWng3h5+BBgT6r7XezR
JPxiRYoru1lHBuLtYBrOdkwfZ/fxHJCK0JrBhKQkadbIrRFhY0gBOaBMEtAr3ZUR
3nGRAydk7q5+qufVjy7JCbN/B4xrMwKGe0t8dYPD9LoYWS6Wdy8aTRG1IE05G4XU
aX6yrEkCEHEPB9alzsp6ShpgBCQW32S9V4Y8FiIS+7fDrth/Oh2hTurqeZjoWzgk
sEk5lv5xbbwSZsCi6NCgFcOE6rAraEz02Ku9I8Mn3jPJcNaVNqrm3veOMtqeUl7i
HwDP9zitaXS1LEsFc041+cp9vUvqBxIGdjkvmYGAMiy5nR3pZv9YS6U23h3Wt0uj
hZyN+pZBqpTcbZFj+wjxbORopprP5yOkIv+Ff8SDauAKCwsrIiOmQTQEUkNTj+J7
DpMX32efqNkjEpsGzKpsjuK6U+/3QVLrZR73O0rfzLFKIiYVBuRZXWZRwZeYv1Ug
fc2jDwKn5vsgOYIVbuJCDlg0Tg0OR2r+zf+q8YBWSk2znnpyNH8A7vbNeSxCKUst
2PcwKoVbEiG4Vu3wGjE02Q0cegVC4Dhr5Zpj3NXbzoJPnCY23ERCIEgRJ0C0IQoz
QfYS000cmCrJczQ8dOuZp2xfdIPCFECEENjhctkjKoIioZLb0OQjsitWs626RGK1
VVISC4X/kJmLaRAN7spn//y2IIegYEvDklKVZlBbtqpBVgVEBH3J2icxcE+Hbede
a7/+n9YwtjGG/EqAWNHCcP3vvu+5DkobOYNh/hNWvjVb1t3fQiffWKm56NBHx4ji
D34saGLOQVH0D8+VYJ04RPh1Bo9ZhAExD4LluNkbv5VALs3LC+XxrUATkNtV4cN3
qh3wpmjRfNihyj2mQghpzhfk2BA1g8zrnyglgI/jVrI7814hDQmSkN0GX1mouBRb
bZQTx1xyBydFPLAEWkzjR3EIehQ3Ix+RhjVuIuaTgpst5WcewmaLioxd2g39VF5/
J6gBqmWR2Jcwj2qdBDqHuapZPEKWFMsYNv13jgaoIUa2V4ufvlb+E9cY7fHRjViL
o7bEreCS7/NL5lWEJr3oXuyZ9a3NnnmuJQDh0vZVTP7elhlEuAn7oCh3V/TelvsQ
FOCni9x621kEnB0QO3MW4MC9ndu4fy6yUbvurU0nwIvO52HRgDrjNtZaxwibxDx2
Shzj8cwWrt8/s5Jq8dTA2W/6+tZIN4DuBZBIx0nyysuwGIFbm9bzuHgwWpD7MeUk
COUvem9KPlwrYy955SZkvQ0sH7jP1poD4Hs1U62f6y2azf2+wHO0hWHwMU9NRMXU
xhKTT2uu5rdcPgAP9APeMArdWxpKqm7MBUW1+2Jus+1jsGVwGFup0LJ7NGf9qlA0
xZEKmjPxuPICstY9Ykv3HD5xxFX5vJZNr+JqHX1zOYI8wyY3a2ObcoG+fGr0nnsE
PoSCzuus935SUk69Mx4A6wC1Z9isGLaaWZgSV+yozeplASqBjPSsuQu/wWq+lvH0
YeqTFyVfHnZKfl4U0mIgw+vFBFLKYBO0aWivxoIwcZ+rK4Zc/OpKCcFgiJmcyzNg
9BSlZfnqlEOpcMu3YSN5OhMXv64I48TAG36b0t468cEcu3SFZireG/8WXlAf+2aM
WMZIlJs2pYh02oObPDemszAHcS9b3gXwuE+YWaoqTc+q0nG4Qeo6VBQsduCzysnT
KMh0fOsPXrac/oRkagPu1ZKouGR+TDLlJqnsuKXgsx7d5CX7/ZKDmQtImuXGzQib
iNPUf91dmZUEklkZ05/R0EypxCVN6VcuM3L8X3k5fJ/XEXOKiarJ33V8KyFOZYfB
WL3SMsFjSsKhQT0udKCpTis/4MhkbBxTn0JI6yjkX2JDxzOD+dSbh8InqNnNQ9JM
Hwnzi3Tcayk6vqxDt9vhQqNdlgFf8Oibt+ah49NOJFpDamWHU72LCDh/lWGDukSd
vZRUWRI151RizrxaDNg9mR3YLvTHEXfSSlpf1qZISyWImbmOwCaBaigXEh/cO1W1
pJ51qJoHVrIecy7y46PU3KFZhPCb4MT4H326Hu7ujkC07qhcWDhmaPtjlk+7S+C7
BXHTFm2H3D+u1P+dxiZjKVDsn8e0609kUtKbl+Uuk/3g/a/5SZXLIzaOM9TiPZ2e
TX4p0mVQWxweOPG6pBa47zHs5C0iZVpfzNOjlbFAyQPH26R1d8Vk8jLeTgCNOv53
ilfXrSSA4KdH9Nb2KTy3r7H0nMYsE8VvgQGkPvrAJbMTt1cNDqkYz7UUpAjhMMFW
JOF9YpgwSb/f9PJa3867ST0Roc1lm5rMTyqV85r5ut1vz946+1LKplxgC7kFJbde
q54kJtaubanfEbUl0DUYq+rlF/8z53goacshD80TI+WW0CKic474U7zDqKlhglt9
Y8eI8ZJMCJ926kXxa7FO/8UY8ZtRakGv9paGPloOJIvSnBCeMVvyRM+K/Zg1ozOw
3PSshWXaSfCRwb4ehsV8HJrdob+jJB7GXJI+X1s0XyCGFV86TBrHbVyH0sDBDUCg
zYPUPIixeFaa30KgsHx60LvPZ7gygYnRNu6iKeMJKAhWBjjVO9mHpz0dbAsxpWUw
sea1iF5a4rZslGbT201XOTvHeiIzGsfUALJGW75SAs/bxtZ7SDYfZo1/ltMFw8WN
aCkvvjPmgyx1Y5lzqRe9upkDtpaU/pAhlbty8GDX7a4cfU4rlyKScwYeE7TxLuoc
0euTSp7o0iid6tBsptC0HesJm7QftHXXCJWfdc6oxSmlW/lVF34FNAOczGamc3/k
P7zUEk3imMd1bvGXu2EbbIFyP7Mlm1YnZ8wBIdcF9UMtPiYlCFWWXyZLMVm6hNrI
Ppfe5JtOFxYKs9dNHA96DnwSEnPn9zyp4Gl6X804qsmrXuXsc69nEaph//uTwt7Y
1Va1YMmfGoyiwcyke7G29uK5KFI7cJwqtev6BTmse6ruSay3UyGuomF4lhTvzS53
gYnhpNj1spZSoD4PMcLej8MoS4VyQlSOWc1u/8WJ/0NOep7HLXGrQwu06HECv9wg
VtrQ5O5pxOCahHPICxt1lH98Q2srQmosZTQ68xTU03zPYvWOngwbVhsJZ+ru3Lnv
1LrROZZb3Y/mHwxrvhrvZI1+xIoeqsmLnsMQqzee44S2dkbr1XuyA9O1sAGV0pgD
FYVZ22ajyPZrWQCZiLowHpsbHvCk+mvDgbiiW5jItDXhuZmKckwssJMYfIh1WCkM
wFWLW7hQX0VyKX5aU7/0MK4uZ+ca/uTTKWg+rTDvv6X1gYCz3IVDtvuDv0U5azPj
7S73n9NGTiBFZP5fvM0/dhNRkDrRexUim1RA3nxvzFtvDY+8oG0sfu1z6p/sal7m
40F+x3N8hinca7Ao2vcLX/dXCCdb3GNtb5V7n6rAcoLd6b7KU2DO6IES0q9tevnX
WIhXwLdwtn82r2dfRpLPk1+Qn+ng6Mt8HkT50wJVxncCmUDMRaQtXCTx4IYBCmnv
pVhqyw1ubbEIBGW9vSfJtzORGnnpEPiknNeZwGGND2YR802ZtU71RkWuD20zruFz
kcKVBChZk0VAd+rHkNKQcEjvjyx/iLFgkXQv9k6ejBztHNwWn1hcPylvbpNJROm2
IzG3ngOjEBh97wremHAD4JJg5z/3ijQ0rOyn0OQuDJDZ1YyvphSMOLZD3rkE35Z/
V2zjpRqXXdMII1qo6Yw3uNPm4Drh9o7f68PcbFPiceOzN7i2HLwhExjjK5cVfjZs
dnSUF4zgjA8xsmq651QmDx1uvN2QamqO7cUHZHCWfdwSzDrpLgPdOwRg6ifCKhvY
3aOnKH+gaKBkzVy9ubUqgi8RCSfDB0qJiFBnwtwMN7sEMHEHq5o3/gYNJ7WIx8NY
YXhwVBtZJ/nISPLnWyAGVPGiKg+rzQ1d31o+BByeiz9IXcYtuP7P8OHnHMTEgdTz
KsGNjL+zY3su1Uj07a4NRsgsFFrd96H6ZJgKGM5A2qMaDYFNBieRM0bfGPXKNpgt
5JbuUWxOjt3qtGklGU+wMZuZhJB7L4rr2UYtcGF07qdHwa7wfge1Og2ZXn/WDjJw
OnxR41YupjrFzdTPveQCbavv4+8I3o7srIF4sGWDQzHMQ8k1r1W8k51US3KbYsnA
zlzqDLbUa7kJAP9jWy6zbMaFJSEMjgbRnymRlFwJXplnNC9TMZOy/SKBVmb+QNQf
na9QNx+nBEQdLVpk3iBnaWaurbtPITMQ9MgjafnEon70H9SivnKAuJrhNgGOpt11
QRvH3hpC6ZfYDRMPXo1pAaizlZVMcbH/FzaQ09Ettew2gZBFM0uKI4ORWPVwaZE0
LgDJshhj0+WyFfNDD5U1pHSsRZYz3GQzpSWu0RPSRc9BtD/20i+X6I05lznXs/x5
r1yycAzH2ikMJqf9MR7pBkgun+nKnzceH3trgRQoWUsxWCIJrvPVAI1F85YlAMHT
liC4xrUKnu1IlnBdxG0nW4Xu32PtvUxswxkgnQ8RQ7Z4c7BE9gIfhy67Ej3PLnSc
yo4RHt0WGF1gl4XJF2OVSZSOVcP4vZZRVAa9P/ufowdtE21J3FSgVqdOg0JS1ku5
yG3pRvJYgBlV2B1E/Ek3HOwrc1KDjSrT9OjYYPYW5+L7OkkUn948xsVkBEhW5sER
YJ+BLugxz43HH44TOjbgZQ5K/vPlf/ukh+PG0cfJutk7sP8bYCeU1VnoCxvtiBIC
XF3xdd0IWaElIk492raq4o7jK/tHE16e5aD87WEZdpN37VA9XrNZh66j9GwmfpV1
A7Do6hAtNjwSjBG9/0+xO3cm36dz0SMWUt8tlNBpYbCbnYLQgtTATWyyNzvDa+Ms
aT2uH1RQOT8ZHtsJsh3trJxiIFQ7j0jhASRXqwpBNe87pyXtzUGu5uiaPyBYMCXB
XvP8wuxuQONNRbrm//tOpWRAgwl7JMU/05xaJl04HHuxsth3Tv7JK2vdubYqgsRr
oThFlcwvPVSZChJMUjvvAi6CjhAKPtKRV1NzWS5TNwsV50ypafs0Je08Q4UA7WOw
NFa2pIVt96H1G+jVr6L1Fa9dUmie7QbXmwuIGMc6GgkCfPfnno/rojeisMw7vpdC
9FqQlYzxvWtHMCW0223utVX56WyDoHf9ya7XUC78wtzxXKVF9f0eifqNIdQ6eRsj
Mc7Qa5Yxg4TYD1hhqkuIN3xkGtQcKquKVMUUhOPMogOF06kmtEXvL2hdV8rDXUGQ
vfw65yZRCqLRe9Q21pZjbZRygz24Y/BlETPyEA+Js5M6jrlQAYjHPMNFK6rV5vI+
uZnBxM7vNos7MgvNC9jlo/ZFjqcjRN4mn+pZLSZfyl/ecHBlpTfUXUwODbvVOqyb
XCmK9dR4k+jdxf4ATvN3M6QVMF8JR/Jf7xBGC6a/7Ir5zzzbLaeB3KiwywmmPfcm
zHZDUeGpRQZQ9j/rz7JiXhNaoJCvDlex+Qw/6T4VqJW6x8lCta8C2YU4ce2mw4Tc
5/QdKGtvKPvSsNXU5qYnN6hJGRqHfMS23YjF3Gm2FJDZqMTdskWhjZxEP7XxHFK1
v9jaAa686OvGbfUFcUEMz8ADCyJkbZmHLOg+inyuUUzGyLRo+X6CaLE9BkGR3qAr
WTKFGzAPoJl4N8fllnf6xyOSLoFYC/Jogjw/LP2cO32VnBFpgG0l6YXZSkS7YQi2
pAGSDDadSn7Pc071xe4Rrt6KZlju6s2vrJ8TPj5h6JzvekVKx84SEHRlyffZ9dPw
QGjKGKiruXR5RnUMq/hcd9j6f6mt+sF5L8xMfAijzKRGadtYg/T4z1LPU9iNPpbD
P/4xcRtaPOctnxiEAa267a/8Yt3pkaL8CvTY27Yzv6ULVrsLaTdzFwDur2vgSlXw
IEMX9jTjyOftJu9M2VjhwuCo35r7pqhZmx2vtTUU3o0XGiF3z4Fkf9RvGQwBqGTh
+OfQDJe/8mmjZFPS4HOWsReeawwKTFMk1gJ0vLgcIdsuNDiAv9s61gtQl+vmegMf
sFkPqq4K3a1VfzoPr0mvKkFJdq7e4XMD1f+msEZAgV1FKNzljS37eZfKvOqozEI3
0Me2DKNald5yY1UXpY49c7KDgpiP0fH1KVsjvhCEmbnez/4h+W8mozxtNe1BEuq4
5I9FUTLucRB5P2i6lEA8YHznr/gnINpqlNUMQSSgM9ij+geRSPVfSR8SMWSud9H6
2yXyw/sS3c+lzk+na6DCvma8S6yEFa85tm9ViHJGqrWR9fM8R8J7WNTL9i+qBnVH
x87CwPw7Hy73olPTL9t4l6sRTBtG7C8ILK0cXylRmmTEDstqLY2NVm2y89NRl7EB
X/x5Hq/b2x8zxYkIUnrMd4Xr6SKLNb3VsGrR3zsNIQtw7mipgprvIVZD2utDdgkl
JaWjOaO88IBya8R7I40jm31+TteOpbXKVNA1iWCyyPqV0ZwvD5SLfUq0Tiu5hQOS
AE5Y3e3PDsFRe7pZ+5TS0ka6ovcLTzrMzPaLEEmuOKJcmaQLZEFiFWp/HvwJeJ2l
EIWMaW/YshGcDNxyM3vn9F5CxLs6EynVw8AxH+r77btrw84YNMz8CRsZPNDkofJf
ukyatAcs6qaIQxpfGPhP8v+1QIfA23voCKHKzqeOpEsvbPc30qLVfjuX00HSX5My
jDHk+HmsaocqcGZW4Ztp754o4JhdE9rVmqI/nOpoozUH7A5PxQ9z/2Qj1d52E/gg
8jUnOVMY28/AUafFFM0Yr0qAj2GcYBZGWcL4f3lvm6GMWhrlbusRxJRxeJrmeiSV
xqbx9IoLeARVfUBY/G+MrInIRZXU/MOnXplMLe+2oq7qFUmNjgwYVDCRb8u7I4p3
T3yXu5aGjZURP3NA4uMs8Ufzp8DAJTr1XC73oX0YvWqTBAhMdvf/oEI4RpEnFK01
5yIo4UA4yicklwxlT+Wy7Ubrf8In/WtmylPY1zIrJhZMpaX1sJjdmaDBjfabwEBZ
R4xbAdDHmAXP4keM2x0UF/MrWy9GEBxyR3siqTrrdMcKeJvi8sECyA5Ac+8X+lco
Uw/CeLmxQnq0InsKqQYjbv5xl2GASkZE5QD2BjHFxVVU/vEsGxDZix1aezWsTRAB
8BosNqCsstNTdvb9YR2yR+RAKeCeEwkzNmNv09hGtBZNag2avd631p+C0ri3e4QI
MhrRcYqHCeQdRxQw0j2VSUXSYj43CdyQvH/OT0UPqR3IXwjkV4fJUQPTWOM68JNH
SmCWshGeFFUAE81RdnUTayWmHjcQ9dD0HsLI7cYATbkgpi17GoqLLfJgmHr3kCaj
wWKrF+YqjXrEavug+QKAPTr3A/YRehXZVLOJr2zAyGwoGazux3P0FGrDxcW+mpL0
mv3qi5HAoajrmnZFoBnDVxJNwogPFOL4VANvki2gWAh6bN4eDrw7bkDW/3rok8gE
T9wChJBpZgT9CMA9EpZjbHcH83BTHtNjMI92xR+6WhsAHXzMiQkn8qn4vYAHx1bz
b/TYFWxosYtd6/VR/UT5TGYQvjrnGhPlM6G8/xxFwysYs7B7+6tYiiRuUld00naQ
DgAiHGTJHA0DPfSeAzIELNWNPYDiSyuMDonHe38RdgzJwoYJeSgtAY0nwfiisQ5/
Y11oLoK5KhLzfrXEVaoDAJ+2g3dpLrjj2T1BrPKNFMcbVWDuzVnQkdNESSSCaEM+
IU4RAN/qb0nKwvWTniIW/OanlS+89F+U3vpspN+bblc1DYAA8+/kBwqBiIfX7gF7
PzcM6cm287UWwebf1keNa1f8nzThe/l3OeabfQQuDXlKgLF0WEqNL+5pwlPBOJX/
oYzeU3DAOE+/iPOSZ9PrvfFOzveIwX0Eh2D2ROjjfQJWvBfvfG2X+74JdzNgM2wa
n5JB23u1d27UfvaB74iyGO0cC7z+9o1OCKaDv+zFnZ8alvLMAbIPpRaVxgnyGELt
Te17aWtaLtaJpi8eyoVxo4wJmUGM6ABs5pASIOKIn78RcQZEWHRIFNzCvd7ajDSd
nOHizG0bvq6vJzrw0QTK1xD93WdqaGZw2jc84bOpbh9g+foc8//yRBIH/pSSmJhQ
kTJp56uRVgCLMvbTM6DB+5tckzT3t8U6QEpsLkD8cwN5bYM2dE7mAOj1tgaQS5Y/
kUT1yWw1VmUpcDWoCr/7bFw7Sppw1BWV5G6Ex2M29E2KFURNYd61FA3ABiaNsYLJ
/JYnlprzukn8Km4dH3Iso9WIT6nj6dOgHGnYT0IOf9C42Sw3z1wkeqIczFNDhlW0
S2ynuW6vhKnkz0Co2yof+cTovk1jF71PdY53MhmeXeRJOY1aJHfh3xLGfJFwz2eS
1VsdZCXvK+3kThncXCrgdaHyof7Y46fK43TVe+1ZTzJXEahARaB5Y1p4AbXWnXWK
CKfSk2PBBvgkQsOU7Nn7dwnMkMHtOHjEAGwVkQ2vz3vAN2prkbY/BOiicCEkMoWZ
N53NlFbgT0k0IIMF9MAPSTlpSbVJxkg27r5fgQoMl4djhhvZzgVZLiFTon6Bx7Y2
NWhrU+XjZSzzqlsb+QumMXHI0OHjx3TdYMxKYy6sjxN2R2u3FaVSzv0QdEkoNveZ
BC/y+bCTiiXsirKX29dVr7o7o+9D4gYX6df6NflBej35RLsAHs4Rru4HMwsGPtbh
sk+Eazcf6HYkYnuJ1HLU3zB7+ueo4jaMStDyHonMbib5aXFZazPSx69AXm1SvCmw
M+aBJEReRjbuhJHBccoNsTGpf1bXxVYo8vuqwC7zuRiEdAV6oA1hQC+JVBr7fsCW
9gDeioXYYVwrFT6oO8+WG9Fq39+6vTuvHry1BxRT9wANxXhKqABab2P1oH2GImIb
RyZw+y0XByIyGyIO9M9HZbf3zjFICjlqiUa/meMRdoKfTQIPLS7dacG1WvkBtLnD
fgMYNscGyjfY4WmSMpIBqDho9sIQ22wCEwyfeHmMCd5EB1UIOO+UFocPSjLMPMvH
mUS9PKpj9uFUZpeE7L37/whB3Sh2lLxnWsdFKpqiC+/fotIL4TX6DzaoD+lkSHQo
lBbShTInO23mN6K5TzdSS0isxAjgXVG3BnmuOQj5tA5Cn+6Y4er4EDhrdsZm+EOu
r8Uv6gSAZOyzeWZXEBXwYUNTaCqiS0S6rrYBFD34Wp4oFAzOeswHsLNJupgqm1in
mDKfrfxMZph3oBjEQ+/62l1yMBCknciIAL+H5KQ8lfK49s1BiSspBB8usX3SK63i
WvSTL3tajBlmoDd2XSpbmsmGNYkgTYgzjIjVRSWZGa1vu1cjjaijUvPTVey7cCAb
uIFv0RVPoT/g2qr4IfHoc1+yyJ64ff1T+LS5ZM9sGXXa/o6mymR3y5FHSrWU/aC0
W5NqrNCYfnDcWng1djL2JtapRDbrRLM/oEl8vwpxUtYWNrx7d9ShThtId/XNsj1U
ujWycMUXgy14LlTws90E2IwxHXrPVUzyquPXVgHRIcwZlUrXFsCuTWT/+wZZuM39
JD8UGUXJXW1Mr2lq9X5Q9m6gD1tJeS6FHjoH/RFUL8Hbtz4NwoA0WhaI05frA489
FmgWDCuSTwT1iz2Be6Ki6mqEiXXWnWr3HpzA6pFb9JUbsQa29G9qAHDvYIRhbUvh
Lui4JcOKRLfo+Cy/d4gIAze/dwYv3D7U9Gvb7SyeHWzf4WrObsSUl5pTvq/r8hoL
IRFJZ0/rS8uSyZTkTSieK5P51ODr4DI2lBhNHUbYr7vlT7PHG7ri7QtyuvF5TWYl
3jlx6Fp19Er/x4IaHY9HJa6mQDtn/ysX9V3gPPlRPkjbggPkBxDveaS8Dl95cZVe
29fNJFThXb+djyPZGKquePAAv8sYgIUgG7O6ApfZ3pyE1cv3PV0LPKXTEXZ7GTcI
BlJrPU7XPaCljO3SGxNQuIlUR5q6KH9yUoECOwsHv1kFuli4a9QpzcQYGVGY5NbF
W1kn6t/MnFDAYvlAY2yfpEWeb/hfOIesHKMiCvtgF8ME/YzbyHxx576LyyoLnzGF
v0z6Yfd1MtCCmndkOgmanRf829+w34KFh22f0k1KQHXVJ5nfv65ZSvskN9RC/8Qm
u3R2SX2SQ/xo+BjB0ecKsB76U13owgGL2qKPZxiVlv+mCDJsmKb2RwV1x5DJ6xyn
3t10Gp4BBywC+ZxbY9lsyd2o2QrZrO46ZLISOC6qbvfRV/rPh7tHSQ3LK1Dgrs/H
PM9FpdAD/q9Rq9N8FX9/fYK4azhQ4td0yYuOoMgZpRYx2/mOFhoV1huuGxw3u9Ox
RNTs+2pj0Kya/OvdjG2/RLNEGec2lhKO0v+13jSqCfiBBN7FECVUyahjwWE11Y92
NY9zzEgz7wqmrCRKSgZZMWF87HXBZOHmhk8XrNtXWIMHxXxaPauu8txtOC/ZvnRs
+Lrvv94heYXnXvKUbJMjQSyaEFIPaBBzF3j66lznF79zdBRwceQFnC9SEit7XqZa
T+4vIO8ECj9YdRyehRQ/n3VdAr45643yazRFUZbgDz/62vo5ABA25P6v8I0Dgglr
PMDnTriEnQu8kOmIPLh2PKtG6ExFTsxjfECwUz3neFOCsHAxI7XsQEwV82oW7zEE
ZA+xNk6BUAgl4GH/RwbZ8k6ThuDdMRoJq3x81J7urbSI7npH7ZwSPN0k/L8nIE5n
RaPAew70f4Z+yieqUGWBfw/WTxIVksiSpKRqdwN/BwGohxUH/D5OQJY3SeRbpCQw
`pragma protect end_protected
