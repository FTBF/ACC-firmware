// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:39 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
iWEuDQPN5bRfzbpsLjphwVkU8qsOvE9IQrZWWdCABrtTK+KZRAZGY6+ZEJ44NdGN
ntPTLuIH0U8bRMKKUrZg4CK/JC9633ATGBxkMUCk/u+FmDLvZLu23YrWIy0aB1p4
jL4b13v5hJ4WkYrqJIY2h5+DoQ/ZD/XoJFBCCFffUm8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13568)
nJABt7LoIrSwFSkLFst9i1jLI1FXPehfDzp+sjoPSbPgrMInWhf6c6ROeFcypf5a
7mv1Bovd40Q+29aYDoEfJ4leBx1T+1GmdjijB63chHH++ycJi24usOJ0FFObxrGt
ibl+g4NQYanKfIweiVOFmh3kMRwc6Dd9N0ao3Ve/f5Ojx+EGF5NwpRjHX73h1QWp
Hh/4BJDhYzXBRq3Qe3dp4k8HB52LApxcFVxPv9YUkdOBQD0sWVHwsS5Z8hygizXm
kS6j54+mr9ukwD9DWiOa9DubSwrlhb2/vC8yId+VWlDVE8EAycTmZXuKfvK8Adqb
5u0H4UJaB5OC3aIxHF+D/psg98ws/J7rjCxHZ3OxCKLOdSCMWg0Msc9z1vKDZEFh
Vp8VuuwXJQhg18X7zWm9YRHQuBmVFhUerT0+aElz1J5jZMxpT1/s0WiT9Xpg4rSN
lsdHLZsaPSw5SzaetckbvdW1yJk7GijUMi2Z5TBv19GWe7zSPZhA+OD8hClK4oiJ
9p2tM31P6oFxEHjXKdlYRw9GkbEWkXNOEsBFHYeDUNdmUERJmjMBMOxSb08wAwAr
NBx9qXUIvXsx+bwsJb0osxu7Z0Jqbnfl4ckOBq49LnUBzjIPCjXUleS1Ip+7OOxB
PyyXdMFczQsRyJlJcy58IjfyAa28iRt/9u5Xy7sP0rNm6/yi8thQPckBBa8j5ADa
YvQ/t2I91lAiP1UPJ91rWhiV17zmtuVBB+9FmF+BDIjizvBw8jWKvPcNwwCyzS7E
ZkSFoa6kGjrHUXKR4lO6n7i2zKC8zCgzxDXKdCUHqkBOf+E54n12FP2bcXRsQ3Gm
npSMlJVkq4PMLljhGYfgE/l9MZTGJ5Q/ufJ+kizeUpLSmlbMLbKFLOjfC1j+3Thy
4XlJflhuyjGfKwUh3EwIEHJvG9RT6OupYF6bucTa4Q2qKqssyO8e1NVSmtGrLG9y
iGCRazeB7UKEeGwLowsiVQhxD2dqZeawxH1ZgN218Y6LJi6spQ8Gk8J96ZFLFcXJ
lgcFln436c5J71lG5O561aBA2WNBKPhIhFBylAtHqkQnGskJJSs8pDnGbxrCWq3H
rZhY/qmbCe5ZP8QNbXVPqDab66JnuTCFUYZSWzCR4xqBJiUCoZ2HuhEkiWJoJ6jC
Yt9Xmaz6T7vszEV24hRfH5+BT0xloElzW9s4TRtICKZsS8wC31W8wv0/WdSz4a1N
4mEqju2V9X8zS8sh2GuFcH8Rs64wcsoI+/8Fu5V9YcHTo+n7lobVFGsU2jQyZkHH
WpjiWYbJUD/w81TczE4toqMl8jDA7cYdRkF3epQDARzv3HbH03KW6TfUXio6QI3q
ByIi1PBD9CdeRYFwH0qLg2REed0GjtHCyJQmCESJ0OKWDlDpzhW6UF8kNsaVMPKV
gMHr7uvRmIyo3HoXcsHacTPGc4hz2WoYap+/8jtfxGM57wPACQcMzZakvt05/vkS
Y8aIDhkxA+fmtusLewxn+7uv3STuGuBP1eJcsa+JBbXfKM6RyaA7mCMQZ+1KZ7A+
Hj/SWdZD4TatigYogn5Tcsz64+Bt0S2m2oOEY3OiAlalOX4HJoRhUVwPDqnZC9Qa
QUQIzF4jgHr2yyYARx4nmnPahdYU2G0YVU0rI6viiQ4uE67L9tYTKWljbbSsu9Ez
UVv6SrXWVYzVLTxSVshLADZ77dGkS652t2vC9v7tTYR2dqiaBYGNW0JCzLw1UL7U
QFZw1POi+d/IK2SKmRNusRJoyDB7MIuRgZkf2obUaxki6LKSS9kp4xL/tUXEMU/O
NSu0c1FOVWJyQqxiplH8JmE/2cTiJ5RaQ9XpGgd1J3IJgMZiTLlgQW3WZ1/cxwQx
MxM7mHVvoB6okM5H2YsE+6Er7FwXoFNwKBYHF/yuNHTH2Nrqewjdo2amlnNCqfwu
bnZVz1qeAJxxsZoi1jaCUacivOlRvCI3WoOUMY99HVDWg45S/gnVZis3nSGeLyCe
ZengGIOyYe7078aWTBtY3Q9vFTorV+3bBAVswdczAA1YHF7yWNifq+ybMUrvYP2M
r7nBOSlinpd+7+l8/lrMqN5B3HzQ+lsxwkugclNbp2aS3YKo/x//sFlflvADLpSA
3ksc0pR8Ydk0f9PTJ88dmbLF9iXHOZvwWI4vFYUIluhUi3GMz+hBi/eD8I3cdwLE
85E9dk1bUjdg1iL+H7H5gMpIIYIJSkImVOw9OWYFKbQINSdA8Mh8Gy2O/BOAdLuw
8sDKj7W4BRVe9uQjNvjPkqpBWFohLXcoTlImcTbq1V3vJpulgObqdSoDq+Dw/dQB
HpbpxQG79fTM/868oHzyx1D+Lnc6TyGRZO9vcdoK6JN9BmRWw5Tl1yK5rjpGH9mG
SyvFE6EiqyXtddhFqnWqyKbR8PjFegVkHwkWI6WIYAm2y/npP7Su3rS9ZcRUYOou
tLQgOFibauU19PVhH/+5HjwUJ4K7sA2Sa+cBokgScxCi+i277jn6JdaNLw5R5uTD
2sbHwDBVFrUGp2tqxFwY7rFmsKbXSMcwJZPkTXhcFlUDEES42zdmuwmzfPnr029W
qIlqCuLUHppkH9+cgraanFCEmTfAgkyT8Qnn6liV6eiVjaJxvpJnvHVsz3IszNlD
Y6Ul/svrwZvxH0jWwcjGO7SEAnZMAdp18vhGrgU5QUAyRyHQ6xdjkOLBKkEU5nP5
cpboHDX/b/ZiOHomcyny4jZ8ktIgQnxACc6v87WzFL2xABJJprsDdNhKFj4R77Iw
oWwpyKAaDPUan7RmrDeQyXU93QbyBibk5lUrEg9A1WbKDS3EY9ro8MmoQ92ifCsb
6W//JC2VYsxoRF1Oel6MUA3rwDi6QMYJyxtFadmiJ7lf2xQ9D2ew+Me13vfqTzsT
V/RBCJ1gAeTQlRtn2Y19doJux4YfxVyJ405ECreHPyosQV56PQFlgTPwY26QWpeR
0wx3yJZp1UQfdUUXLYCU0qhBNt3A2XYN+20KgBrmxM7QRzls6x3BKc7iFUGlKfIm
4Bk5M9SKP8v86tZkjq0jT4nUsn3L3goSdJO8vkH/6dQ6JY7sIQeCPQiQ+5zhaNkY
L7kK2GLK0dugJ0kK5reiA80TufZCinOqQhLmuEccReELBp0YiNiPea9JaTGRtQyh
R9UqIPWmKQ8anSeVlOddDy12Rs4GpaV+WvN92HdANgwMfpD9PSdmwCEqckiDahto
fnAJm2LU0uVHrwjJbLvZw6k1prurp0PWqNkeln3SU/UWiQX+AImIT9Xw2/FhH+LK
Um9Z42eS25hc2bJNKsbi9DQj3/5mBtWgfUDrC4h84XIVUY5K5AAT0cyQWhbSvyp/
gBFkp6JBjUYkyI27kwAc66//or6RjqBEyP7klm6r1d5ZBmFI/21hHfGrOF/iWPbp
tbNe9w5UrF//1rjsQl7IRwBNc3bTDvg2gI8iCvzw2WNZ8ZFzTYnBNbh4vtn6qN8n
A4XYlkCvyNXsNDFTVU80qrt4ox7crwPwWf65iLiZ40KbPvuPGneo0lDpA9skA+0t
K4ZjVZ+oSE/IuMvrSpoGPaUqhWKVz+BUAlpixl93/H3iuwsnw/GW9g9QsaLLmdsD
FAszft845Bt5ugR4BqlwFqHH9QYHrqxEYjhhFmlgGthoMrkl2TI89TdcTQfKERaC
fJcm9XWuQARzcfw6nn8do6p3N2PTV01FIMXE0ZAon1fTjtoduAY35UMFGGlPkW+J
abBdtJ6TbBlJsoRRkFCp66L6LrB7v0pNdNes2l2euUX0Kcu8yagW60GzCPfLHB8w
VJZS7tmEB7P4KLwVE9O37AFyUCVm2CG5OojfgLmVvXzkRGSbtFOt2D3g6FpaMu+W
yU+uyGYC9ORUHGQe/KIvmxaRdFAGx6cHTcRpxjcBzcbU+vcBLHZRNYvQbyVn3sFY
LmvwtC9lGdqMCnueSGyiV93t+EU4FfEI76cJ/L5Z6uGpaq1oMymEERnkzvkou7U4
QsWyK0HDv1Susku0h58vXX24JNA3RLSjHaQFGd7MY99s8Tsl8iUywIHpYTR5BwsL
XlGSim/GxoFGC4DlCbVbN5FG5pIJBgTPRBt/wBffnVvvsmD3krjklLoS53TRALCN
r0EKvLH7NRPA6nHdtmX3yR9y1MNZbfczQ6tqgWu4aNXg+xQ+ALKziHZGUJdNHWCT
PROGT45HmfJigyC6iIu9x7KRq0s/eltVt/jEUakpWnU4xVT6dwKIv3RdHvbYSgg5
yFUlEHZTkrKbVT9K0rkTASMQv/6NtBQjBrQ9+WSBSSZtHDBi1pPjMqSYh/amoBUz
cqkiAmTdkhWqXBoMxpwBkCGLMaJ6/EuHgKqLBUbLL+ERtufCa8or2lp2W0aO/A8r
N4vbiacW1Fh5I2Y4Vy6mRZcmtNrz0mZ8ReGjxgZ7LIUObFbTyzLhcjyeNr2UPqVG
egJwlmSMy/PnhbNfZ0CmJGwqJKmzm5k19yDTQOBm+kpH/IFebq1sFzmf2rfX8E4W
snnKRshTbOGtGl83+H4STwnhPc7uf5izapyBcwQlcwKLYukG+hYkXC4sEoGN69e1
LRR+C6AiFckwj5D3bfm0+2wYjZcKSMYAV6y5BhmTfWQlQh5tX5ARAFpm/fPagnTW
oLUCRO0D8h3xsM+hkaoikUFeSo1ivVdRhKa6+UhjqK6ALYjHyjA/+iz691l1qNFc
h6ur3KgqyIgJCa31v/GGiN4/AXhcuXLCMg3TYj78s57ammZgrALU3namt5yxuMUn
HXQnUdEwn4VACGQBGDG6UZdV2OvsRfEyzGzpXCrUYcGb0cgtnFDD1qvgeNtx0Jws
niYRKkHtONchH3NQLGJqXEuXC71Xa8zBAt1hr/NT5UqRyBmK3kr09B2HHKvgW5cX
SbD62CZerhNwMjfj2LT4FJdLuGjp5kcCdISdHa8KsIbnop9KMdbmgvpLui75JRey
C9vBnTbrwJTGZu4r06iqaqUcI9qD7WMHONJaH7IFOumtRmwzabn486jfQK/s/CTO
w1j5QOg1i3OmcoqafoCH1RdM1VDLSZoetJE6YaQEc4ZbCeCgeeVIF0A4kGDedCIY
5Tr648j8dszko6dJi2cfskT5N8895vSvB4M8DGBpdEtfpSApDE+ZFGGaa0MZ9Xmb
HHtdHshgM6j6iD4PWH9u22rOmqvZaZ1OoLLTMyw3PN7JXk1m46Ssm4o2JBnwW5lE
drHQr5B8jsUFtIf14Obv3gGpWwcgNZK7UrA8VWMePXAvUOJxHR6QBw+kqJo4tvcj
hRQhRYz+qfn5R8PXX/wsh9a7ZWb5mozpN0Z2IBSU/XIM4yYwfObfF3utklOdPcuu
ze81SHr7xmuVCMMtFjuBcruXhpC46M7Q8Z0faElfJ0ua+txlXl7ePhL67LI5nFdl
YqBpHZaVNcOKL12qx51QJKfVmglmNj1bSPxoh80gA44VZk5LiDnkHyUo4/56mdwQ
sN9d1XIqHbRxX54juUmVCjzDT4kPqVQAapAyrl3ioGJ/lye1m2SmWAJ/KeT24qB1
TeQPwCHh5f7dVtT82NJVohP5yWLsCCCcIIWz2Xdmgz/KnoBJPhNPRgIHkdvk01FX
bx38gH6G8EisPcqv8fFEFyWDCXxitgNNXyPBudN1GwoLxZo2IG1ktm2/TeHENrte
Bvd1l2FKjBmGrFhQpAgc76j2Aa/D2H45q4+sXaYJUS0lEXRsSJUhc3W2/TorlALh
4SHEt3cRxMYbce67TEBAf/9S7DLUoieh881Qq0VRDxV5ZWfZP81hZesVoM/IpYxB
Pnehq1YsFWLW13r7AMLEbAI5rOvHJSYn4sJYMesXQgXR+tBXptJvUfhaSpm8sNM+
N47kowgU//1tHMFWkDI6W9aYizMzY9VUueB3QjgLYrn7jhZmMhGAkMhQiEjJvHRR
btHrlvnr4aZkschCSTlnbOJrYg74/lqAsKDPNRyqNxrKbHEqZ+CKNdR/3B61o+u/
VMEGYiiwo4UDTRRxE43JcUCF+4HpqcCcleYkgMniiOckIdm/F9CMnUp4PkfPLMzk
ohCkcfqbK6I1BYZv1V0rJ2vvR8RFEvNC8ZOYpXkOdRTqGWGfxAKm0ap0APRZndqF
zJVgiqVEjgdFhMsTzTa14xH0S0U8NWQRSjRfW8MF/7D6+XyoudU/43EncxblTQzq
cQpwO9WBYjj9JCAY35dWl7ELiiW1kCtRzFmpySe6IBHJONNMeC4zn0PvKRlIliYJ
p/18FfqdWGOSB1c9QrvtTZLAaNJkNwFzRVtMsWY8dEm2NO8Pgj+Ve9vaUV8n+s6Y
Iv+Y+k/rI/g1asTchNxKUEXVjKJG6dbQESEDe0x/lijJ5ivQTo8JJdJuxyqHE5AZ
FPpRxtzisSMKonhJgiuFmres6ROgyS1RgAYTOXcyITpbXLd+xKxsur2qKrwLEfgf
eIOCLmUnAqlCYDs14jBaPYBHe3KncC7jOPogX5TrdwVkDXPFxJ7D0+Ic7G54ZKl/
SlrYamfr1/C3o6J0vsV+WBOt9OvVuBGV9qy4YVWiJrmy3myeVeQGP5KqpNf2eBeA
/5hea+2c2NTqqkW7DAcbc4Q2vkchjTqIQb06/iCPesaz0OqTjHkGPK9QvpJt2H2s
qNQ7cW6mQyt7WOSqKMzYjUhJQrQuQZn8vJO3a3W/n2Qw/jWbblvlhyXu2sXlXVDq
J1v0A72CktYA6pO5Zh6CfXCnqx+6RxySrU/pNF25xKWqtBMJsroTIDrglF4uRUFU
TeD39rNf+DkctYauA6mdhvfcGIP0WfeZctd6lWat2Ho3QFh9cm4W11gbRkh1DspU
Sc/7e5hd9IU6pLZys7ATiSkdnQA02d3n5R6PKkWcI7AACmYk2+aRLMHJdTrKYm6L
HSXl7/3rat8f3gGlyJcnuQV3LWAMU7EWRC/+u2nQxswBMdnQ7oOt4MXmYmJLVNI2
awwfiumHJEJI8uhOXknTxc5SkU3rq8izm8n3vyYWd6GXQUZQCihQpvWaLIBETQfa
Ruilaf/o6ttj8cS/hjgu7lHckjCd62o0foCImdKq7Qv+GZNX9Cqk0Og12ngovUAW
KAJVZkg8flqAylcdOhl5wp3yCzC8l/pdmGbdRWimul+IWXay0pEKh+nydjivYLNQ
TGjLjiCGcXslDKnKqz9qyqxArOrMiZTiyTi8Jj/Yop+IA9ZThQtUtCPCzDLSYOwJ
tcb9kWZHbjjZUrQe/aqU31TifvMHCYpMp/DRMi51MfXwdrft/NWtmn1XsCyDxUBX
0gtZv2TbbJrtxrJkxxv5zUHBvsKgMu5Ad5Nv7R50XrT1mjTOSQ2bh8usnQoyVKsK
2nJ89nKfOhjTlJX4rsOIzE90so1Q5CPKhPI5ezgm/chmsYMScDQwp6njVX1RrDaQ
e3gqKooDgLTZh7ScRbNFiZVJXNwgFZqRD/GfZHWNffMBzoJ2wQHXrWW3xK/9aB+c
GL2BPbwXaoyhYpudxVV5j3blcWhKMFunImikndURYsRxfXfm/3nfSDsp5jY8sf5+
ZHNyJpXlRMxIgN2Vu0TYA8AbOoLw7kHm1YGQh0ugivTy6i1ltXvoW55BXiGyKhJh
yeGkFgI/k3GJhYU6hn6w+aO21KqZLROiuPT0aOqZm7AYYNfj7yMUlHZz6x1meaR5
UKyDHwoatMDy5QzHfpp/OM+4YFlJacnubiskALSnZLCesFl75IkF7i3QVXMXYi6v
p5ysAJFdSze50VfunD/KVvrU1Gfh8eL9Rl9+RkC4ikFoFAChBx/YYJJBbhpJRrW1
fFT/Ass2nC2YeK6QdaudODvwU1bcDME9wnsrsy/WCohoG1XfLIpsVHO004NPewDy
B6nIzRomj+vvuPBPVaUTUw9AYF+htOUB1FMd+SP3DBQi/BpcD7c0HE7eBzrDCQ31
K4xCM45uLn4QWGej21oiAdPwifoF7LEprEa0zjMqiMJtAoM5ALMbpApGqZdVezsU
nqr6Xi+ivPQVH1htojUF3CC2ziQUeboX5MaLp3G2x/KC2yJMw7l5rET/Xu0Z3SmF
INkypfo+a/31d71aLMTbypIiQ/hfYAV1kAUxQuMbpc5uGlhvg9KAueG3+8H6gngN
xF1bNPyVm04eMbqOV1wzNXIEq/GgLEnSkXBzy6xGCVV1txMktHua/BmknSvHuJJL
k6Q6aQ+Kw9FWy0qEIGWOuxVZSGVW4JN2WJ0GSgP+IPNjR4qvRaSwuDyy2ihGFDuD
Ii/4ma23uCQAZjcl7RqKY2y+BO7ozE/n2I+wYd8PDE6b+i/B4mg+tvmZUN01LXhT
qKVVT/qo3kI2ht3pA7fiEEZKiZyKm7GRIqq9/oNmDf008sZE/9hZMsXwWLpp4FX5
bIe35jIovIMvqwf9WavWzG8cZHohJyX5H8r8WnoIQbbHY2qJwDPD3DGhcFxd9LwD
EUi2XZ+0zI5QVzhjHn2h3DX++reRbSuADvwBs5rp5wv6ygObDGD8D2ZXdIKkdd4o
cHzvGLmqEtypCdkWiobf4wU3vw4OKFmqAVOEFMNllIZYKolZzEc+mVy0CYpVLqTq
Vi4CQe8SUq5G0d2EciHU4Z89K8eR0i2trPivpfa4CHrkfCpY2Xr6+pe4ncw+p3EK
mlBk1VRtPjkHsUMWkP4/HrRFvN6S3Ud1N/Amooje4nAwSR05tTxsQBlXqxxkYUR1
Fph+jTkZj64cG4cmoWvOEuwSAluim9teXsovB8CR4nWemhXZ048plWKRyzrHHCVo
uYH9uKjFhGNw1uTyMy3DjJk1Ol0lzP+7nf39v0O0/gDN0WjpGfYj2TeHqijn2YUn
oR5Qy3a97g5/aOWTIrXgoW1i/5J0DC3AOeHLj2AscRYHqyeLpftWD4xHKE6Od8vL
1u3/VIhSzkvPKWofSp3cDB4tEqh7YUQPw1H87Pa4V9tH7Zg80cLPvcyrp33Wld8M
O8YWZncv8kpBZkBNRlPe42FIHM7LLAnwJQLq8A+j3Uq2dgpd5F+67arMaidKjJxi
tLgK5/0aYulWx2m5BnQG4yUPX15/sXCJuBwH4aqK+Mj7YSSxgyROMKZ5udZsW8qe
+kf9xZvD1AnPKeibK3TUNvQ5346CEDyRIVLsUs7e4BbItX0OTNcX2hzNIPc0m4dH
p+yFijNadsgL6GSQohG/Ry1LMQC4YzMAkAlR+iOOlpC44T38/+LJMMq0+tAk8lCR
m10kQUbNweObeaRCrZtswAhFXGM7mpv5xCIWoYNhWmZO6MUhtjaZqNKAHz7UnHeN
c1WSnNeX+WSmeioLJgCBpSKlCUbV7NhIAoCxciK31QJDOKdfjdubcksTJw5O8dgS
mFPHW73bQw2/rPwq+0+Xo/PsVwLqN4R35+jgZReyaQlSUt+2A60PyvCLgC95Peks
32MwMAEA4+AYABcXGJwbTyw72JlydXwG2gkwAIK0vMRoYERCJgTgu1PDKRIbizFJ
g0djhrhrM/dC2WjHSFKdeyvGQ+jz76Y9H9/vXIKwC4xuq1FgAe81jo8DTHHFEnia
oRmYnvIoZ3Tx6FQl5ucDP3e5tDJb+I9NEHEsO8WNy1Qn1iI25mUKnmwc0YWQxyph
ykFqvsAPOroD5lv6u791MylFNL+heHMD4F8w1MV059ButF1a5w7DIGrPd6hb1tnf
zhvASY7UucBRpHoJsLvnunrEAHOL3IGGEnFhedFxHsFiNqxy5rz3aag1pDQVkdhW
em/ZlESQkT496a5fMruvXm798aXeJg/23BSeB5r0uyX0cZ6fIaksGjACjNhmqstQ
Vx5CecBOLccV5Iqwoww9cL4dZj9wV32RVO00P+FpQ00ZWpT1ekqPfGfkblWTi05r
NDUBh4glf9b+w4YMyxugMhKI2aLN5ja+ZCnNSdZ8kO4w7IBjSsHVLlF3JcBpYdvb
ACqefG8GWtbbxL9dOorOMqhNjroO69nvxMonLXCxahZwrCfJ0Pq922muJURSAfLX
vr5MFHRrs2TMrki851ApVvltt4i/Y360lQu2X7mh0grqdAJdNOt301R3k6rQPov7
GFWo/KK48CydkJZhHQTpBYD36LesRD7dg6qCBKanpvjkrAKxm0y3Ol+Uzi/PW+g5
KlLi+KvC9k6Vax/nIlVf2OYuKUamZPK4IAOBawBNpboUCw8S6XN/p7C+0CDLUy/+
TcTyDSauhyevsxbhWohHlzAoKOC7LUdwXjJ7zXAbrIc3j1gNoYSI7i3M117DSJh6
ir8Y0aiX6gDK2xQf4hdzNanll3Gjd7sWjFtiY0ZoEFynwRG2u0kHFJpfAT21YRPj
naRV7anoJFcvUk/YeLUVtEzxIvtqtCeACHlfIyzE7hedOcPjEZtApD/AGWtawGjK
Sb3ltASRsPPp6quNhoTYyBOe6sL7gL2XKtfvGrjAPd//Hnx38rsAv0DVRE7hlseF
TNhiZYcynZuU7+zv40+/Yka+RghMtwcQ9eKWNu7py4e3nFzJEqDaNCaEpFq05caV
yaGnKw2strZlZe5Zh6zkvJIZHV0sTIEVR7vofbCP36rtola33ewM5rZIBZM/d+H5
m8dT1OVgZpiTXodTbve7QYwjPUlDhRXj1ty+W46oskNYqLF6AqgpNU00ar543C4u
Gxto4CrwNrNrbeodxCphmx3Sv0dngvni7MPalqFYipf3ZqDsYqzxy08PrAVtzbB1
UUsc+rdqb4Dn2xtsh7cn18mh8qGFawPYsdUidUBqDxhcf97RORoxxIyk0ZkJO4rQ
rYL5AdETDjY5ImRzvxCA0ThKnfbN8W3XSXA1oCJuj6wKOSWmtBlOBlt+sLyQOVQO
n1xJB3qJO3yeh9H9rCafAKzWP7iOoli15coC4HKyorb0FefvVHh+h5S14u2Z0+Dc
UlElkNrPn3TyhhvcDkQdohTgBuohsRwaR7J3uPsBbDgmPRXvkOmO4Ld6i3TmypRM
PS61YoJ66qrisr7uh/7GzdaiPQEZwsJaak/rsr5ARBv0cKzU6LsaymUQAWS//Wu8
mOeSWjM7ou5b/ZiB+tllSqTeNla95cCDMXBIjWFrV7AHzMPqImS18RYPb3Yv8GLn
hvRWd3EiLhJp1FEF0VQxZtkZSvEe67wo/1Gfh4EN4kBd9xatiwVX+RaVOZRSdzbu
zQeRcALm3qp+iAvQL63XlLzwRNNVnJT8NAA6aJigXfvk5vs4dWduNF7LqMrsosr4
aa7NM3OWmgOZtiy2XS7h+d9kJnEvq9inzXIHe8Q4AlxC2XK4MiUK1/ETf9oJs4fj
XxraKId0OX8fYURzcUEEdRD9hc0nlTNk7IfLJKOt3yZR8BaLIEPGJRHPWlOiLL/f
x2X+2OCg/WJ6EWf1MRbYde+5amf0Eshwm7T8KYFhgLy4Jusg4F0Lju/mnLpil0qD
IQVMC/zkNO8f8sjrns37ziQTqciyVrUP6dilkYxPcEy4RUfOaQSbPz48rSgojk1V
q6UrIwhUYzJbq+AKVb3dR8TYhtcu4jGPnQnPOEabyIevhKH4iHUXXXqcD6F/WzkI
3vAFnk8Lpmh5iufjO76a+vYzscSJtfQHUdImiWi+z5s1UDsp1sYP0+IVktzOt9rX
VElYbXZ10tHuXVHZ0h4Ntfc1jv57l4Dsuzapn57a3kH7C8zM6N6amERSsN4CaH1g
zqm5TQDPs4X7/W4ViAckdffpy2NvZLzK5twIGNMfdrNr8LJJQnNkZWe4Zv0zvvTL
acSlK2Gxpg8KktazPYmku8WyIq29Fg9eDW+tXi1xZ711yJQ5I0qmPD9HBSAMwlfS
83gXDFqbFc1FzT+Cn+gRgd++paEBPH+HVlq46Wc7Bt+YXkv1BNtK8BdOX3JHBcDH
+p+9rdUOkK1vZoaREo8Ny3pV7RTLNgvM7PqbGZc28n4PzhUqHyHOo+Kjc+//S3v7
DyY4JsOm10bqaqpAdLo8REfh84LkaYC8bhf/CpkbaNKMCeKztRcs56DZuK5Gahji
POpQBBnMCnu8JXkM7zn3UTk2LhgY6KB8WUSVM9Se54GgnMAeVGZtQjVeLSZgTZu9
dtgi+TvCDp6nnQzCn9/MT9VRrEOVDDPMlA+o9PQsA3GlAZJIB8Fs6MziYY04J56F
wpCVB2Y/PdzreE808IXEpvxvUi2ynn/njGdYF7uvrCZlMKlI6BNqdFuZ9lWE4svu
QNjZdx8rB8FpP9k0pX2E2NgpUOlbPb715pSCY7LJbIexXROxwN/fckJ7GwAOLHZC
a4YfelJVD5jWR6/D6v60L5rEuxchDmQtlw55YpkL9OIm4NEiPi4A4p2jZRxYPTlz
pwIAPfUWA8D7zU/ttayFQDCLZ9oOYPdrngQeyvM7cXFW4V9dNGBwXcuK7UX5OwLq
XycdOPPlv2erOgo/lCKo58S2KMS5CkrUcPZXcwI3DtgRUXqFf3VnVmpzLleaPIc8
g/zlNUMec4bQvTlme/3sEXVqMRIL9tcftyF1J2WKMr+LjNY7p2f4drB+C5riI/86
uJKDFgtAeAEATAUD2uH1QBmmbdQ3+SbqhrxkHMdjyx4eVcXyEpciSmHAYjZt/Rm5
aujLkHsIJBKCOpamv+Kf39dTfDELUvBQgqZHjGwHW+Pa8Kr8rrQnHYdpEurFMrhz
vRxJbONcK2RfNoBQYgxv7q95KtTAUeih4uEyQEp+P/PgQotdqvLgt0F+0YCxsCt7
356V31dvSmbkjNs0nQjZnSOg1dYruHLu3tgCHXm7jvi5cHdcaUMilvoUzzl6kDuO
LUYEcw+yoI8ncxNgbaVUwTJNPiRoAfg1eE90tHfFs+wN/sab9WAA0ZojWlYeQwzn
xp+Fu1Nyk7uahWzkOnKJKGJcnB+BicGjt20uI1/jKHh3uyg+xFXSfoAWBLFgmnI5
P9J96tLO6DNe35re+DEFo63qOLieBaXpVye12lnQG8xdxdSZAnU3D6y7anzOgjZV
HXHi2DrZY3lin5MyRRpu1DTk6T20Sv9BmBmOpvOoJ/na4ee/gKK3tXjnIIsnnLjo
0zX3e5dsXuHBQ1MXsoKK+3/s5ibNQNyn+vKiatw3Orx81dP8WBNCr6PPf0IxCwm8
7yJGEg3fkwM+ouCDvEXhUgAe3r6wg2heKR4WDFlY93En4MMJYiJVNVfNjH7VQRoi
of0jzt3OvQPZMjDPK0Hsjm0uCio8bUl+joYkTUxa7KjfnF8ZjVOkUZ1zdhD+ShtX
KB/J16arYFfceQmiNubtxBXpxvxOyjQSLuvz24T24rNrHf9plLNr7l5jj9ZAawZ6
u3i3KWRfWSkn5Qcxhq5gS9u+y/rzLtpQ97CcsB1nrrJFGUL6uT1CArG4sPaJYLQg
gzy4IQ2Vs1jbL2lxttrCy5TBEiSnX1sYNsvvUjTY5n47Oddz8N68vkIvY60yxjZZ
I2UzCgOOomqCQ0k3O+KtjYVUqTNE/iXs+924DUIj4oHFp1w0I5wyqlv4UZk+l3YC
WIFYZRkD7ANzleyaBxMJIf9Uh64UqNiftPfsxAuWk794YR9+uYQNrh4zwEx8TqT8
p/d3ocRqOaNTzeWiU3Os9pqVSU7sKCv966ivXhLjHEgS60BQZU7+hxGOhhsC4yKS
ilxZjMcVC6teqXzMyUmAuuNzHJyLzlq73bu2L67APRGGn57C7AF4KpFNCSehkkOY
b1LaYaeGJbU7JUQfd5/EkeS8Lmh0qkoMx2SHlyrzmMT6Q2NhdCxXmAlwLaz+/1dj
zqMrNHkA0/OJPFoJs4KA8Vwy8Q3Oy96xcf3N7yqB/WODvUpbEZM8q8bfHB3kBwMC
FroIvuv8hcBXTRhz2IBdJcYax15ruLVZod+tg0tUCoTSqv0TnoStHddfL8/H/Yyv
rTAiBurkQWt4/Ix4Rs1MJwikaDrkIHyBbGGEb2zeWF8EcK0+hJHzhcHMKeN42AXw
ePXFRXFazAYdYSKe2aG/oTymuT8aPvv+AElQjM4CIR2mk8SlUn0gGQEJl8XVoKFA
BDVnxOY6dUv0waVDXfJO4kX61CKRIU8NKeFz04N2qOqNnkM7njKVgxfABW20nUOc
F9HgDH1W/lu3DGXPIMCQlrfwZQYymlU1GFuaqMIGed2ltyPr9zRNMmYrSojKhEfb
fFq5jpRKVHzD5zhfp0baOoLP4vJd9mjEbmahzoOcQ3wukh6136ZiP3NaKLV0foTZ
V5FTFXbN0FSuxgka+ZDvrLlTNAd/Po+ga1I22sMegEwnVkoG8sNnUQTr01KTbSv0
QzU9JQ08NnlbqST5F1YuIqGLRlr+Rpt3qg+rM0W96Qq8RrxwHIRFZl/z/GuH79yj
/f115jiojEU31DkGi3bPAkMYVlhdQKEgVJjSyqEi3ulwbcXzNgBWw7GxMLALTy1x
UJue33+/uTXN0vMFu+TXj56k1kOjF9882XI320Yd0GnbZqHoNBqsbzDVb6wlzAWH
oB/yoLoM/h3PjkR2Deid9Hd06zSNB8I1y/pdzBzX+gvfp8lHzhiK4H2D1AU6RYzJ
qZ11aiqT+of5/JT0wBCRP2Q4D6wAdfGpLOxJb/wiDDh4c7JEeeecHB1l0tcYHf1k
FIOl++4RmvJU+cIHby2EO7Kot5opZ6icnMSKjXzFgImaFMAmokt5bFzXyYKKICPc
xJHJkTn9T61J7wX6g0r8vdp541uibm/JSl+JQUz4CHHClFVZaUC666G2rpkAthJj
l7HmjlGytNmDNjuc7o2uI0I7KcdxmNlvTUISz0kna+30I7SGQQQ2g4XFfpDKOkKa
ZKjm0uEV2kgKnH8ZXGIYkMh1IDw9CQZW3nwZidOiL+BXPP7wky5mM2s6wZUa+hia
SVCfb0rRvjeVzcr8UtSKkbIeDoYVx7mXZOrWwhktAcBDgY89DsdJYM7WgU1sBc9d
DorMN5xERj8irzChGQxEcRWhkQ8pBkjuEevxdr/Iw8uRLXFvX56LU0HJ1CducNQP
shih8scLjG61sKPehMu3tjaa8/Dq85JUXA4iB5ptEyD1JaH+fl89uI/irp47GaIG
yeCw9CGv721lSZl3GG/RvNpNPt8xPPQYl5ifT99Y5A6LfTgdhDnyO9dWsIYygPnT
yWeBC9mOT/W4Aou33nzqK61RCcPkloF7cPlyv0Gb61O8ZEK86LrjLwcdnUsLOb96
I60NFJofSudsEHl9WKl6YrCelBtWwtPs42MpjUb7CPyizMWTluIHoc+wq6taoryO
V24uO2t8FYj/TE1f6H1oOVZ7gBaq8MIA+qlINzv9yV8gZvZsifoS8sg/25cuA1qI
6sgO3e2V8pWjxKa/m+/coS2EcA2+u6qdPIYGuo8mOIVlw43rwW30dlIvObgJcaYM
5bnUlrjzhAsiJe7GUmYu1cwBauMCO95YslyY5/poM8F91W6uqBtI7T1n7FJFVUKE
DMDtxh9YJ+eYAfaHQ/VJTzYUbsoa6OQGQNb3KL4R1xgOecuzbTLFz51QRc678d8s
ahSN4y7XtiRhGzyJ72fAw+2WmZCJ3jy06CRSgHXlpk4i3PRjVPT0ZxpA1ot8n42p
wRAr9RxEXd/HmgIW46wUdIglCZaGDUZNztu1guF0K6dVd4CQr3oeVa0UeH6NxOs8
8HU4UXir3yxR4fwXUB6h8g6UULSzaG+gxT94Y3EA7tTC+2pddqSbnRU00xtqnQz/
ClPlD5GphKqvPgnSY9u51YBBL4+uNvGaRJaC24zLjzHeThvbpRM+/Mkd5qBJJDIW
38kmeD6hUkUCI9ydzWPDe8XYMfKxmXIDivh5gikx5kRQIwcL7SufpbnmyhlL8Uak
EzNA16Ts9Zt9I3/DMT/sZR1n6qMw3+sHZ6TvnrH13IbgX4uzLQbiEgzdjJucbwQ6
mtEh06SSyD/rTROqMVKFekJC/nN0erVJe9fSzjewgCXaMEVuoU+NQ4YKcEh9lfAt
IiMKE5OA167NilK67V1E5dISGyRyMSzn+UcBEVP1dlqRvuUDeoMip3P0eVyRFdnv
/0L9z65F6eva+7TeXWWfArXBOOGIkIKRW+BLuGYEL6Ag2ItvBr8YLB6jf53/HZaU
XqXzasSt5Z0RkCo9THchcZAyXo6JX6g+D4de/g/cHA/+W5rzbI5uVEEorggaUlZe
0X33OaEDg+YFtQ2areZnkroHiGu3gWsucNwe6jSFfu9mF8S2SeYvknHTQsFjE+rD
u94Kq0Dzs2vq+veSCA3xcUxCE+o3fhNLM9ak2wGyFL4ELT3CawWON3nvFm/Ebx2J
4+XCoIVM1ysapR7YpGswQdXEXZtNPu/7b9UUqfFDHv7f6TPkvLaIdBeXJUuyuJdg
cEy2HNDvHUIAO0VU+3+G037FabE5z7FI8zRqK3ZREIJOdcPlXvWM5dRORyVnkLfN
d78m7jjgAmLQlWzF+bWNqRq8CoGxAOIF3/fs2fMveZv3duEKa9PKq99VsjaO4uPX
uc/EOjfL+p530co6QDOYtnCJlLNi/W88o2nDEsbL2tCKBSEUJrrB6p5rbeO3dTeL
jwb+/ZxATUcGcsf6RMWmMYBqsalpRcvVeQ4rE6Owg9owpXICuemsX9YUCHA32NBT
/PPsys63X/akvwE7oTfA/3nJd3DCoSIz82v/aFywvjh9EGWw4Z7Pt/aDfhQQ1QXO
+x605YvXfxzUEX4Lj0XIPmK43vNB33DwEqv99gLZfCciMwmoSeXDtI0hIMFLtgHF
WeSz1Ac/t72HfKrYFV+hAXflhLnSIPZeQjJN+vg0Fd9isZAIVm+ee1ZhKmxvCE9G
LbDs23ljw/zSmF4hznoH4qgvdECEOHp5WeAI3thswXCmJIjrSrld7QunJ0foESpw
W6S5/pAqcSk6HLhU9+TH7x/WKZoQPs1JuOy7LUw5vHDvAj6lwvQP//aJ1LF6JGx2
fOe6J9g4uiyWgRNfWBZwy4g0ec4K+6gzBYQlFPbkDw6OtwoemZ0cysZTZRJKJhE+
f9BN5rMwbHdInIIEczqjLNEpdDknwnnvv6YiQtCdlRwzMwKePjIEAu58PIyTEh7v
qXOCaNDnjv/hYc4/8q6yZOQRfqeqPpjfZjFGyB9bgBeJRXge+X7exWFYpgrCjLrD
02E5+J3krxGymC4YX4c9xVZ/oelpgOjW4A3kjc2tqrY4nhsgOopm6a13cJkb0yFE
XN9ehPT9vpqEXrxRRKufvH3xZnWJHEtBcr6rGGHMDzO6+szuLy/8likePxaZgl3w
deK8+MqBUZgqoWXz1ocuNZcofNM7MlKWGrNbHIx+ox0SsQe5cd3Lq81jGR8qY+pR
p/wqX551hv2KMD5P1QOqguR/cx66t9IWOkCq5URF2EXRzWje469hLHsHyUDt+8ru
UBEW+VnXogjGkP+J46XqYKDOqF/U8rXQCWXGKCy6nO7Zz0B9a66TeCI+hwEKkmN3
OtFnG0qSVQ2p8s8SV+Re75WOw0f53SebZ+aTomcach5xsth2OsGAEimVBzNclbsp
/1gC4QP4g1fe+Xot8wBghK7tuHgdcV5JLIKXim++1KK8ZoyrLXxP31R4tL8DIiGP
3CS7lWABjyAftn9/LCOrPWepu8x4sqRHUskKt0vbO+gHvSg8GOAR+l2q9CYfrt5D
UehGIaLT5BKYzn0c912ZNZUHCxcUnT6CkHLE/82Wz6IBs4d3Zps7w/ITV/RiHDyO
Y69bRAIFIO4DN9mG/m1zdU0aFWyRoO9uqY1gIoa1wN9H8MMawCExI4ZcgaRPLuUa
3dx6odk9bslY24Nhg7SL5rrwTUlx6hGpIzTB4lHTAx9CFrE2QhI+alfYjKJ8m7wp
yFBpWMvB3oohMks06Ufqxat6agm0cS3NLIIbDzkwA4lT/kHlERoYqdSPhi+HXwJU
K3/08Iu2xJEt0LAdN0PRJV7u47aJnT05ZN46crcOMOKB5s7DukOjKGjggeUOyPml
gUV2nhhMWzK4coOfUtQz9GLq2Idx76fO+7mIF8ScWR2KWEvZ9zCBpK+H7k0O9xRT
t5bqycapcBdvwleL4ibv8GWGvJwc1mw5KVWysG9qt5OmKqmK49Yvai9g2niyxhwF
LbjHxr8MHZpYev/1M89MnTHzW+maZBvTVJRrq/anxSmL7TUlfvPR7zxKy7z8lH9D
2RQ96dYlW/PhBjzuEAHRLP2ETKA05ZbxfJdQi4m2B5Jkvxdlbv1LnJExtD+sqiMp
6rgbzMlmUHwkzmwmJW4GJBQE2kp1CexTQ2ddiEs5XRY=
`pragma protect end_protected
