// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 03:56:54 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mfpOTHmRO/WiWKQfdEcOHabVW2fTJ5KX/eGdjjaX1s3jZCFdihpI06OjjE0v9tKP
ZRzawKAeFUGet5c7YSYyBBfC9yJ5x1P+c6VBIsKiiOFX37J+JL+gvk5wFpS809YQ
Byn4LpzTUWVzSOJeREAW8CYnbzs0W9YYqExnlR1Xm+c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2272)
19fCA6YbldrzRKKyLrkiGSsbd/ORhvpBLUdo6bzaAeOvx5YBYKxlxrRQDyPL5AF3
EBSVkGmsabR5OXUnwMTIxXd8G0koLDoPVebq97Fn0K9DTVnspIkks8bgyZeiMLPc
SaQWUMkiZt4FQ6VSOA9N73fD1S+WYAyahvTirnlCmCVvTQkituhHllE9t7M8kWEM
MgWjvgZA9AWalhVdBswzV1/AXrQI1viTjY/FsvFsarq8UGI9raWFeOJBIH2xkRMA
kycwVkTRBNmMdvXbS/U5cQ7SPZYy+ShDTs5n8RkdlxBgXPDtZV0u9EvAueu50pgB
L9XmSh5alurDT3u7S8zz8CpclLlPQ5RgBdEIjRrNiinOvU5jUAPl0Q+ckwY1Yt0Y
0PXvn/c0v4KxDahKbljPFONWNcAdlXXT/TunQjid6tmeWA9ezhdlHYb1/ZLc3fiu
AYsO1hPux6XilPw9Q3fy6tOyaDwY2o6frGbfCAH/g5m343ectKXuEMT8S3714m15
BfG5RHSZsxY/sCI6YQwpRBMcfKZ0pLAWJ76u38OThfUyz4O/vVMZlb68X7Xh+WVl
+4T3aK4lFSerJB+iPu0KVlTWNlba0LIuCJK2fO4C9ds42fSAvPkBfhJ4vFj6Q1iv
ul9F9XiB0x/RYqDL/g9N8M2J1QP6Nf4mw6klUB/olYV9suW1PmZMB0TuUPIki/xV
+oAMGPWnxhSGuTVJJT6nwuwNm/Av+sdsX9jeyBQtefzxuJJ1eVQCIV0Ynrpw6vTo
/lZbCnny0RRVD1eAfSWTW4r8M7DZT77qLju+oPRAEMbPgeHBPvTrDriPcyj0zJQU
fDcD4F08X4gwNEg3cRKFI3/iVSrveIVEhX9xO6AnOXpbufKzwywFcx4ibtR9yH0R
n1VYTTUJKRdgnUoc+KGXLF3gXZmemrcufDCfCTmpFMBo1Ds8AWHgNtNsJYw6dqvS
q+rHQS+7McAJmkql+T4nuzROKT1/PxF7HOAOq9UGZzMmFXp12AK4Fc2EbKmZ5pB+
ovbdsxipZNkfwHgNN6fuAl3c3n5Cp22vWGIaZCKA+8zsWvgwsQfYbbZk342+iyCz
bZ94+5kN5koer+Bysk3cfxO8M1DeO2wk5uKRAgztlQPVgwsgEGNGV43wh78mDFyv
y8BEt+YGjJfMHQipjHSzQkD0qpK+EfbjCT3zCobOcUykcZaIArbdLCvMcwOe2PbZ
UBy98Lb/s+q8lDRBXF5lnP3jcPcOdB9/EajRwwXZ88SgsVH+e/+1wa2Sfkv7RtxI
+2Vm8ffrGkaVaB+DBlcwON1OIgPYay8M8tYkqoCTP+oYEUPbpp7iVDGxJSFgLcKd
kXrIDift/SDjME/18KlUzKKI6/efjT8jEwv9RhDLkHlr7S1lgQ/RbE/fDbaW5kp+
ad6SVQjRT9GsJY4zocfcF/QqG+H2DrGRqNflBLZ4q3F19XmSs09jQjzpkpa2JJH5
MuX+1vFr8tSG6FSv/eHU0ssy8SV0abTRdoEtfKy0jhIC/YBmHfmU+hAf4TgL37VG
5lF4fFUIxbDh7Be/5o6j4jNsoydrPA3qZ51R0IW1z9L5OMWbjUkN0mKm9bNT22ad
6aks2UHF9uSgYsTjcvE3r+MB0MPt/OhHnh3mGSuCdy7e4iKds1x9DGA87l6L5yWt
X32DyIUi3i05Md8U2aAqFLorsnPJ2vqUo9JuPIXqG7Y5H+hCA4SkGwkx+kD2xTsh
s14u7fcC468sTke4qKR6l7OYNkpf4wUsnjmMlU04wDQuCaIJfIGpsETaJQqChoTg
9AUnBJFGLQaOsdMewWXQ6q6RcZzSQjXNPlXNB7WQ3x1bQhUx0RlGLdmclWi9EWsY
9vwp+PfXyElBT2mLdXZQBz78qNOiPy0gM6diBXAqqnpMrrgpVyhkxrZtwNSxgOb6
cEo6VKyc6UKqXgE2KRzCQHqu7/6JmFzvAlrk8T9G0IkheUNiJIN61DzRJf9kOyfC
vSPvr1TZNugnmFoyUEQKeyfjtxdteF0vHmZaS2nngXswjYcU27xMLGNooT9sMImv
l0aD1WUovzTp65v1dYeYo1dnGj1zZi4bi9p8HG29yM2vTcT2HQhUuPd7Cr9rgzPg
JZog5Fy4BdFXkVP0TLm92VqBAipWHMCKofmJWshUDIzUspFtMNRI0TldNjYrInSm
6/69yGqkgB3THWqzQrBDZwe/ZHualRcaySd+r9gqNaM94QvEoIaBNbs26JvbPXq1
07XpfkfIfNNKiFwpJSALZA/UKTyr2KxGKxSaGjMhh0CSou7G0AIhqZkHpKL1y1wJ
EA7am8WZyZcslxjxWxp4kVPco89ZGnmhSg4l/bIALDkLgy/pgojAuDxdx1V4fhqM
UKxIAfqL0mhuQRus1lRwZhquE7XaOM0rwXHcnQ7N1KX2mZ1oMYWVO9y3dD/lfsY2
dZ9wUdaeTe0hRr9OdSTml3pXVRlzE0RIs0LWwQl94LMk1QNqJkJKVC/oq3VSvQgJ
ys0anVFald2+8N7QbTiasnEjMZvlZvuUooXr8Dx3bDgsnQueB3fk1vFWvx+hHXOa
+/e6y8GXqWUBlq3WzWd1XMJgwkUnmPa/pfFau/XOQ8d+XH9cLSNv5YGvMSVZ87nk
KDHvRjlSRLtyNQdJDWbDEr4gpkrnzMB27tODDFLvpphQ7ddp7ky4jd6iToWfuWJH
KGWgoFVANvP02Vdu/uHGD7NwSM+WAKN6dfJaK2nEmTs92e98/r+bJTXc2iZSlOtV
xBu/lrIT0iotjE7dBkMnjdk9jAp8u2cVutLT7n50slsLz+DUtgSjKxumNsyjuXID
z2SilX976JjAOSTVI3B44o0wX1cOpUT/34/JbvLuOvDw/EpDMmzrjdO06ZySx9di
UCgBeqIFvUKvlB1+SL/tJ2ik1rOblaXowvbxWXjC1KIjwNUeA6gNTceSabWxc1pX
GHgDQjWv4WQ5AKIlAo1jN3GaK4vusV7WwP0Ln9jsgXNE6i2X7wIGTw+5nH5jAjVF
eaVDhpDbpfLggKyjpDS2sQ==
`pragma protect end_protected
