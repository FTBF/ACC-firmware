// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 03:56:41 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UoGCgAIJPG1CJFHWgfuFAgssJIwDb0y8pDsy4O880WCRgKqtR/p1kpfkimXRVdIO
bVCeqHb7wlnNQCuwn/EOEDelY6zZBEa6JAV0e7zXPwArQ3GIXLeAlwdIvv/udGCB
hzmLD/8g0O0cjnbdI2BlmP51DNnrJEPLywBnCSIj5uc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7088)
BN6uMpjTkgb3Xq5wpEg6kSjDQZVq12R7/c3Es83z8e/DXJsDZgWs9v/hDh5OQApm
SNGg4E2HuCtYKq74IZIiaYF2PZiJX9l2lpRXrATZAcxbw7UQRmbCf31SpVO+xyIK
80ZedatbzeXX1Azemki8NG/X62IhGiQ2dYr8Ia1MXHIvkBsQEq47+luAskUdG8cb
+84mj20LBqVcQeaEMN8aISug0klAMH3tjtSiJkGsNGb79hacDa4aD7NAbTRcXYIB
gnwZPNVN7EVAWybWfaf/LB4jBvMOWoKRZSLdlyWwyzYaswQZDotCMzL2XUd0sMNY
53BqeOGNJegb2cO6z88GfzEVGxd2Gspzo4z2CkGd2agLHog23xFfCTqUI91eXhE/
p40BoW0baSX/St770vF1E+I0Q6S9bc/mplJqvE4yvc9Nip04e1RGTt06eHRiNjbg
50qSKfNnLwBuXSaA5jFBN2SUTfUrwnfARlQK/B7rQnPxYgOyR7L8MwBbJMzF0D7p
ee2UCybQ2BYvY7h9C0gWUR0+927JZmYSlaHgDD2EIgqzj9v1e5yjV5fsxjTXUtSf
hULcFjIIhNpOw/YYw3SxZeuQaEWfL/AmmtTlx36DiJRC956AeNLi6b3iLdW5YGZ/
FnOiHNOW7ZlQV71hdQLOblSKgbPlZwtqIIWvPgGd8pgr/imBdWhng0LLqE76QYMV
hk/jwm1fW8r6jhBi5ZTu1QvKq0fFuaYEvt0yZEOpS0cC7z0XxVVRBd0jWMdAVQLh
o0KJ0U7oDyQ25caLVhZM3aRWOFx5TvcHLMNAZCTwrLYW/hsDVlms7Fu/FLmidCyv
GbIpVEQo4nQfTLwbAmzJgDVGjNwT/hkyf5LylusmbNX6g1kSO1vknCuTshWTyzGn
FQTJkJBjgOB1naNTqq2IAOXu5p/ZoXUCulVBqapgF/Z+RHyvgZJTreD1MGk5Mheh
t2c2KaHJcelqlsrxltuu3OOZBqSri8XBbQmYvAYY/u58atE+XR/u2Swj8TJaxns4
WGEiDHnNtRX0Evj27ZQOna8i461ghZ6j6KBYt2r3On13XavNLFDYJv4W2dwymPqu
PGJmSt8tQi+5ZvOjtJzaC1nsb9JoqoXzEI4ZzZ3DScgLVcTtO24zTAL7I5VLt5Pg
T0FNpR1IxJBbK05LFpQiIhHgX0YIR/73nU38YDhgz9l7isP/aczaJqtwSsj7/J+k
iy9W0tQXenA7zNCMp0YLvEXMVUfjIm3LEavlPcutdAfYiEwGJ1tlNnKtuqzz4SnV
Q4XTePmAjiQulc4Iq5EfU6Z9vFPr2/PF78y6z3TbNc5ApZTMfyeInUhjuCbGtxDJ
yLDHGrMrLtcyaSwoSaNmGVaGDJJJLnxmczafLPLu6vNAeqUkeyyLtCmOeoh+z17C
J0sGGm6e9/03+M+I6LyFjecJkxQc70Xpqp14FZcEwTs+cTQpKJU9Z6Sb3N8UnZvX
ZQNT5wxAUoycIvFxOjrkCjmNLIqCQysdSq2TkQYnR1WgUaxrqFUircEXEx/6uE4p
W/UJbj1E1UxMuZIaQkA5fpvLxZnp9Qm8rluSB3N4VwpvDo3V95nMqpeb8YCS9RzT
PJ++opPxyJSQAUuzxepC3qobZMXSzEAuH6KaevaPbaPn1W79MyZOzbEkNtuLLgMB
0fZQ6RsgJN5hNDscoieOaHNQeDTq23+DlK1Yxppy5zTZmmkx0hDqGeIGOn8tbbAk
+6xwWkbziF/jQ6JvnCFgz79OEC9v0lkAKVW4dy5Nz4y/a6k0E9rh7n8mSA5SdxJ4
NOJhRMbt5LaifxIzqrUjtqSofig8d34Qh1MMArYK/h4QU+CilfNV/4TCFY0HvTqc
OIcKXQ5QvRaqoKubHPRC1Kfgh5vALk20XIIJlT8sL64lQKtag+/UH9GkOUhyem1h
UY8R8RMIbjInA+GC86By9uVfsyN3k1Dndg+ajxfAb2STKzwNIVDSafAMXl56089u
BlHFJr9/fTn6cU+oagzqE1/p+shCk7OPbZeEGX6vH1/o/ct4CJ+Khz6pSPtX/Cat
FFaiMDlwFo0gkBbX9XQra4t/11VZWrKwqAtyKB3hCxedjANgO/7DK3n8/tWpqRKT
9p6o44vmBIM9SGh+KrtV52B3S9EvZNCk+dgsCv8cbRg92Fb1X9VLTGlE/azmt4/Y
lbHs0RnLOSY92HQVKOMeH7ln+TH3SyHgQFI95I91Sq2dk1GvK64H9pm2H/BPDjdv
TlvpLbeBHksU2NFlr0TTnvT0Wc3MeZyiZ8tge7n2dATHOdDlsud1QTmxd90KCn++
W8Ak2BB0f9dw10PzWc6JOFqpInPgqC8ZIZjCBhu2RFvbS/Ooy+MqddNg4JJZ19aj
uFDBPsH/Bcq09otiD+3vaSn8qmyT5KlCQsC3d/Md80fA5F0TnQMkAxu0EzM+9pJp
GnPyZiOZBXM74kjPloifLu+K65ZB+PJT7D+qeqpO3D+HH/0EDmlL4OQR5Zofjflh
4M45lsn5zNkYYQ9pal7YlLqh8LYva8JcDz1dGCqKVUMNWThdI6M7XOfRhNm+RYRK
w7FwG8+OCH1x6lJgtHPXdeEDa/n+hn3KtmldXos5jmN8QtS3+cXTRE7muMJrvOsP
aVMydRs9vxvJ7cMjNrdDoiy2T2fnn9PZsaqmW5tjCaApNX+vFZJNBAGmq2BMR/MV
iRR6oQvzCZoO2cSrsFpVnn4LxgwKnFJTADNaXDa1Ti8YPr0c/Dvne2WDg1LBk0w8
dG+MjwJ0MMff2KuWXTb9Jc/i4Bo1JJw7TATg7bMJtS/0dXlBEQPCddqFHbGxeohr
B0/FR4da9akGyp79bjOVgkIXqRW8wPDzJNaeWeXoCsm5PBly9w2tStkK+Dq+jwq2
1jFjHT/vy1N0AGqgWkSLRAKZpvQiTT/dndyNhiXG0V8R7WWrRBbdNdstFxzMH//C
2OdiNIxWESPPjcAZMqV3aoMwhhyUWP4uD1kt1UziuJZPZjh/YDQ5m4wHcrPEudkU
M40QeXLrrI7k6OX9VD9xerPZmrMYKdmbh7OcHdQOGIFt5zwE6tKyDMIj8IASMlk8
wZX97tMJ2WsynalHzod14soIEnDpOo6L/yJNo+ExeZFu3B3S78WmY33h7joPq+zq
m893BC7uYyCivyaLEOPPDiyp8aVcyUu4wIBSoJ7+jJwdTsGTJ41z8QTsn94peEbZ
g0/UGAePasT4+CW/z1QQD+CxQZRzUHbw4KxN6FWcAqsr2xkFkltB5Pas8gfz/AeT
WtDQGH27jaOYxCBGWQ67qvDIUENsPGVfxTUC2a9n6UD4lwmdWLSpvfA50xib8amB
b7pr6ydwvZaEgR/4YPpZLOw3C6m0/S+qlR52AmSwBCIHP9r5DoLPGtcFbgTlpKyc
7gWYMbDYUsksFT/GuXd+e57wgPeRM3GFRPUI6XQOQ6HRk+7ohMYg9JIz885d52ab
muLgiX9yTxPrpdDlICI6YXqBJ17BLzaolc7zgWR9gXU6QZZk4+/weUK5DYR0Lq9W
80oQ66ksonDzOy7YLKw0NXtObQYyF9NQV52fo20SCEF32Mu8RC5kz8bkqeaWdZJY
f2Bi6FprdA785ANP2WECG8UD+43MoHiz2Yj+Dp9+RAwzfZvQX2ENNp1W70TSyIB1
cWNhNeWmZ3GUoj5WlGcVeLwYjvuQ4oXTcfHsiPQJj5n9AJ6U6xSxY/i12OvobBL6
nTgnpz9SsevPFWF9Yj3/+nh1K1DHvJieICTT48LZqPzRjhjz5S7w0Fwuoj3Cgack
9vlk6lGeO96+HWYsiIZn3SepDxqDr/q6rOoY0yYfDjn0kWB37S6zkw+PI7EAVVIt
X+Z29Mu18Kmw1wWYyV4nlcDlFuE4tBHmQcYhwyqoJQ17p1gCmo6+rZQLvinIIiqA
RcGhJIdxBJU0OoUSXBXYzYh+izVzz6ylJAipqSqxOfwVxdkptCtJQiY+G1ixB6oH
ok6RuSCS98cDA5ykw5T8t2NWwf6HQFUTDsOLAj/edRhwcWtWUspx7yRDBnxcbc5i
+JmHmnXv46gUVRWMj6dXYUv5RdsEz98JYK0sdup0qurEepUdr8v226Tsgk4DNMe1
OkPADXXi+W2hHomyoX3rzeJta89jyQGP9FKK5Zy4oztB12okEEBFvAMVvqD62Tze
a9P74ARqHoL7H09gpbPO0hWbY4R2Jt+v6tsdIKk9aWrqCoyyEiv/nP8NVIR+whbv
+gp0Bs7DGfmta7jV+2CCGEUtQko1i+2poKuHwty25AZDcGXDn8KC2RwfgeIaI0KV
mbseMoiqpx8mPkwvXifWoWGo3jcqZV0N4MDHObbcu5zJ5iAAFn1htDhpV68sb0fh
NsBoD5PV6mxbN6qTnhUjqzG77ObsNzlFZCxEi3oUlp5fxpJo5tEDSRRsmoEWmphz
E2fajz0jKP6LYmB0cN2CRVBYkLVPffLvU3S0xWnkZNk9jL8kxRt5LgC376SmBBV0
Ta2g3rIXdhDawTxgSa0b4hrDVwmpWha834Eh91s/ZOinWxLSRmspYE1n7Q4KZGIl
BDoHvSax73T5wzmNTH2KfTdqXxxnXLjNbhI6ABwYjUvRYrgu3NW4pgfet+DN4kg2
P3riDB0/UySZqQ4/757XjfJzHSp/MICAvTcUNC2BYx2dHpirPmdyxX5zoAt0WjuT
EAuowKgE55K+P0k0l5UN23k0nSTcbpTk5FAef+c3a9nOwjXWgQ5HNwsuTC5gXI+B
pg6mlWkflDbccbA9hzZNJ3CI57D9XOIUux8KRfjn7HTWnVWL7czJBeNyLHyEVFR8
3SyIVIKv1MP0C2VE5Wix6LDPQSSs5LMmj51blSrZfZCroGvhru/pvOLmgAkK6q+q
iJGhkKweZ0NNzywCVzDib9ToPKaSgRQF0SF913jgWvsVkO1BjeG5WriIRhJVC4dW
iDzPouDOktGS1u6rqQcp4U1/0u43qCIctV4NT+BQ270iGKOcPAzKxKd+s9/Wbhhd
Sx8P65s6l0FnY/j35HjHEN6zY8E0p7kOvy8omLFq7vzuyDC1HdGTKOKTzVDa4Wdr
Damj8zjvQ7LAJfnUg0/v5ETPzcfTjd8T+b44AAzqFS01uFNXEM5J0phgnm/zyGGg
pujvhzUB1lSjIfgT+TEWQ4u6c1A7TB8c8HyunzNMItWerqSFB8EOWqX5HKpPJhk1
o30IdKzeZNI2PeoIi586ntzrUi8VuO4oacMslXFrWvUBJLGSBrCNZVwickinGu86
nbBChOtWB7ofQOxANn7PAB9ee9Kdhu2p7MyRG+zo+qWmBM6tuOjgZZhvr6H3PtQx
P2b3uM11r9lm3+JozqwL728gwuGuf/nEdmB87mclActQPDX1KEQrvLC8o0exDQIK
BYkRk6TC2lUdRMYsqBaam5Zy5rxSXiULE7gI4/wR6bDtw2jfSCCS3ZCEU/rFmijU
jZRyCJW6h1NxUz02AkBxj9fPZQtG0pLJw5TKR1dssHaTiHXundEIso7JeCCpMiXo
8Ub6EMUfi1WMsbzHjzlYJYeLT/glA1iZzy5TlRjkC/fx6FtEPpAktVsszoyrIw5+
BAERvXuNZ43SnEcPjaVqa2BYXBXfQjAoBIywdRazVZQdsCJ/upVpffNtayCPckBe
VMBlO5DoiskD1OhR4kzRoUpfLwx5AGlu5i9ynSjfUnoe+oyomc5lOFNNayWisfnm
6/Bt1uoRnba4PzrfuLn97k/CUAZsmvj7m5YjCiq84i0HN6sCwNdI80NB+pjACR0O
RRULFpmv1RytPhlwqTsGxPk86ZmBP0m1E7S4JJoEMPo7YEXtnfnBM7MVmbA+3iAf
qodr4QL8O60FUd/aaIROVZaG/WdRpVkf8zk3QvtNnHHBoKcbxJjejOQeovCYvxl6
Z6TY5c2rN9vDa+aiaoclhbZROqSV4ruTr2LNESiWgdwBz+o748yU1mWLwbXC/4TT
seY7wbLs9oxuzzZfRXq3COnnSTsDRpX9ELS1V5g9i3GODqigsNNFDjucpLwzM2S3
YTuycD51OwO5YIt3Fh6gj6hhPPbt3dwjURHib08ZlkEtJZOKEEe6YxFHM6P+PiOZ
el76gTJRmeQ9hXChEnIQL5AFvc2cHXj8R74V5crODrBYuI3vvbiTTZbAIdmu6UHH
njkH0I7KH3Au6DgnAqhruFmgZTLm92GO4uj56mo4Fph84A1RyRPtYxT9MyhmYBz3
UPVTz0b9G8LgnZCjqtMJPNLGlSrwd5IvzoTNfh7JHH+Fz/cJNCJpXThpWe72SlrO
ob3XiESj+Sk8/BzaaYFMQ/gd370EP7Hs2iiwM8Me5iIq44S+GrUcPDMI0T0obRKK
6ZeFiF7POajPpaEnJJL53kc5KY53otOgopYtr7sDn6yt7Lnpq8s8fmvxf1/JhJhL
QAMT3ypWWQWeglAm77PASPsxpJm7WgnRY8wZR3RjGfoH9MiKqAodwXbmxa+7zFqH
Y7oNFMq1PL+Wheekj2QnAbieeI9SzvZagV0sfLDeAWGQ+topxUkUpE5D5l67rQdD
cHVJI7PcLYSsST/31YG08VhJyf1Lzu48WfSugKzZR+TZQ+7oMsG9mD40ZwXZXrHj
LGfawe0kxdrO7LI7IFgIpur9CuD+8bJCwzrp0pOhGtV4x++65oYqwJmKowLvjc/O
9DXxHwala2Dqcf49JWekHbZjYPrMV4r0OXrK8liutWahN7H8yegBBUqJOlAMtLaH
wLp7HRHpfdFfZjV2yof8NoLjBKvFTV9jQbTqyL7WW8cXOKPl8O1JxKUdC2llgFtd
+y0FX5J7zJoAtd320ubUzGdbvDuC/P2WRIMm03okDBHi7qHfglGl0r0oZe1uk7Rl
5ln9WPE6T8kJ7yTTEvOu4qu9iZZRsnPbG1XoLWMgSCgWFk4NljsTcdBa4KhEj7ts
ElZrSjPfJmK+F43mTCs2J4JCXIQIMw3em0sTstBwHT0uFWnxl4fhPXtjNPk0DfbQ
DKtfyBlB2QMuydCOhMEewEgwF55rWu67rUUgH7b5kL2mApXkL9C4BulcMmCT+Mui
zrDCnHcDFc85kfkWfT10wHE56Bvizwr2EYl/k+6q3hZ3z6fsLxRd6gkqA9XSBIzA
N27/UZGrRTF/GJTgF2WSeGrFoJoEsWn4gk9CUUDD9xsEPABxnD95wsqCiZmVcrJ5
HfdP1Yq6TzGOIrMgO9jwqNnKfi9USm+74EtQ8ITxHvZRlsEsPYQCa118xW+EANWm
srLSRVJu3eHPmioUkIIU5VFxeXUZF2pkA2688Yf3Kmo+cdycDbMtKGr+iYrF2Rp9
efXADuki7hq08nuEvs8QvZReP7fEgDvWuR+3GocteVg6bpCWNK/n+XJRSAm64Gva
ekLP1+fMb6n2v19ZcgZfn95c8pu1Y+VH1mQDJFtVus7/CKYHe2wuAX2aUtCMjQe4
BZJYiO6d5kqMBhV80Fm0uL7ezQsQV1kAo1mDyJz4vboDXIrJEeACl5098RGlYjqe
jcCJ8Mmbv7C/OMO/rhccyx/9BubLGBP9d4a5IhBeo7QTgIGQ1MHSHNUHNLtpgo3q
Qza5xDon/3JumUdLsUneutMBBJ5+FAvPgcuUrQrP7HhO4kq3HD1ynl9t+ZMKs2Dy
TAFPwXx/hyaV3vRQ320qO1FYhYXVLP/5eEsV1Wi+aqEr0ja3awSRoH0EDARoL/s/
Sf5q53NYBWsf3EJCj4s96Qo/UzlvtonJTHuNtpkSrX4xFlt1iTgq5pRf8HfaL8VZ
kwwvgeLVQfcGfSk2olgtPAoXR5y8EtRxDeAy9XyZ8+EBh5ibdun//4lbRzVPXQQl
tlG0XibCyg8+UmI5nMWzQ5czqTfxnoM4MGQ1D1PKGdii70XmL8DTejBry1ot1oNh
9EPZirdr68WY/Dk3Nkk+VyoitESYWjmHknVzMzyUKQxFedDfUhbo/A6AjFnRaX80
VYrXADmGvGseUGvZE68esbUHw9+7j1WyiHIHmQ5+9XS5tVynw9Nq2DNIUoYoEqrM
Ipn8IpXeLpWdqluw+S8tupfLFLNlM0k7XDgbWIXx55hx9fuXpCgitGcVx5a6i2Yx
+t5NjaiXWkthGjk09b+WLNPjth+klNr3bxKQ3uWTLkPAqdIKPa1Yh3MU1VEJ/J7J
ysITaZ1Sh3C/x2ur/KEf2gJOIVtb9jXJVJ7iAHkGap2qX5ELNB4RRaXgRH0RzXNi
her0mTvRq5NRF/iRdh9kXJiKeyoho0NCKRgR280n5fFTiMJT11nJO+CGu8BJ05aY
VxZ5zjYXV/Thx6zXbqi1HEQq4I/DTKgNiRX7Wrt9gYWGSKta4KoXoAogyUTuRi7+
o7of80qYmZiJ5WNYpaySySnaf2+5dAkzMfUbSwdNF5CGuJlfviKV6eVFQfE0WPds
Tof0VRkTT7HxnIg5adFVWQC25ixUM5LrxYF/MUFZVIXnNSggeUEO6RSKoMaU8nCC
MPa8qy6d7HcihOoeOgWRp1gbqfaF6kUN0PcwqqCj5kVKTZY930eNiLfSyeHRpIfW
nYumQSdaGno8lVA7HQSqfgPsz7CJWnkt00fMN+V4cCyQkXGDVB4UaC85VH02Rn/6
Bph/cKiOwkrwfzEtTytwXkm7cgQiWzJsRuVAUE8v5BkqhRmgVxzQUS2UxzYmv0NS
gKhV/YshUeseTf8ZAYnJfJXdUrybla6gZCPUNlZj+riKp1z/RAiVLj6+SxnmPCRP
HnsTSk1bmEPQ4e6r3uA/67BuJgNkExf1M1Klg8N5anJopZfJ5zPV0PW89jXsVV1T
Zs1x/eANPEfj0bpZPZ1nJEUXAwMQL7pLc026jsSTLE0dBKImi0r1m2COY1H5NXsh
cF8/8CNfC8alJHCSbytjMI9EAOoR5Ao7wSHwcdEgm1IGrEInopzBHaTUJrImVnCD
i3/WTn5mFRJJFkLNA3b63y56a9/bxc1OMqj0UgWmVlt6IcKSA0DXptF+Jx1J2UlV
AGD3RyVxzHV0x08TYdHaqLZu2eOSi4yfHP0DtDuCkRsMEF61DMfKSjH4G6g/b7kp
kZwnQZIvq5I5ESRH8ZuqUBt158m6i/gmakeQprcHjo9soRTSevUtlQuSwheyAz8k
ojdOtr9D86Yg6hHSst4zQUf3+EcceOP6R0GXB8TD1wKyomDkE/2J/GZQLwsZ6Xdx
w5yP0Z6kI7ihLeaAn6f/I4ntULAY6WlsIx8ccBgm8KBDtDxugesSICp5j1ANgigt
laakiC6mGE7CFJAGeroGEylJ4ui7nA1mN1wsmrbg0lI20hKvvzIOcmT2IP1n6/ef
bn3j5ceyAITh7/7soCaUmhsNykf+gcUjWvaxJndaDDUKQW/Ey552WmSdGkp6++NG
uViVMH6aA0wjGsShyRzairr2/VFhRviw+AWoqyXB1I5LKEv0CVNMDk8+g+qNkuoB
eN2qlh4JShN92mVbqkoawgp+CIESIQ88MnE6iP6TqLE=
`pragma protect end_protected
