// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 03:56:44 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cJjflmMZvIyS3w1/E3V5ODvEI3rqjw6xkk41ISvq8TlCQ+FMxDlWiLyrKTDhc0Hm
OgJx5+kEF1y+22NKIcu4Y5+uqyN8pakiiGp2pUi/8xFIdG3JwVaTYzWZF0rF9THg
wxgWNeq5US27T6ovJlhQDx5kZY+SFvt7IETecA3EMBE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3280)
0TrLYNCR/rUhfX8cTMR1K+4EnkijDmpVvxrVs/oz6q8piQPP34i8U6KPchkLQ3KX
A09UP5LLTieOvhC3NdB60YF4xCo/XAIPsjhcLwvpkIzIA6tqlMnQ1VEPcARhh4VU
Ad/LZC2udYanH0cCnAZAiTUaVVod9Cr0DKiOVP4c84uHr533BNJsOTB6bE7nluw2
Yv0/7jrhfr09VVp+5bsdMqBwqmQdgFGb6AQkkxoPH+wFWRGlfb0HZbbg/QoQJIlz
8pdnwBSlzYeOqgw3Qr4FbFLGstOdDvAZytxeBKdPnGLZKMxDJ7+WNm1lIKGBXup4
YnhFpbvg53T87wp9gHgAcqa9DKaasqD+D9f0BHiDrvTqp1zAZrhi/TI6YvqFkncQ
+CI5n6Lzk0ox6HaXwslpY/9OtdoX+yuso7DnkZo+5zzteDCQsYl5S/0anq4Lm9nK
P+esTp76a56EyAsofewbJFfpm/gW5W2r7nLJWdlMQB5HGWGiA3vSdJX1OyfspoDt
FR0StQd2Iq952THB+8DyZFGSztJdaCz6A96tgFkOawB1/FqAWEbECK64ABjxMlGy
0rK+2YsESEhsOVcC4iRQZEvmltj8A8Zp7bDfdfhRG53MbGhjUV46RlIAp7rK+g5J
ybdiujqRANwy9tfPUq82LPcAG3rZTGLlG7YDoGfue/n/Pz1an654krkKT8t9cGVy
Mku/NFr1kb3475KVFCooZdwVh3lYmFLuzFzomrJtZgWA4talU8MAvsuBelAvs6dV
MiVoc6vVoqRkEvBOWfszUmO3q7Z/Xm81sRzxa+KpTId33HhFzZivZwRTXDt6g1qP
a072ypEz5aqxLhcb37mIqFt0kYOLQH3DYxt2ZJYmRKlB1/gNJZ75R1euHZHbj34v
tDe8cvh1cs7agN0ZzXAlKK10Bk169Jloz6PEnc3VPWH3mcSk/xE28PesM+bbF4vB
QIIShZTna9c8REa4IFLRDJJikijHH5W0d+DknEyvNFOJdcZmrTkhevWvbOjzaRgi
o4L3FRYx4Nq0+kVJV8Obk651MI2YxZzUpi/FmYTyAE4WEdAZ5vMhvMX5EhYAYkNU
VV6xVfc6XVL3C9lblMm8onuUvPYsUOVKYJgkVNSNsgHjvFHfnPkxVyIrd6gKei1C
vP3eGONymSbyVpaIxnXZkOzvbbKkW+77Xv4ENs0NvL4tJjZT24hChJr43oVFAQqC
SuxRWP36YUrUCq4ksrMUuoYl5ibHhWTFNXeRau8MOBMBD2uDFVvVwDm+EjGgRcfq
Fviz6qXr9d1im90gFaK+pIYJozlpwVuCmUr08MsrjKTC+Qo4WsIpr+nPeOXiDKHd
oOZgJPvGyZqXa1YYRRtX6auBUWqtX4prs7uau8IKdNPNIRf7QrlQu5avCtfTnmHv
LbPeac10Uo1KUm2n3Jc2l/dYsrE9Br013kpeg5D93HYuMAjbMQZJhU3HG/B6pBC2
voCxxlDusb74I19Gx5Alo6Ep8g6CC+N6izjfAB9+qzAjXJKgu8EmbRViw5OzXQ0P
HxeVGYnSZ6GWninOQuy+hTkHeO6MbZHzzcGeD7H9J3Tbjp3+zlKn5iWzElh3AAow
qsB+xScLCAYBN9eW/pwnGNL/VEUmhpx1lUEY0Gp1Vvs6eAvNWCuMnS5JjtgVjGZn
KH+RMUKpsRipqFwuPf/dRhYYzF8FGbl4voP6xlcdU8pwGtW9TRd2V8uN3SHf3Rl0
xj8976EG6TGfIM522iudD8XablHZCg2o53ecRrmbnhFeMsqaEMv2JsBYv1grRX1P
3jAvbbYahoD8dhUYj+pi7sRZjbBLAZSYRphy4Olz4k+Iim7Qs0kRKsxH8C0fsxzi
qHKh5qDTCw/7CT0/22Cndt8IWB7mzzemMzMKr24SC8n5qUc9Z/NoUQeeqLNXdyim
H421FPW63jeVYeQJd5QW7MFbXNGPnH70zKX+sDVec968iGq09ulLCkg/TX0qaNSc
sUIY/XwqsEkrShdOXZ2FcJwRkULlo0StTfC9VNmAuy6EnnmQU1KUaXCuSkYchTY2
DchqW5Zf40cgZJ0v20u/WbKcymnCNPVN6M5PX7A5dnxR1i3Kks2ENQdMUcGebxXC
mK4/CgIrgtIlNztlYDL4ZEDR/vV0uUNW7IPrPZ5JGHvcKK3fGVSue/mXvd4jw2nA
7DomfK9BRg5scRhZQZPVlxVy0ooeUCHgrzgcMYgsGiWj6+4/xHQadfoYhW6auQmH
XdmlYYVc5hZ7JJaJhfqHlhfTlwKPvRo112pcQWoQZD6QOEnnm+fSHYDWoW7DSvr/
WvS3yJWg01+SZYbli/HAzJs1HiAHtMwo4abOVcWU7RfppmuxCVdZ1/dSQB9sCc4a
KETxCI2RXQZF35onWo16pDBzakmjpbxTy7mXUxrVqXkZbHrtSh9ttob1ph0XV3Ls
6QkcMzgwcd78usSVwCWQp7Z8mQns/vDY2D2fP5IU2FwTHIpuZqDDuekY3FShsiKj
faYFbEaj2KY0KXr045f9qwqRLTKUvE57O7zSVEqGE0kdIfwRpIRL9Gli2zYAQEik
+vd2DMA54co49eG9BAbqs1A1/mlQEvDbzhFtji7Sl7AqcaMA7rZ8uOiRCrfBRqSR
wlC/8BX8SKXNulxbWHUkPZZzcyTMpyJHEhQCrE53Cj3IK2dotBahFcTEaYYiaTk9
l3euNei19erRM67LXN/AHBSMDPku+Y3KB90rNzQJDWAGbF2vsio/0Hm6ac2RpGbq
vRuwaB0UQIaeh31vMoYYD22X9Xla5DdmBEfuTUWoIKBa0GbKn8pWMq+URQ17txtG
LjQL3Zwc8/kVBBpWWYmLt0eEdnKoazMLhp2/BJwUg0wJL4dFJpf5drsSCRSb3/NX
4iZtu+pIlN4/56hzhmenPf7Sw8C/bZswGVHmPlWB4lvliUKmBO2xCWWbkM15j26y
UQiOjYVc+BRavNYSLta60JRU9EHIFvxCSE+B+iU0NxADCwt56h6INV2SYVIqj8gx
EC2+3yo9WafB7JC47vZ591r7q+c8ywE8EmDnSO7dejnBOkoTD5FZqHxxHBwMgarx
Ct2Hp0XAyK7bRfTl2OrOmwrMX+5kOOB8keyt2k0LYy9Nq5LQe7Q8HRE/Qf9w776e
0SoGfFZRi8iZxtCB3x11lj9h3friUjNgdT2n+WmWAH+sAj15oXmt3DCVy6MJ8Gx7
YJ1TFuw573gmd+2o9l9Ybg+Lc4q3Qhhp0woBeQSblLSvDgidWJuo+Zoa1AGNdhKA
UiYmu61U9wdMbJ/usyDYJRSVaa2vi+mZBtw4FBasrathkrWaLF3lt6ahpbmk6f1u
v7jUXMgEtjydMWszDQvTCK1QalZhh9J/nr1qqpG1Mn6ovM1DNTNOZN9TMY8B7vdG
s05hmY8u7O+cA/OwdhIQRbGz9v2LumygqY9PxGecQpaIJTO3XymL3rV0ffvuA3LE
l+tLn3Pey9QjuW6oPCUkWi8mLxxlKd2O8MxP+wpUK0bweMvHVgqpZ9p4hpuW1ktP
Vnfj3jbnn8Xk4NkVnxRbo2UeUIIvDW5rgNTPtvHA3jul2JgrF0eLJmsml6Au3rfe
Bmh8aN/r93AQttO2y15ye4fGcSo/JJeM8ApFPCIds1yZadUmp7sWjn1SMTcEAMq0
mK9eauaPeJzjMUD5+OP+DNG9lpW0oKSO8aagJnFX83aJnrYA41I/NYz0uwwl9IxZ
YPc/ZwrYEYphnhop6V7tfwAk5BVTnbJ2bYSSnKWo2xbHk2+WSoKJx6caWqRKOSUj
oI4a7yLdj2ul4tP9IxkqmiOWBgL8UWQdGPwuk6E2qEUZ9+nVPVu54SmZSXSBQNYL
njXNw53Qz7AYT8UiyrJx6RoSX1AUe8UGILDvz7MoLiVIKXAUozP1Xo7+BsvFhWQd
2jCjnreRYkV9VG4wuiyw2iUxqS9D5l6kbV3vLLH1kAIdUyLtdyB5+XjFRs4Zo4i0
r3C9vdOHi18mBDDlXq5FWrEY0mHURENVYfa7lxEUJN8ax63FJ0rnEnOc4NYFpJ16
Ys7ktUhjvocfHUFCd7r1d0gJ/IYWPC3kN0IYjwMV3EAijMhcny2CF7nfelxrXtKU
lg4Dl8wOJLuoHwERvLYJE8yJVi2UgvSYoodz11vB8tttRfrFzBsFdOGhc+UILW2k
bCtOPN6Z8CsOPRYH50nEgExsAUVHq+wB1wygzKwnGOT5+DvHlxFKo1HtNju8A7et
Gb0sdJr/vYHj5geVdsLSqrjXB4xIUrBSozZocXfRqL7XJYWCRKqHsIjj7FHLbkWo
l915M7Taoc6ouNgE844gWTccc8q8MoL9BoMxbF79odx4z9eS7LBZ4chD7gQiO0F2
Wyou+DAyQ1f9AmgiiesDWQ==
`pragma protect end_protected
