// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:24 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MFcJoUDbBpSf5DJ/i0H1+h8pjqVgQb9fhnp37Up1eo7w+JQ3fmHS6UEjwG9o6v7/
pa/ZyOFbP+BZh4cDbcOLFNw5cYjCq+4uVMSt+AmNMy0frKbGbFmhBJsgouOu+1xV
9/aBqSFMps5/JLdNkhJpqC1u7SnY4NwIok+MaSOPsIs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5792)
YjgxYUvcMWbuLYCCYi5dYu0Ck7sf2TeFOXr1h4iYsNe7vncJ/XRa4dplS246G/24
P/u9hCmkmhgTc9I1VHjKXy8zhko/8ksNQvgWEeu9VcFtjj3rdHbHsjPGQbrXLSSs
e9NveNRFIKpc6EokDi2agHw+uf0VN99wM+AblyBkTDeFHYf0EM5beEe17mSxg4eU
b5aZsR5Q7Yg6F2QQlE/YgWXPouIXu6+S6nYE61g/IzNwSiQD4hXxOGdR1kPA1Udo
juBfog2SL3I7R9y3DRX8HrMRrgXN5XQ8XeHMDFHs/wqr6OXasvobdZxCKieVOTaQ
ifZSeHfGta4IrDoQp99G6Kcc5+l8hJdmlgRxeZcMJhK5h87e6JHOm1N6k5/gjo3h
sGVTraISyptJYR0LjO8/RHhslD3777+FcmZNWGcg0/XMhWs/mGEiWknT52Fbfjog
MGeVBeoPUneIC1LCjGU/81cZ4J0EKvRdaOKGl65Y2hcxrzlXV6EtBOOEiF1J9Lsk
R315jylyZPBFKkw2M8EfIecvwAHMWGhZjkK2hu4VZYgMQawlPu6hb2N9x9s4g9Nv
DMemL6NiimD2nK+MDPJUpiBUypN95v9Clcrt8UprjoqFo5NAi9sNQDS+Gim2phH8
TaTx8KBoifwAUmd2SnvQE0JVLs1K2DQQcDb6oCV9UX0yZOeNjOJUMOHW3uGnLkEQ
y7sruW6jcbUV/T7samdYGedR+s9caO171JXn98+WGG1OJbO941VOfHLIu4e2rGuQ
sRffiWtRf24+cgrSOTURAuwkyiTQ/cYCpLjGshoh19B5TkELrxO0UnhnGPCaFVoC
d0u50qpGxgAnz9W+j6p4zl74jCxptfRzqL4yG5Vgw4ZqVIg+Pioqc5NWf3PSzMza
kw2qQQnMbOTxMPed/jAprdDqkjyJovKbwp0Z7koyFjiZKiI6HJNmp66PSZre0RLn
fsOF7jEhIEI+DbqYsLVc65CcPzq8Vn613ZtxOzLXIMEVG4ZGVxFvkvCmjuFXWhe2
Se95fvYydl1gNd2CdxOOqU6xtcYCvn3t0x6T30q//vjq8yqhRTk4bSaCV1PWQL2W
Wfj78AJDgbjiYgU8p5qHfdjpKYzvom7ekmaRbPO4I5VinLR9QeiW/B5xfph7ShV6
74yj/yLp8/R0g6lU6/+1qLE7UOOgkQVcotae57OQKZpbY8BH3Xskl//DDDn6H3m0
g0z5yeHQEmEg6kB9naO3zfr/dDNMhGAF7vOXutkjP0FZwJDZrdt8ZeqTxqPjqmOt
S7iwLXXtXh0//fz+mVe4qsB8qoKO21hKKNu/wIRXzfXpskZGA1XO7KqEeiAQZEH1
ZALE3Or5XzjaB9nXAm3WSs5OPxrBfgPkbMbFBUzlGl/aX9gT7ZeQE9UwmrJF5udn
iQxt1XG82+Xjp0TIZYGQWxzSSIcXQqLDF1sYDRU5aWfU4TTWdRwC0KpCpnAELAKS
JupIV7xWxaEZauPz16Csc9GG8YKh6DYqkO/YcdX1OqpJ2GzWGu19YrrF2Px4oKXg
7vJ5tQ2R63p2VXwpW3ljxZcLtI46VcxSOLfaxru/322j8inF8Tq1+T8G20kLdl7o
mMtR+M+efgpr+RzXCksecY1oVmJIItX8SofNzOi5XTa53BZ8sUGVzKUlxu/ZoPM8
uuoz7x9re10FkagA5fRLyVsiRyenJuSjMidqGRwPqxe9SXOGdbf0YHn3Up90jHdP
tWxgyn09Uh9SMrte6Dk6Gnx5VllTJRdKQTF0eX6qgx/HKdmxdfAQt7SxArqt8M9M
IoC78Xblar63WQmOlgYZBhavm6/al8GYfmgyC1HJnTj4DbxjyunEOsc3Apn9b4UA
kHidENwxMO+AzeDik8FZp3+b1Lwloxp27KuYPNTEr1JGfD8cyYPHJohmvoE9rkkA
KBO1qwtDiYNPTEZtEMTh90bqR+CmH+cL5xeIHcbfmyTnw8GRlANmbpflcOlfdpH4
rc6MrjkfX7W6PUwe7rn0eyDLn1M5Qbd2oyFNBLb3FbvOC4XP6jpcNCtlgFh7b6td
3K6OWl6p9X2krALrjM3xP+PDKhxcz6cLvQvwL9f1WdP/eY/ZKULLMdRkO83uBf9y
5a1eOdMOPsRplU9ovnCww45MfZ2KUKPCvkesG4/oo/VHk07wisYNEfz3ufbalULc
FsRXW8UxXOwyAOjoyCJVjrJXNqhXfUg+Eo58iInVDSvRQFt8d7HTu2E3Qe1AyF3E
Cn0HG4Nxo293OHRXFNdEhrZFI51R0U1bLVb8545d6EnlaWH5eCquUlJVCS440xlu
IHD8clOgKxkZNwHKJewQympuloeLmXapklZhvoSv0ywRjwyt3qP62OF3U2pZzoII
d+8ayidrJkWOExXKxDIPbwVTrhWnQ4R9oqSwRijGuiug8QUZqnK9V/SYcIxhdIbi
e+VUe72WKtdg+t85gVApsTyNAUc7JDfswrixZ+KD9+APxa5Z3T/OziLtWREjvULN
HX2cvc14zODyoD15o5+7w2RbMe4ZJPde4Ku24luX6XYYS/gJg1zIA0bjwfaLHAfS
56tbQg/brquf9OPBFX5B2SrNJwGi5q12I7xTjMjHjO1H0AaK+jCb+ghLpIvTrKi1
Iv7NPM+rKhPRaIupyAh7YoxTEP5FyUy5yOlSGOt6qASBs7dkWQiWD9iksa/vcZd0
sicn2MNojsOjiiYtF9yW57nR4vHy/Gnpv9O9xNWLECGLPGeRzTt94/HNCg53CHt5
jXYHZpHpkZ2oO6yUMW/oJGxpVbcS4I/Ml6XBDK7ZkghfIe1sqWHNuSV95AELcnaD
ZNbj0EgCmxDwzvHXey7cmjNsmmSDSQkVSBpulmoTeGS4gS/BY2vyBDkqgcRlCz+S
vuaeDX3mrx1fJn6uGB4FtBvxDwwA921c9BQO6LTiKY36NfqRS5UqPzi4ugAMhRBO
+P/KG3+/uEWfVlThGnlPHdpYjFnnYc9IhDhWeF41EdtxyZO+EftUk671IyGJvMRV
YGIhtpgTHu7DZN+yIPCGdUO1SQ0Eh2OBDSZQ/YW2O/Ji265f7YVJOjAa0Nio9Wvp
DPOGb4Z3EWnhfIkOz05IfupStcbF1NraUfX+pfOSClGq1c8lOSBs4292o4nPqkA5
3Acr3KhVutfcY1XgrYFe/f5xn3f0nmFdfWg8IvuEmYJFJPihxq46Y0oxB86TnZNB
EThZt6Pvg9glnr7nSpnBRleDA88yaQ9ecTJ0dgCDeH9vpy2EHW+80Zi6iQuKruKj
IXkjHEjoZto2JXp2BrnVT5KsEnQHItv04c7ccN20yB35bfoeWDYYogbGYZDTEjlp
MK2ANRZ+kfZNtO8hdG/idat8MepEApoBgcCmAZRwnZSfbR7xLG98usd8AT0wcds8
+ELbSSGNgTSwAh5Z6AGcpuP4jPEAIdJTBP22meOG1lB5Lll8FGvVS+tpctPvHFa2
Y/uCqczS31xZI+mxvU1Yv1lFuh9IBUNRiwy1W8t1eQ/LVIbOTnLfLMh4+HsMcf3k
lgeOtDXZPuwzKq72nacoBJuPmFCaV+L8wb9oFF7uZU43uxlRdzk9v/lHXcr4pLph
oFy2GOUw2vlbMucEhKe7JNyJroiDMGs2E2c3kl4rRi2uqExrYrbL2N3G15ZUku2g
D8wgyrCf8lcr9LcWBB0t7+6uJc3Y063nZ+svRd6uVZNUoYj2Nii7EjCQJjBaPPdm
ND2bv1ziM6HzujoQ2GzxpPiPKMvU6lZlcgV8/xpbA924tqBaXtgDAG1i+oEkG6XL
R4U9V7B03c3fS1IcAyYWnVt74RQC9L/fJCRySAtCJG5JRRygotnAo0fF45N6LwSc
4ROBBimXCFXT9UJL5+vlix1Xh3APPcV1uGc9NAJBB3TTp9+kcObWNtk8awhn+30u
4QzLlMl8wutxBsRUotGtSNjnayqRJgp9ZitvwotBmQ0x5HV8ev4QAbfPhVgRKJ6u
2+l4QbzFyrUFg6BEO0I9AWXE3p+GNHtu5KS/uv60jHzDuI/FerpUNKCfrdT7tyi/
dNBt4XJq0xZjefeJByNVqaN44xPkHiOvb/6Z9+DdG5lmfRnkHCnJ9cxy5NiQbsjK
heheGN/8OmE4T+FQSkuG7Nu2vrZ4B3ELOO3ZONJ6tMl9TiSWOlOTD+4x4OQV/eMs
jr6H3fcugjYTdbW/w8fHmZej66bUfj6wl9PNFJ2RG4up6HwcYF3OYO07EX3faagE
TsXl9zPkk/pzzZuWU5eACAOWU+FziYHo7EYKKOliBBwRujzaIOkMwFcbKSd1BR1L
9UgZec6Nhs6iFgotCmZiDvVulb9365BM7QPrVe2n9W57ZNOabosSFj1PmE+IpRE7
J5bwuXeA3P0nlhPd88KTptCX/hXthozjCv8IyeILSCwzXxtJCdy0wG2Sb9s13cYU
bTXhksREgECyni29zpA+AHruAAEIvvJjvAWQnLOPrKnCW3zyZQci0xE/VFKBOviU
rrvKSeKIH3P32C7sMkXt1XVu/YqsTfQpA2DETFgW2QWWfYBHMYBURZcHzecx3JSb
hprSHsuTyBtBJRVxpNX0IqpmLtCZtgEmGTjMHO1qo8MYiV6zXYgYPs3yrAdnlICH
XMNNQK+bzR/8eHuPKdE6MNqIrgtK41eaHgD4NCR+gxAAW18abYXKBuPXzlndWNZk
3wkm8rU6cfM5KO5NPkh0x8GlNQKHVsmhPAVLKu6g5wFGbwwNMuJAIGK+E2mFKWuX
Uddw8BgNrKcM6yF30ZOaTwiy2JaHnUw6cWMN658igoQB1v1KppiFV3ZmV3jCHAxa
pqgNk9o2sIkMnIidDN3QWlCL+C9U/pHJ/6psLtd2xoexKErVLdSeTXZHyoH5tlFJ
xjJLFj3heRagoR+codhrcR1BbfDWRCrMGBxVz1UcU/sToatUSIKC8p+ahI3CGpRP
XuBkiZF+jh1tH2jC5Iidoil0QMtopcbbAgywK4zZ8dp2aBSW2m7B1ICPhQzxwWua
KIkv1yvbRZflRqox5SWoGRGTPyKEWLASGCrTLTID+Jkdz2MhEBUCtu4eaXpu8bX0
pOguXyNPEMZVatV3XU/9x+NWQ7MkQUo+hyx8DZLW4BPXpH1k2i0daQYIp2j3WD1B
QYm8KY2Mb3oafSXMClsXM2cGXKtXuF9+nmrKsS0D4z8pAO2EKhq+u1yGIFWduxW/
U3Qy0toSOVe1tcYJEldSeNzuEsegCmnt8LIQ7NangUsMRyFFE+3EMM8p23MMC/wT
LOwzfANOLZee376iadd1ky0Ydb3W5ZQ4ZLle/BpuAna+1bGXWE6+vc5DeopI0grl
rq6ZAhO3Xb4NcX4Kq7fJ3fk2C3f/fo3rIRi7OQ0sTBxdxAcU35C7u50ePBiVUl5d
lpcBAgruxdVYMAt+bbz8zaED40VPUXTE2rtVeygAtT14qiGUphhC/fmRm2NbNk2H
GzeLS8Xo9BvNZdKOsf8ifTHyDMnu3Nzc5kfqaBP97ZJDn/RJcektQPIms8y1G5Cd
6UmameULlBGu1xhbRqaslXwuBo2B3R9ylWQXTduq0YCAm6TxJhweuyRbSpMf9TOT
INFQcLGztesjighrb7EOHG2DiyGdZdhIm/yynUsJiNiJLRTjiJ33XIzjs7ABPqOb
lKHXlolmoJMkdDVECenojrvqA3cdNlxXDah4qz4St2maxkmVvx3exw+L5gfK8KhI
V+xETBiruC1p/MILMwerE402ABKnBFY9TybHtpG1/6sFJxg/I2uN84U3s93iHUa/
6To5EA5E6zXKCwYLCUoKWFhgXELvc6dVwpUMs+R4Fj0JVykAjORRTnGsIv3Bun78
2t/1sJeoapHEilVVKy0HdyBl4iwmU4N0hMTdEqA5+/ogf8ZfxIARBCOOTUn3wLxG
GWo4qGhJ0GatWfXwphOqdvYMFGLE+p98wyPF2Pn8c5udsOCRQnIOY3Ra2wwIIBTX
Qw1V3wfZYL2lZeGaA4JeEsf8hmIGv5/q+ha6b9bDcElzG9b3xg3ty++3ghpSwvBy
pIrlLnid+uxgLzu/yX6UrWZpSXS1OOJDg7NJdq3cfrEgMP+dTktmO1u9fptMYkSG
D04TI7dSLaDYiHAJTCF0td5bVgSIyyMq+vAti+S03ELVWMijNEyrfIcHgNH3yU80
miZrSMrlke/VvErpv8ySCVtZCPQsRIJqw7TZmTOGl+DrTVznSHCmrvCON6dY2Sfj
JvjUsx9jMPHzC/94qDOEiW58MXx8rPFXzBfnRZV8hry7DWC7BvXeHdBSL/wniLEQ
jiHyjBOumUeBVpiOnOpB+ER250HFZ2MSIX/BGW6aDkWzfALNxi6ioWM8VAQze/Xd
2mKogCWvoJR5lUlYZLvllDN2CtbhiMRUkVnE2yocC9gikhExsfkVdfRx5DlOw/pU
9qeSRHk9K1cls3eP4fRTi0Z4VNpGzqG5HxjxN7Dr7M+z7xlvj3XlgxwvmjyDTQ7u
kK3KF8NgQGBTWjL+zGXfvgOUMhgijaQs4JMXotekNgAzoSXmyNqb42K3K11EgE/T
Fvu0POKuKArFk385ze8qB6j9KXk7s42AnVtMnsrUjkOf74l042KGWUZWATJTrtXe
4pdf1H5kfH2IBORGR+QWpOOdAcQWbYr5/aIwK2wQqgqCTRbLvoiQ8QQ8frHLCmpX
CnEvAITVbPu5Qi2DNNNonRuCy4WnOPAfthMjM4lt7o/qss7NZzBtoBpWN9vsXGP8
xZ1qPmORkM4voummQIi3ICnlufDKkHXERfBWNB2iJRjPgbk+TDTMIVBj80doJu3u
AkrSRCzYyyDQJs0NmAgV8ODl0rkIesxUM47R5+J81seP2xp6/arP34zZdUai1mG0
FDX5x24BvDuzNhRHSFXvJUmitfP4WHaNRhQWY4F7hTJ4j263kdv8z7hPoSKtRLBo
03/KC5/MZ9YRebmwN1+Ml5KjVZ4LcRTpKYObKo1TFLUoxUnufQ92u2SM7JLeLMHq
4jEpE8R5udxGFDSa7Fyi975YTLl7bFbKZFbtdN5q1F0Da4XZHabUQZptdZNjo0pb
WsMVGcumXMtiJUxzfOnQzhhIgXPc2fUOsjolzhGbi5LQsjQhJWhsdXd05uHVVJtA
YTu4Cf9Y/V+/KBOYLPyun4Z3/qIXBnhPGccTzEMUOl1VrX6VWiVZ4Q5iPSwodL3C
VJAlZ8fuV1qyLIZm/KJ/MPI3Ot1VJL88iFnvpoPfvplpftG8VhvLC3prLalEmoqq
RQaddtDOkm/Tbtt100QkUvqJh+IWPOIZDOx0XQ/AO9EzRRrvcG2nyr6OCWTFVbic
iCe8RemOAohxNPuJQ7h5Q8C8jdNO+a+kWP/pTzwsHwMlNfCCaY/lY62KolIMcmxh
8ps+Ollb/hUH/0bl2BvQ0NB8wh7uBPugoT4xjOwB8HTPw5adrMTkD0hIO/E7iVZS
NnwEq/Ks3inmPcXHB+giDuNsWzBcs7F0OSl3uf6ctXYrQxjoFhPswVt+IHyoHHbW
zbWFJmIIjYkxzgEKLm8dgP7Fr8EekFOkcGZwTqmK2CvDGjspvVf76AUaD7jPXwCE
c+hKvKvAEkHG6H+aD2XRsSatxfQ+KTnhQHTh6XVfs8L0HiR9VX/FEKqeRzWgCkEL
TngZiv/vz3zX/jaDRdQ27JYxp1nQmYjPS6G903kQBH2XR66tercT0zWaVPA34gXU
6hk25Q+97Ilhck7qKlXznKCFyf4NgknF7CfcS7CTsTc=
`pragma protect end_protected
