// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:58 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
K45PNuR/vhJFIiXt7Z01uI6Z4NLHl2d0MiiNRFI+Z0uPUZ6AAfEOW2NTTkmJFT4O
zFVdhomWHAYf3/KjkbTxtzpe+mtEHVyH7T6qEh/cWLpHaRIfSlqz0rQNUy1fWWwn
vL1QnBfavZpa35LaahGmmt11iRNmRSu/ReQ33Ow5HCY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16304)
xAOMPUy7KcY9MakZM4XeTv/fh8ZEtlO/iJVzZysBB9Oc121O58poEdFSlSe1NSWd
cj6Q+8cqlh0wLL+Tttb3OYQzgiKvF+qhfzut+Q2dgiUzSZ6MCtPFKT570nVzKdIh
EUbIWs8W+lvOcrKBMxT3DwGYH40SW+4lxAKOjOf638rZh1ApH/WNIYU7zHHW5jd9
jLdMeD62I+jHYMTsC3m2epNvRp2pGxvFf/6Ubiw0LlSwue3Z1tKeqbabO33ciuoY
82fmbgPlYVAWhm3W519Bbb5h9LREoLzpkD4v48kEeLT7zO3JsV45/n45+4VdFhv9
5l2ZO3RPaBDV5OL5T6RyoIQ0YPZ98Ck5PK43V0RSGhVlo81wBBV2LJOsPUP0CFQY
2v+OLqnazVfFSLywwes4lZxyye8dsRcnJFqb22SDhrxGskKlcOJjzVEZjq4QjOwX
biWhadktufzlBmzuALSQMleURxjtsXZa8lUe0iWIxkTC2gVIA8Ef/5OwjbYEMV0e
NCQ64OTPoLQqNm9oTJUXCpylVCnvk1uRKTXfIa5qtzTMtPlzTyoGrOHN1vbKRgv1
elK6tDNjUrLbRv/ILg/IOxPjxEz9G21Pny0MGvz2I4PMUB2mr/OU+abat/jK5bvC
eAafFu3EH3bZwka1TDJ3ydMF+KzYMILhmoi91nGCTWl7VTPOQk7pxjZal76t5Y8J
UEqe/SIBNWkuqNUXaolSs5JqdCVqnUoduYE4fx+byxzcLCK5KbVC3iDwxgvE7sA0
9eKkCXT//DLue174+ReskDbuEajDywTbD/zvo/DZEMgEc4bCv5jZYMhtDgkRGb3V
YwCq+m/c76IAySK7jVe3PqwoMRW/IcmI28JSCRBlJJJRvh3ooRal5E5WRu+o4N8P
Yp0lgcNSw37Jqr8lh/piIAhhWKui7NWJlplQ149LbZVG8IZsk22yef2bLqaa5IYD
QhHl5XVIbjLjtrVTi3M6VastFgHhLsj6do6df3wZYCKgSy7jNS1EKhdsjSIXYZTv
xqXDQsNRbsltkwe9S5tJ9IZSzdWVAnyY6S97kqHOwYWLcvO5r2oBiOUX2jeTJad0
Y6hcaGaXLzvsnByZMnoMZ1OKTnr15cMjcnPN/1XVczVAx/UGdr+HlkELY+qVwC0b
/RKggFpYS+ugcTNnbSiwUKLM41/T28QEhTgVi+T0PBhxIR7SOFj8ZHoe4rTfaFyP
qLjpIGh4fFW15AMLnJCOgIZS6fuhfIwWjYnWKbUztLCkVg1TvYcTmPXkoOkQaxGS
ewR2zOV4Ghp6M8bUlWlh1Za3roT9Nhby9Xpbaj0UNh+DqIDljxJXsVItZpZgALt2
oJK+KfmgCUZS1RY7UWtl9L7PAjKiDdwkBLQffybQdOuiJURnAIz30cFf4Fdpj1tj
CaB4Fu+Rutgsg3mw2waLd1OsWqnLaQFqFXQF7FJtXnHri6cmY8f2iy+xvacqOyDT
+UF3wIPSWgZrvJGM1HHzazImf/y+mKHfKc1MGZKlJI76Uo8xF/mnV5uSZmkoL36F
epJn0j6s3jL0FXoDpTp+Q3ddnjD7r4yaR9Mv3gYLX3PCrb6Y2un0dQLhzld6UcGN
Q1m21jBAYr5bwekq9yGd60bs4xgsblZBktl+e5/FKQt2Gd4MVK/jSZRbzvoh813E
+ImFHMaXf4gXLXJu9EWGQktTnCUCirF8vhGGafDMf65LWFdsNsmMDxDhIIJBHIS6
rl356xnuNaAgrprzDGo89jZH9gTPXBveACElwMsikVQ18SgLlmtEhiShne94bKQ+
SsoLcxAAVlrkFJkWN4ODmTdqZM5F3ldrJ1cccWlCAuvfzQEHhXjn2hh9uNkVYrJU
5HMZLLcWajOpa6fna2Xa1Zm6xiatpW5K8GTx1lORhp5CWKFI+K0GqlcwChP/bASo
5DWg/Y4SRusTezqybkqXZr3UK9MHeDdo42+SO40QLh2JBjBatrlJi8uwBnhTo1ln
Wti4zjMABSu/TRITVD0kh4A4ZBDi5IwKNpn/9NlDn1BZR7hpSs1Pb6yU5xoXYVuJ
pg0cdF23kJ9E/LGup37LfjfHlsxjYMewPI0LggsUOY3C7Nin7w+pesaT7ia6s8n2
yI90hb4nE/BaG4J13pYNYdJaV2FAum6GZqKvAFRZ4OyJ/eePNtPSdhYCjJ1/Vzg5
onHRmlMgvlmjIUBxdYU7YfM8E+JJeXRVFQszsGehpOUvAYQZ07rwdSmqlX+7KSwR
+EMVYs8qwNqAYJpL4i3hOLL3BL9TUMiPOnSU+K13A4CvNnOm1vg/MyENMHE4zEHa
JDAm3mkneFjSvSIjRBcFC42Yi+2YAFKECz/uLCSsqHP3xYhyiB8cBG7Usfzn/1Wg
487Eqp3vMRTQcFGp8nCCTkJM8ADf3YRUDBIWkJ2y6ZVjho5JHDZVgQUrgpybG+Ga
NsqSlF6Z8xKmb/TmBmwEqSzpbo7e7DahsgT2UAlYhK5QG6af9JLFnWI9Uvg5j3ls
/Ysx8KjA17SZPTTekZZ6bKCAmfPwN7wn4r7TsDjqy/0F3ow/uxOhV76udE1SHfTB
sCxchOgPj38yfgEdQeK6vkOJYiwHPVkxx4xFZ/ESDGHlcFxQ6oodrRRdSG3mzlBj
OrNoNxdoXWX9q0OzIcpuSg5z1xMklxKuNkm1WxePP6SFFFfVmuEyHgmQ6e9Awv9/
dFwV5YCxwP6LNiwUP+nfnJ7FBLY1ah9NPZa89HBsJtUG/fIngxCj9YPJE7nJSp3G
7JKMZT7pMwCfPrEZykM1iY4ejlbG+aY8Yo8W8aYlppQ1m/0chhvzjx1MFaTDsbIL
S7PVuEPS4TtLGdj4s+1dUHxWURF3GJGBBORb5t3fW2qeV0zf3atlp+WUBd+ZXDkb
xBrmarO7GlsAHab1fDeO6Aa8tPsmcAs07B7fw7gukFM2fNQE/b8kFOodHKg7Ndmh
SORIvpncecDXej86wibEzpg7g7Nmr0gPErjCZorkJcrTGsMuSsYnQkZ/DW5A9YxG
Qn/ShmBH2OU4s5ZOI5btrwJZbjLPl/lttrmhwI+9Swl//ulvX5uyOnZz//ghTC4X
AIrte57U1dL/e7W2j0D8CYP/JDOz/n89XJYZ6rzaINUZUkbXlYFF2KGGDoJADHO1
1FvXn0+eTbw0FfkrUEDIyCYrgpaurAXawd4dg6iCGkgCl8YnD9aTffqfzkM2xR/I
jtM04vEJ4BbwGwBLcTk/dVh73Kzuy/bSX3FCFdkCqxPO9bsNtTvf3oVZoq1IH3sW
Yllh/H5GkUi+u2w1ThYRtm7+tYMaYHp/bUMx8tv5pZKLPiL6sGhDIEQbuGVnb82n
wIZN4YtgqVnHJBYjzDs3tzF+kPxMoreQCco2zOGWDbFgNOZztB8gj3lTuiN95Wi0
aPghrpj88hZezq8HSeopEO1+bR7lUEMiyT0EDSEQZrrwWGKiXMfrZLOwxLDBVnUY
jY2bDbjNQSUfT5IdARV9XsO+a1cgTvwkYWP5ni9JRczustQ0UHT3Cf720eWVpohH
BuzPfg/fuqZRer6wwS4iguQe1YdQW28gSxxcJIhM0zwpMJmT407Cb82rLSzJ1PSF
vWwqzL6bQYqK3oM+X1mw5rttF42qpQ/x6S9oun4LO8uOexZMNzXUUN5VbCuY4cp+
3DFQhRKdTAlEXG+Kte+eSRmvWiw7/Bkv2TG2Y7pS8iEdFhHTz/5YWHiI1xmJ/t2g
UlQPnZmGh+AuLvk1cG9Urcrjw6MCWEwZG2uK1Sjq+VyI+ixc/z1TLR0QMM5UE+kp
gs0uzw8xDiAKQR/xVkT8nA1xcaAaGzL/2Xy1A1GkFpQlF+wwEqBJpoM9DLr8LM3g
KdVbG+IrCxj9gWr4rjwsLa8EXA404p0clnzVic//kyDeGQT8JcV3QKLJpNQ6LPlg
offuTdH65Dkj8vK4U4txJ+sgA7dWWYvaAZxRM0kZDcNHtnMllj7SrqIQ6N3BmCgf
rnqwrGqw6xfuwQdeMgAPLJ+f/nt5pEu6DyAGlEmcwCB/MnXl/xAeIBaTjduQeKjz
fOfFXRyt04NqAHFTEmw88KGKVYPJvKZfeb/U4O2ikJGyucvbXSaq5fLGbDrVSnry
Ct0sCn5J5OlNEvbqeRPSk6l3PgKzSb4m+qzJ81sPOrDCk4DFcRarzMwNiNsiq57h
CSTYcERjZY+1JkaJqXJDEc4OaAUFrR8Dv5omU0aksi13pBEC4fN9Jg04a2lCFNCa
n83/Z/sZqLPOqcPHdoktwxMe3vtjYu7notj0XGhSjHeegpnpjkuhoC7BPkOkX3eQ
CLj2f9/GQZcYnB9b1XrTDUhvD1eTvfAnVOuy8rxjp9MjgIpShvyw1KQcEPk7j/1f
DS9gC7HrOAeTsH85sZhkGNEYv/n8kMwoEkTELM0abdC4o/eIPvAKad/SRMdITgg4
UOI7ScphIE4Bjvm6FTRkZS9RtfC5Qu//PjZOZ30UQxePnqOgBM78LYCfPuGDiTXo
YjZOyLofHDIizqbR9ohqo8PCieX7wedItgAqWeplGpXx1h7fZUExrCPjanMKXdll
bv+OkF/S+tj5owAN95A7GUeVIRLIgEfNzQEZQqYpxCAbVYbDNDIYX5/upKRX9uQu
6/N7uvVe1Wh7JATqEhG+rL7t/bBBOBRxeTv3boNidiyuWGksEwr43AiPIAJbm81P
kIzBy8OeUiMCVCnWEVWMG8ZfZkeWbdYuW95SZjCwV+IH94Bcxr7+VM8UnxJNLeJZ
Z/j/ajS3NJUx0IqQgwgCUVnbOGL4k0QoOLa+zFs7yLafQhCr4MPvJPO2jGWBtSkb
mRbXRq4HBtEzMAHR/QyBGY1HdN6j1Ny6Eg+sBHuEGE1WY0GF3yQwgBoIcMQQDXfN
OawuRxXcTkiR1aON7XQ1xoSnjBP8KUz2QGUlRssQD9/CwBKR5LyeXYttZa0Da1KL
+c+LWp5qupNGgQkSwxx0ydrH8X+7zTan/Ijs/ga8am3eE/AABunRs9doRyOkYHpG
VcCSJpKoULH//ucV0t/fLARDR8YfWsQ6w1JFO4ozbc8f21UHSLqmB0M372m1C8KJ
0XLMcPttq4bYm/dbFpkBuKTFOYuviTWFpJZmwNqPtACu7BFmUqecBhuyE8x83U/q
KjZkLS4Gm6ejPad1RMI0lCqs5Xo+uTeNtsrltZYmw4MQGtGCQ4A3Y+KUi2Gl5o1A
IXbBHJLcMmraUCWOojNhF7ypgDDl9J4cwprTUe5i1lkGlGquKuqZmvfr3Cd3ZNUz
ojj+YqcmP91WsLWLJhpK/hcz2a+2rWgvlHm7yOdZg4mFEFQozEYvnDmqw1im2NlC
Ti/ZYJYatG+41bQZiZG3yj0O+j59wxE97LnE0Pw7Qx2ZkK/Qm6mLikf2DorF5bu0
TWecxBXbx7aDiH61DZ1fjxFjmheVGFsfQiXC+K+zraxOgEZTA3zRmRD36DfkhJnf
7MYMQudJmZoNNfEF/YbFQB/mDy4BMebrAjUI3pDBPiR7WC3lNkylIAuaMjWZne7M
2cb9Lh8bRYd9KhhEAiY3NaMbfqfjplZtLw0rfirI8jIV6tGSeutMggu6vFqQ0ALD
u9Ob1eClpqmC7Vh5mCxBibbNAt4V5QUWb32CYFtSFrpRoYSeAxyaKwOLuGChhZnS
Xrpxsno3nws9gbOaYDnYaiSAHi4xWjLQtBGD+SbsylE5ur+tCJx4r/jeTZJ/+mnL
Wde6JY1mz5/XdxN4w0bY4t2SVUcZrpapa9kMaYAgCKbLr/zD3ITDWckE5e75sNw1
TF5KeKpNZ1oOeYyaoaCv5TlY7HkqkXxWrF1Q3YOjGlmdamB4K9CMtSDPcRvG3gKE
ioiN5UrBn5jdpUkjrbLOWTyYDRB8S+DaleIJovVZiZAFr5mQZIv0aKeQCKzkWVzu
U4rtz2ytwK7L687MKM9AXHjUo7Fv+DOronBf91Zm8yhR6JfvkdA/f/uhA87VfbxV
9allsuKNxdonnESCFrI6XTaHBCqOAPEgySkMeKnVg0rqW9jyheHLcPzrUPzlRQXL
GaD3g2m5MWw97dTs2XbGgm6yxMCWGUgjeonPSF55SgPPg3RcMPaiZ7qnmxPQrZ38
eHaR8hGGpmMKz2tZepHISfRwCX7BpoTJRZ0l1RZgejtI9wdkJCfxjsVk/XTCGZad
LYuJtBzgwF1MqJAvHf9Ryc0i2ieWIufKP38ljoUH+EUUEPcQrSS0W+bTeQnUOLHg
u2xJS/KqCg5ZOh5tufJF2oo255HzQbwl1+aPbeDzTfUJPDD4/jzm7JtWWHQVxqPd
doFyKxaii3TIPH9b4gN5SHgOqPm0sw/8Y+iE49/0C8vYzjcac1rUz3dGP7606Hrx
bsVwqkouFtQ7EP2Yb2TWnEW5udkl9CMNdCPP1kArMiuLYR7d7kP4KzPLo0njEavL
NOaFPVSLoQemMi9PVZTsVA0UdY0AbNYPbtTCfVU9X2X5qz2TMSMmdY+eHTmnf3ya
9k/nrrwy3F3h3gBKpJbG0hVsoPuIJr1TLiMtfPkoCnGCUvs8kvLTeKUQ8aUmAg0U
I73Ra6PP7TGYib9R4BEbinvQCG/O8ay/ddAlsiGh+1AEqj0v87ITG6HRUFbKQQCm
KBYHVVqL84HIL0m3i89GZCeLb0c1lPykSfKx2UjQuetyKW3bhpDjW2QmEV0mIi5U
7lHfqAek2B9FQIk7BEfvJ23lRftMlknywqzct5UpqqEXms7zbeoQvd+kkkEVvdwm
57BG82LGE5ZFd1TOrtX8W08RPBsPxR/TFCuzlyPpCD7kXnZo8UBU4iJcTNVr+um3
7Sved650r80MIVov1QVZyvH4dlEGdwB2T8ETq+MjJ7Avev1OMTpFuYBQcFAbzhb/
rscm2nM2LHgpukLD/q2YWeunLo7mAJY+fipTtYIkwKzIomw6JOGEseNpT5k75ARd
RdtVpOAuP3qTT6US5sN3P16VY/p12ycLNh76u1kDzsTYFyX3rCXp7dPOphqM0xoC
6fYnCCfyN+gN+E8WMOIgjO8wzOQ/1uj5AmEwxGD45RB+0XaS/0UjUppSXpR5CCyp
/KKX00ysys20SPs3LX20GqdYF7i+sjh90l1mfvHrNnEKw1jLi6jXesqT63n7lq1E
5ZUMg93Qm3NG0lQpXj3kGPQ2OJoSnMZDGcxeHlEYL97I76l7uOWvxxaD2TeQsK/K
8ApcYDp+8CjY+9x7zKAfNcYAslADjNkuzgoub/A6Olw1Ry8WioJJJf817paUULJS
/I+MPskZO1XMDHlcPjAx+TEejTkpNvung7pXQO8PSCYPAcPpnGjCaHqlsSL+oJJl
KERelzovxhlu6P/Hr82PyIKg8Z71F1dOliTgtlJoLoAk1jyCjl6H573z/skCAYqA
ypExA9dKO0ZsHnIkqAJ1CtHj30RmeHqK3wh/07ORY50jhBtRERqUNPxRfN4b3v18
7jCH5Gfney1RkcWb14H0nICRKNowDTd59tzmwNfkdyMJvGhmJGy0jVvFcMIq20FZ
UsR2Sx0HF+gi7ptM+wGRNrPKTKx5dV3SOlp99edOnh8qGbufhWGIBsh7JafLhgG1
J6fI5CmdfIOoJA3afME526D6FUBxjipuRnwn2+DgION7RKBwGlqmWiwvz1/RPsbN
cHoeB1DA753e++iY3G8p4jNRzgg4fYgbHagdlpHcdT7kXLddTCOzzkwnvYsmHVxT
9ojSzurSHav7Ro0BP0A2nauF6OrY2BPdF0Pr5St7bZiYN3Jono///SYc8KOgqC//
eKspC/qypP40l7H1Z1CJiDAMRxERRtTbIKFx8sv7e7dvFA3zj2PiojKAs7Z/Palw
Yvgm2E4YYRIL+vjaNcV4toyaRrixgL3LBetGIEQO4So5w2ijzjhozsJW4IQJONQT
rN/V8UR12erD8KzCRGN0leA1k+9wYDyY+1UWibt6G4bT0bMvFDh20s+VTcNf/vnV
DDbl2GFgVWdDfUuiUWZONYsrQjMrVOfnAIlLiaYuwrwFKaEPtWHNzMjaaJZBvbDy
+4zXyz8mgenyk5FY326nvZOhhmmprlmKmNIbuQi4AaVlwZHK/tV7a6p0jQkjt8DZ
YEJuJEYwUGkI+rEYPymkmvWG15FpsLISizrldu8upwDxrVhMTJbJiFYXk3+rh2lu
IOKMpyzDp1Y1HbsyaYQrp5Ci0p6IsH6Dmib4kAu22VjPmjb14kVOiDjj6RmM8W5u
nJwPyqrLfUGLMvukZAF/CPAJk3bpKnPE0VlpkO6WVta1uQdkf08mVGikVx3k9UOB
dqYswRpJIlLilFXX7sA5rFPW5jHPYXb9jlpe2nnaq0ENHuO6OCwYCdLYdNqT9H7x
hWBYiOACudYkEmBl4eJvLM0oRW6FfbhMsnl+ztk5YnzGzcdsvln8iGPr//69OBoj
/h3wuLVUlo+Au8ouDBvB09GLKxPyTcN0Mkfc3SgjwhncpB1YRlJbV5djYdXKzu+/
/aX6EljLX3YzzD7ZDejqQ65HoPP/FRhasXPI/P/HqBPz7G3gziXLneErsd9s6x6Y
JmSn68cpoFJbmzeyVWWlGhTdxIBxTYrooJXxQCXW5l8v0CUC6TGtuZs+zCnD07NW
RvZYU+xyByRmMNy3tdx1tORKyNsWmr1VemB2hVnqYlhDuii27PEAP/p0JTLaRSuC
ZpoR4DJGxv0t3OHAQ6Bdt4FgaLe137EZeNy6mgOQYL4Z/0ZvyJN3newo7wUQy2HY
sjh1QICH61OtZa12HmKNSSOGxiVU26A4qTz1ZMoGzMwFOygElpeNzMIj2082Bdza
7dCq2ZRG1TmAh9feD4mdvPhsODYImzju81J/uxbZGFnJOnBUCIWonT4ZyZMtDHaf
FU/VHS27fWOJ3XpytpNDhUMmvV7vcwiuBm2jf/w0Xdj27rT+/opdEytGTpBczIq6
rW+VaGEqA04XGK20m/IsLG7RWaLr9rU5XiT06hfCwTgt0But8h22v9k1LGChbe+K
DI6+iwIXxDhnuPCe+f5Q3kUA+DquOlIxFcCzjRE4bUgFExzlUMYCWM7xNLoymcuc
4yogIRnHODtuMGjllbc/9d8nsYEOvoC4I/YhL88YzOJf+SdcrdQTLmeeE9+JbkDN
lqbfxU/sJjtSvBEEcg9bnCjgFN8minG2gFD9YvTOcUyJ1MM8smQ6HjstHaZeyq4N
uEKDl7+rULhQq0F9Z/uAVRRQuZhaYuj5LHBma8pAd+OgJHUYWhniO/m7MLk/PSLY
zgD3uj3huoP/2uSGEzul5itBZdcp2byVA0rW4BetJUc8ZqPCpuzpiJrlG1fbid90
c3ZVw8kvez7Fenwu6uB99d6fN2UXSjVyuiGEEHENVaVaPz7mK3HfnglSscNmXx2w
EckPN+Qc0SeYcEhyvLxfKNYbJE+KZurN3mkF2vF9+1n9qlueNZtA0IaTt5StRQgH
RRBjhM2qa7rgemIQH7PyWGSjint5mYEgMraCIlAKLIQzhHvodgo7Vkhc2jWP2X3i
eg618++p82maJ9O77xN+eNqi7x1sN3uM5Eo3CRaHetxZfaSjQz9mKLxAAfhBEgCK
xWFpMcCVlsHVo3dJFcRn18k/KIFluw5kU5iIIsqfRe5UF9+ranwFTBEtjOEou9dK
XJyuA5Usca8kZ0Po7SiayFpdPIAIclab0njezRMPDNFHXWmzCCq5rX8LPlyX2SzP
XrEY8WRYHw3vK6AxzFgkBQVmwHUHtYdmM0I0vAP00pS8OGJKG6K9lO19eQROvoQv
lFUG5cY2OSUtOSvLWlygoynT4fykt4/AScpBMrubBky0zBGsKDooeZg6zQrjyhkq
Sj6wV3Xbrjs1r1Gr1o6vrcWmHd4FuhU26Mz6aVTet3wiOwXI+TcoJUMwL9q+T7WR
MEiaHDePujWJncRWpnDElE99zUievclEfxrIwuOfQuZYvGv38IykWyPVgbQyPE7T
ZmSZ7h95C4+BbXAg23u4Vk7oTGs5fU/dDHsu7SNR8BaMk9FD3qEBg4K2Avv0Rp6/
bY4zzlED2195EvYhBe0uWrjEbUA+z3jpWw5DQIDARrrckKvih8zKwXfeVXE3jcPW
fOl6OiLm6ekCjF8s5XnBVWRz1jxPfGCqA++3glXn5YmceEC60vOByN14kBYATHLh
oJTdIVJH3TLzwCLJcFu9xt3/0O+VtrXayWh23L6xZ7HUpdd7V8ZpGt8LlAgai9lK
DHh9OdMGZOZT2ORbyYwxwsGaxYDnQpontVj1P8/eG9Gsziau8Paem9c+r01BquH1
wz+lhXlpUoervGGUKa6Y8fOoNFR1Pb5FGw1H6zoIoQzTJ1KTcupey79Ts5VK9L9r
FKzw7SaivXq+pNLEIzjfnIxr+0RCQwWO2TwPkW8eyFzLFfD3HOvwNYyuvO82HJlF
qX19BX1AnQkxOkX7+lcSNSh0Ij4vdt78zjnkYEQZWvXiRZyNXTPKRmV8pljrh7Fb
H4cqdgwGlM1b7hNi065SFQNNDrYSSLos8q4WP5fRVwWwrZW1mfzu2B0RlxddY0n2
6CWvBoYiPDk/1FSeRBg0w0EKENezhhgCVmhItkGwixfPqK8GnKGbQaou1k5uPc8t
2P2dmFH/gg/5mBtLmlDZWAQRod2ZyKuJZFL1C3RlApmgBt+h7w15z2XvYrc0TE5T
t8l0KnST+POexoz0oqKKHc1OYcaZR6l1fhWMFhKzz2crQJ/pz14h9bo5AHFn4zSE
M+8Cw0Q5O1cvh56E23GWp2KC/tMUyxz386rFs2/OnOdZhMu/rS2jkso4ZxmYyF/m
CwWDzmM9OnRjili3No0qrQFOYOcAo4J202LH91h3b5Syd11GkIrqt31eaokFbFBz
QezjUy9sif0WstlBkbiqtN2WFEw3BrZSmSCzqMj+WQKmUjZbMp5FH+S2GiVZZUFr
09Jp0qvvqgPHvQZMYB6suhyBe+lj0DnORZn0DuapbuBkNuz7nS3SEijA+RxB7YsV
s+Cndwf2aqSbUPvSaennGnhIcrEN1DzAzSHlff5XTTlnZ+CCDFXfLR4FpyXQFEWS
G28l1TBsLmIPnsaP+vUmNoznZsDAW/o5X1vKcE56lXc2BRfIUwH28lI/ERt8bxV1
6M3Sbvh++9WKMeQ4G8WNA+rV29LhI0BX9MysW8CN29kXr/a44xQyAJlFXNklYS81
X0g9wezAfYNMFC/7M6LsDsQdwHW19LUmXNCeFNzvAbHrhYkCBoAjiLL/K/wkB4em
i99hMONPxorfE+EjlUL2uHcH+Ngik8BFFHJAeUlEaYGAgXh1ZrkVuwx90jtNmYPO
7kWaPH2sMkq+gioj2mTM/pBvPIhT3/ZwHzPBwOUWhO54z8XD0Is+hRPDWsJlluk7
XVzAk5X+wWfXABIRvoSHSNWqyYv99JRMmTAsDnedkXj2kMopKehFaECEONvI21FW
omBqgXaGnfR+JeNT1SjLVltdakDD2Ss03/g8/5Gs1rwmp7JdZoaxoO96hVCsZQNx
3fqRb3iTmejP6W8KLu6wn8Xt0Xny+IBcajvcvmo5zgmwuGagyQSbntsQ52JghsT2
qGN9LUgsKUS6wplzsZaLC4egPCIcL32nj8NR9nc7IaXuS4A6keoMGIXwhyl81WiE
4n2VNYmvD9ER4TftaYCWyAv9zDdzB39vx5gjecnb+WxFdMDz0xdv5HVDpNjyhNrk
XJZ3N5s+iv4NJXCdwX73drXDnAagi7LFZ1xSSMFCW/1H/L54ojT8aPv5QhlODz6Z
zMlbw035WgtNH+IQ0HONshgTfLu/3s3XxK6CgbuIPhyRI1xdUX38VKTDlaJQUrwv
KzYBSsX1sEuphN7LrPk/0MrV8pEf0ow5T3DHIl8SF9yXhuAW97Behmj0mYLsxJtd
0atwJqfFajkB/1bKjAEwPfjmnjDXM2bGf0DlTHXWp3ut6HhmzF3LVGPVqXC8gjV4
n3UdWPN/63VNd2joOXPn9vdigo5U6W+R2RRNDIymTIJVqthZESqcp8WPdDWK7rWe
Xw37IF0YguGLb1Jm1kX6JZqA5aIr1DeMvjJme2XgG4Sm6kdygaSkHLm1hPd9NuA9
uR+iBlq2uTkmzwcGfIpoz8hzO7ORsfpMS/9G/LOyHgWsFTn8aexTLD4m1l5mKpsn
6z1cxkU04EAZ0l3aUqahVtzOBmyVQ/O0hlbZDld0mxnJwTqddytHAaYvC7n99eYq
kuI9OFM0QtjeraXLAzNrRk6pv9hLz4lY5AneIG6FSOLyLc+BwQvHWUQIw4R7EkkF
Dsro9iE56vT0OB3z+0yjGFegwfS2t6u64WUYWvvQThpCyZSnK8RJXd5H9XMLn/uV
NISfSbB4D+rM1UyyxpwOZX/4BOo7KkkoAIxd4HiFXB0f7IKuOibDDUagGEXu+7HY
L06VeURIiS3T2O03cjE+g1JIoin9fxPsRkF9at5+QE51aONR2+KcRwDXNFWOmumT
NnVt9YU/0pmsWG2N1pkLwx4GOi8lX2dQ4qFB/K/VJVqaOd7R1CHdjDrmyHfEgSLL
idcCaSB8aQmlhxSXdgngCT7YLt95e9gK7IGyeHMMwLz+4NS/oQP3a/w2oH3tjQjg
ttj/cdDXbl26e6i2nxDiwj7AHq1DidXHMpUsPopOnKnWccSTZtR8V5DNK84uXqsx
dJtloOL4OOfRXlWLAYe8TS9UqWx6VFgPeUkMKPJdJeJNxbSKxfHIGKoULMBYAt8+
2dCJr8nMUeMFx3j7OyLIHJHrW2OjpH8Seh5IPJfRHX+OIRrehUm1qokEaIPMsc7k
Z7ZU1MwPfJn6KANkmxJSKPzZBV6p4qPfzl/iSpkvGgN+qdnEfA5GiGQNf3a3CUvo
V05MwfGmV7eSdpQD902bOQyltrOP/O7ozO2dLPRNoc86oHpw/UuTnFlsRsa7GmiH
c+tS/ChafraNslGrAAA1xxnRsuzsEa0U4p4FBTeVOzQLWBEKrDvYvIHNvzmNY9s5
gF1bt+jNwQyp8I5AYNJVSgFpIfgSmLKgllRZxgod62XJgP6qjPJFq93EduJR4xyz
l9ex7b2izhDiGcXnNOdHnonru36t0ff5l8B9sU1b0fAV59WgPhonx8nzXCO5GCoD
zhpOoBmJoSYmCKqDVPYwsEM2Airhl4la/eBaOMObn6u8mei2NihOHlubArEMjV56
+DwXjGdpDsTeJqqc3kDwOYvk+WKCOd3QSEBTpMruEg63uUsrHcjvb6jNOhlvk0ln
oq0bCz107hl3nBCKlfkskSNIbqIv3iBKqojOiK0nxTG42TckF88Rhn8nE2So1bK7
Qts4gNyFyiy74qoe2rM8sKdyxJZpHwktDB3GLP7OOYP9wzKCy84BrUIL0DLfr65D
vPwRopi+8fIy1jSsIIA6tOZI+JpFxRcslpKnHppzAzw1os+EHmKNVmxqHlL+b1I1
oXflcqGGhSe0WAZvaA5ndcTO9gi34igIAWe4/UsRIhyFyP0WDnHOuIKG/nOAhMyS
LiCZa7k2sabaZwaVlcr4rHEVceZxE7cbD0ciGINydRap9tbCT85wouv3d8rAnrRe
c7evwMTL2mQRtp+e4xRHAIx2YsluVjIex+l2JvthoMMSbyBtJvQKpHzKGH/3prEL
0UDIJ/WfQQDdYBYTTWOMY88hSv63G+KD85zkwMvFegL5nHhLD2cwX3PBe9cBdcZe
n9iIQS5BgAsU9L0qMu4Q41+YJgmDxwQzU/EYZhaKoFH8rwr+uyUFu+Ka+t+2wuTa
WHKtvRAvp3Vj/LnJ1r3N+ztykONC80HcHp3QjdbXTzfrwsr5hDhpulz07U/DyYmG
a3AnX902PVzEroZOBf7CnmEnzh2DPZ12tfcpdL2KUCXO+i4q3HnrirsVaV9IDnxd
f5LQFvNUwfmLdROzv9NDCbRIyNZzivSUhNLfww+DhyZvnyCUoZphv/HaNKgSAkVv
7b3dT9jgMKjyFMllKnpDAY5vAGU85KICFpIjFfJRLDzrfxIOXdm2zHrkqbUwgaO4
3a1VPiQDw0Dx/en80MACyckgaYH3iSlgSQg0a252hUR/Zf4pH17JTvcOp1Rs9uX4
9dVu1GxOEPRqkn8pru9S8qHAEiv41zsR84Ur0kzBprA7q5DH9YUGtNNymyfSjxpi
HXqSFtUQHX3Wyhi3c+5azVznrqopP6XLtcyf0OWXUqP+92Z4YAGVOw/QZyvBiMU3
q/8gk4Nyb4fUML/kf2nZhl2Hbzgn27667AGhTYliCVccfO/tCv/HCcSDEPJsITjW
qdTZJ0iLzlQhMBuDRB25xUHfKVxkImafhYJAJ+oLBKkFjQ3a9D4Wycn8EjTLUSLk
0tAcNOGn4d09nNZ0LX1xt5rpATjG1QXlz7YMYGIBy9wUM5jv+h4Da7HcJmYFaRUc
MWqWIn25msS3Muk+/zhceZUKb9wz6RlHi3xZIAYLFCBKsjR5D9Nd7Z+rOpep5Eno
o5LKbexaq+DER3CPmTeA3EoNXLBRQiaicIj+cKyId8dBMPI1Mk9MmSdb4fHhDdHL
olbZvOZKp48GK4OpBbpObjg4eGCZorDuCSHjPby2H+rHBNUtEPKkXwvosvY7q5nq
9gcDBIW5evqZC1QAtNP8cvU3870KEEWu0jpJejU0FGsX2Rt6p3kQ7wX1r1CW5S2U
bEeiLorlOnuE6dke4Cj3RvAu6I/Jr/xTtQgb1erDXZ86RpcMRER9uVYVp2a1Ylqh
cg2245gLmj6qKynH/+chWkEE38u5Ix6LHdQK0nrgVnsZilETwKr09C+QruHKakPj
XsAVAkIXAtNC0TZ4Xjc10L4t5+rY8EUR6u6iVAFmXWmyBdfbxxubF5HfE298TncJ
KAUDtKgQB4TMxhpsyGUBHW4tS/0oZ3GpdLVR7+dNlcfuwtkpVwZQQW+XomUsVPoo
bKUdi6retS5yF4XOPfZqgvCF0lliHK4nGH7JOgZ1z7lGHbh8OjT2ezYOocgtESSg
hRzLJHDXcR5ddjgIqGdqRAgYYcRcfJTbHLqCYAThLllmXXOf0zBirLzPmaPSBELe
g2uJxSIN8mpgMJ6PEUFYCm9yX4gFDdVvt9Rt56DOsloCj5UwnQj6Md5ENygzW50s
IaRcjLzNhMzKcFnxylv1NtcvSiJZ7D+01sJOR1I/0kjXX8ZMvLHbGuXTETx7qeyi
GmtkYHpe+di++EKj19IT2LaeLSzDD9oaRJqdbQXGN2T5bJ8lvFVm8V29OVifn8aJ
0GhfLDLJNheDv+wu3HL1nseSV6bvcwlYlFUYH7a+f3MrPHo1d3UXNvVOghiMM+RQ
6qRbCqKepySt3BPqiCJv8WAIO+kCV+lEFM9RsdPCQ8jDcOchMnbrWxRBoylrNvFC
KGv88gKr3xstJQ+ujMKuLIUZJFRWk+7BeST9vSSaNk2HErdOqh79CdYHVZb5p87I
tNV0GTTTgPayb0Mv07YYIVcS86FjRgAJPLXwIU5SLftNmRInXY8NgbMhYReH6Tre
qG4c0M8m3lWd4XllgMUpLRpB5S2TJAWdqR1aBsQf/+BinW8NS6yoRgsSfkgsbwyw
7vCWwFwIIuobPGA8eRDw1FEFyGJI+sId2QUeVsbCxRlyf8QqbumSkl50g7f+Mre7
prLx8nCfppTAhpo/U1r3ID5ZRTQTxmDrv2jEzMY2sECL+bngZ1T0GhCyTX10uL8H
x93KMye+1jqZXVi68DuuFdpY7TzRBbEKx8DwA9sl72asyM7/BDuDKD956H0baBd+
+M5Fg/sSy8BooT5K++4rQFicBldjnrIrsuz1ehNOwz5MV6K+GQf2YQpl8rhQW8Fv
ivelIZf3WEJlsLOKDAsZF58Rz8gRXVZDAeoGIdDIXiKDe5Ki80lWXsryFEQpDnv3
pflds7hqkBCo77MM8Jb1171pV4aWHiB1XxP8aJNAECjwE71j/7HbGL3ndOTlEa8S
6LaCMflAASA7C462cSQzhDo5HJiDX5QN8NMnjyh+JxcNV0WXtZV4hUaDzYqBV7Ub
OJZmMGJpr7+XIqT+ESSlkPJkkqbythjrxeQQhtD5mV8rtaTypW/LCLzsq7ftanfJ
JvCy0yOrkt/wl9seROeqaUsRxTlZ5nigPFZAg4lGBEpuNiyG3/cBmLZFcv6vTauS
THUjWf26XKRNGG1JRqWHN5J8gbiWOYRIyBWLf89YU8gR9HtOLrWasFz5qSWlmQCa
mgRZTEO+IkO9OGZCfgqBK+x0BOEQCEvI3mFB7AFwBCNE4kOIrKZ+1v70m+rj9g/x
v0sUtK0PyAJhqbeaCpQGRrL3S8yzjKn+GjZCy2NuV38lpR7SatZ7yzogqoiMmDl0
qxBsrdej/pMaiKjy3nwnuLfIpg2sMJrJG3CFjCLEWZHbGgpVaCCzQsBRo/6e7M90
0O885uvzXbo15q4USuh9AzBXZzkE3JABuYTOJ8YoDAUWKccuhjM1cgSyj0fmXAzv
1Lia0NTSm/p/f9Pd+TUBu/hvQrrz1OvL+YssrU4i+RdTfEZbEOhft8b3WbvEFHVX
Zq9EwKA4+0i+8AS1eD1NeZQif9iWbIqRQ+3zLDlN/baM+CCSHGFyibz8TZ5AFpUV
sFhi8CtE2eUz10uTwwuRlWx4JVc49ePtuxWSM/uuYRft+0uAkV7x/SwUHkFy6xwh
qmxE3LOBZmosZdNbk1tMOXd5VANe9BcH2f41joSNyXxKJqQrYWQUi4+L2TemW08t
OrS2J/coPPQAQe5JSMyUFg3JqPXcxjqKQp8tK18BxnVXkOXTRa39WMJPHuAhlrR9
KSEGHjfJJi4HZidP0df1NTLTvopVebYbEteQ7Kk0YCumhOIidch3h5LWnUQEN2d9
BWARYiXjUp4eNMmupKKpDwQkIy4+v1V0z8HVLDdrISMcj0H3Hej1Gj/6XvNyjOHi
ENDZnn4P3dMnL/UonGfurNCjNjrYxM1q6QFZxJUfQd0y+U5spGdE4579fsu1FiTn
rlldH/2/grxD9pWimKYNpp/LXewePsuSCtVVTX7Wu/kO6rjwHyZqbo3gQskDGFxT
ZAegra4dRw3BUGP0fSAlay6bTeQwxZuweQLxTMKKn+9SINdyguFKxoGktu0MAKgN
xwyBzZgEX805+PqnBxG4LD9dIlGTEUlheo/aJ3y2Cxg6m92HInK10D6gMBrAGI+p
UoamFI77VwHPoCcFipkjNeheTur5mCFrSL/LK17ZRzvz6Zg3xdmqCq95c3iqQg/n
b9p4GC2E+/EixPXETgPdUWAFwIv+xayx0GIim2xW7RmD4YGpqKDaErb6D5ooRr4+
CWd8O/adamfHW/l6KLGvRic5AtRuHuwM8xPyUhMgyw4VLHYxsCW6LB5ytSF0IWqI
4Q3mui21LfIt6XfmEZTDIEezAX0sFKyBSPFj3xCoFCdwYxE2G8LmpnNQHMfot63o
eI2Aquh++UKfB/qNoECVlA2jjoNvVD3S3dE4Tbyn5t4bHTLBdphBffswD38M4Nyb
ET+2bdY++h3nNN31HYBnsnPTapcHKs27bK2vso3POUQegyQkzYZOubdYWPffJwYs
wA99h3x/kAzKboCMRFKg9KAvcyTVZYWgAbqPLYfTGYXt78cxNUL57mgvQG68nPMF
4jbC+es6yLZHsdO0+fGYkfihoiA3DkXGhMwaXAPot5md/uOKKmss6Am4eeiE2Wj6
UVelU5vsIhgsfMD5clBzyZ+XHmZIIwBmiViStZulCyVO7WzxKW5fH/jQdJnrJJoy
YSBI3h6KPeOKVZsA8PKyoaChy0klIGQfAmp1Vtqu5DN3MZ9RAk0jO+Bl0Lizg/pG
emb4ktzpXnB2E33wOnVqaAoup9ITn/9rHgjgnbldDmLfSwIwKqxEivQLumcsuWE6
bj8bAmgYNZ/YxDoJBIk4O5EQ9x4JmgytXkdLeMUbN6h0mSQJsO256DPCdJsp1yE/
UHCSA5axFX8hLvPCOWGUslpwU7pjES1RfMOMNMPq0CR3eZbg6FpHGdGXHUgdLc0I
Os6GXb8hZHz8KLuSQ3FsivVIKAcriojTdf0Wxl6xCxlkItcqHi/eNwvF+Tsmzhcj
hpa9Qiiq6jVo6XYCGqkJeFjlBio60+ZhcaMSOrPn255yftKsSNTjAO4i1tikAC5a
ApZaDpAqcd0SA+XlPFz5anuBSrseH1cmCGp7tbXrt36ccYazSsW9ZkxjlPkx3KCE
V4W0WQc0J7y1YyFCqN5yYSBf3j0wbfmF3HxPS/swucoYg47ieK+JfvNZcouWXw74
Rm6GztEdMEj1bHPRYRayHavSLgRdDETWoZtIH4Sb3xJrmcjrgjZL2VaxaPDM8sjI
tu/sm1gSsIDmTglF8uNJBWe/gAPMEU8lNzIbSeyuhkJRYjAvHB1mfY7VIrYDmSD8
O3/wbMdnJRaOBUy28kdrWR/IB2pNVFleBB626qBeB8Hv1xWtKHRItJwucbp2eYWA
p0M3MIIG0uE/evPF/exBL7bQghUjP9AbCWlfWv6y3HBYwV6RLgwnSDbs8ZzjuxPe
qTz0bczOsSt5BQ0ijOC2ESMaG2RKToEtm9dXqN0SlTiZn0ApJA+TgovrLvTGqiqq
QQ85HvMH5jQhIH2Efc3EH5NFQgR1ir1srCehI8rGRCL2C+MPH+LSEacJd0nKAGmn
y9PiHjyfis42dx0j7YnhP1D1kQLVH5TnHw70ykPQBMMGzJft1Y7VZbKqsU4YvPU1
wiJ46Z/H7rZ89+tAuuZKPtApX9MfJG+8oBBlR1OdnQAvh/3s93dPO7OZsIPUcxI7
EhFWzdO7Qt7ghlfhyPTSTMKdrvEhtSaGCLYadNocTZaC4+2Iu2lOskrjb5eLWugH
BD5krgI7eZNM+/TiYnOnFQe/zSiqmg12nJQUutTvfLbnnOnO8sMERLwnz1Oo/hMs
F18UNfsqvidiVVmaCiuNCvWif6iRhDOmLH2O3uHm9MktS9cczxmwGiRhZeCLqgfO
nGnAYpqaPpWs+KiYznIym2g+JHoOhrddWsBRPudjFX0wHmnaDUPWX/sGoX9cWeoz
Ug4os7XkY1/zRuRnOWCC81Lrw4XdWEI5EI9x2oU/9BqszwUDR79O60hCUk3IGnhy
oztQb3PqdFAYQh8U56zjdyv/ddFtZyvEUiEDYMoTicP5kr/BomGd7WTaSAzCrLgg
FLH1WXTwzKfu6X6O6+pHlQSXScYS7HuGtBwpkq9y8jJaCQwV3zF5AD4Q6GJ804/f
Tr/MB90u9lt1+EsIkDeIzedqluCFsr0gUO64AVpB7VuImm4osnKWCojjdr6bHNeS
kfMtdOw6t9HGCqjDZkBH5Qc2HUbixpihkFR8bDVUYC6Xx2I0NSUtKTOeTdQCa5KZ
MfhWz4FomszH4/OCeURkNwWyuqxFsVEIjVlqFk2ZGnR2vFfd4bk057IawazUmx1T
L4KVhhjGg/rFgcNnGsgFtk/WZAvCYUmHUQAWMEdxwqTzPuso0IR7FYDzJ5qhQIPb
nlNELedxgTdbKbOdAjnMYb84viiryR22c40rinot2/CoxRrn8VmT1Z2MbX1Hu//T
Yki7u3gPD2F4mvIrT5boE7D6EATSvd48+4eGqxfa5jWL3l0NEssc/465MEerNxLb
d0Y18KEMk1HsBqtTwojMOPl2XGYxsc5apOCENhZtnm5JnfMu0HkA7pstF/Njza8d
Rb+huJExf+uWPkz1j0VyocWZ4t4EUAvDzDvsvDKuRJJygZRBsB3fpUHtT82uLYpI
QAJLMSjmNNHV4lJgECzCUPPhj/839YsCP1lLmovvi9xE5sApQwx4W1U7RzIGRN/z
LjYZoGKeyxa9ThOeat5tXljPllSFzTsvZ8d2CdGAa9xzHM8jIVOIMmgDYoM3J9PJ
xiCdixpWFZBYU15QO3f249ZcCXuS5PFlWtamWlIay2VY86M0brqOpepm56kq7Uu+
cJhfIyM3iIsdRvf50ukg3HLcrlVsXnZrdZPqAwSKrQJhuTy7XGckYp/R9i9OuG8m
5+f5gUntHzQshCWt3cZGGZX1759xFfaBQ8ag5Gj2eXzkEs5uZWvMNjkOo9djQkBx
FFTR+4PHKV077NIF1jPbRWZxnWA2sPR68IHWES8GvbkksTiaBltc0nYuy/5fKuC6
kUUm2cYPBXMQ4+jjbWTrzE2dAE70JL1QljTv97dS2Vc11EI5XtYyARrLoFNGaJoE
A2l4kzCTKEthKA1/zM7PngJiPPyPBs4/TgwLCV5bNX9xbeGJ/GAUQDQYluZtmjGC
/3oh5sFppp+ySYAtYF6VKqbQF9i/sVUli0ZQ07t1hg7Oek21wbOUjdvCaMFfHIUc
dCU7IAh2j14GrI6UMYaOCia/rDJqiAqFZ4LfP07RcneTVn8TpPBpwu30DfdRGoQA
ljEPSmTWWtLHvAIyTeZUA6GO5JyqTrKGteLzCdWNYd8Ttesw2veqF4e2yhw/ziZA
54hgm7TAJ4JJO3hbgho0RHWU1wkJb84jLzAB5eTdT/AORwUi5UjeIMkCKRjhXGtu
0r9JJK3WLEWu68RvshGgW5zEAwhKTMfTri6Qu7o1xzxD+pw++h6QEr6R38ICt1L/
FVGeugkbgtrznSEAW6Vv61CoMRiHUPSCyHMYn9aOKNnNQ0CtWHewzuSgzDkzKs1B
rHvzq6IBM15rGA/Nc/9uVBsEsNmJ4Fw1TDLBQSYrSOOqlpHQPV8xTgCKBpT+qd+Q
3H5tI3zeQW9LaoupgwpUaJXG6EHzlMpPr85lliaoPKEHJ8v90TAPoIx7+FOMz3Ec
pj8TsoJ9sby0Igf1bdNPLdbwNg/RuiNV0bujURg0UH7yqTo1VhlpLWAP5jJWGq0a
YztguaXQXcyo7LDNR8oYqfRx+hmPH14CiIwbjRXcH+0pjJ4bVALND09K6QVF99qZ
FCD2l0GAhrq5ID1dOTIUkLe5cm9+PlMu6xay3aYRMX4D9VfogEJuaghzYomhYYw4
YSeMVgVjMF11UdKr2UznT1CB2HBjN/JYYNh7Hxci2XwzX2yyGXoAjVwxeNSImyxg
PSwvDbHdAYzZgxa/+NF6Hi/K2A0bHc3+5QTais21wdJdJWITPL61qcJJl5P+qwwe
p/ImxMjkK6KvFp0+q00/PnHVBac2K+FGgBLthlyAWjiUxldF+MgKRkL6pwQY22A8
xoEUNp3t9yPtp/gTG5mz9O9s/WxKOr3gLlvRsvhqAA7yFb5vwll/6JxLFdrz1YUE
D5+nSaLlz+SVrrANmYc4Z/30JGdlS8WUDD5bY0DOkyr71SJX1UFbuLqTaJp6CSJm
YZATaCT22LPi3+Tz1BsS7Xx0lWDCca9tA7rIDFyaDgW6oWIrJtXYuL0XfSZZtT9X
Akv4l1QAQvO3wQFfV99OY08sAmfhh3C7Q0GHjo3aKhJgRqKR16MgsLPOtm+BzAxI
+a2JR/vBFhBrbbHyVN5LCT89R8UV/jLKCPRGKrFVdA1x9R0nF/I9J6dZETw3a+5C
b+JYa30xXyc2hsAaNQeX0ptsu0//7hQON6i9yYGTBAIhXWiWRo/ki/8bKsFbVoWN
/DTtdnm+Fl4vUVFGR5Zsak/fR8gAFNT6QK8Bph62AGFdQJ+moW3jFbl8yy9Awb2j
6sRuxGwg00t72BTUSPJKSl4Km23r6Ih6O7J+efiMWvRxI0F274aPt4rhkFFzWhiz
5OU1/yr7I2slIFG+ZdTy8Y1nbQWD9vsAsHtJ0GlQwe2SMqIB/HWa4QNDO18nPSxo
oduK2udYHoiigXlmRqVOsRdlM8NnRoA5LePVz76Fqw2PeWvwie5pGyi10OG/R1pE
N/b/ECTJ8SOm1418FX2MJqidJAK7cr5Y/TMJvEh0dJQ=
`pragma protect end_protected
