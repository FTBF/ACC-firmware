// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:07:03 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ItbimE4P65jh/WwfwgCqg6PDIjK0A0RHGrFGyZJxvMNSfqOOiPITWXTLNKEtoZuY
60jgQmguuJe1M1l58p3ksDoLmarkLHHjJBNlKbPXSSTEjKTDHLL4vvf0PdY5Lrr1
elelkPsxTcvPfnqPo7D/S5VkgNIYRmjMBViAs5ejU7I=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7920)
DJRaotHeORT1mehWpCfO+XMOBY7lm5zUqEcran9v6M2m7wa+RTC/h6dQQKIEVots
D4aTnrt7IUB/ADEQDSRe4hypJHq/70q7Qa0ayvSALyORVfzqtEoEaZGp2jo2UlCN
w/V06tEOlDp40GgTF5jJC61E5LtM1aoJB6LxUVo9MI3ePytxPVND3yMHiQboIf3z
6rdI3pJtf1LBV2KiNFFqZ+VlAqeLP3f2Fc/BUdhxIQn1MS3NLptasVB8UuZv3exN
PZuXaTSO26kKMUilgIiXT+OKVuqFf7cIqYeHzSms2V/lfxfiB2yU2HVm766Z6zmz
YclIMrH29zCU0b+nLwgziGg5KmiJKNhUi0QkpTJeUsraqBb6MMWXvdF35IfTuidF
qxMZOtXUiOY0jzp308FqvGfKBC4NI3Hbk36JuAVUxaP++neaT+PxWTOJcogB643E
Fmar5L0xKUuEPGjBzZ4VLuYF3PWP42tosabyy43cRY4JUKaGKnW0p2ifrgss8Y/T
Tt66JdcE3KS1wUQXKPNx1yZMmnDo8YoBv0Qf1O4vyH4w8d6F+qzbRW4fffnfV432
YnqlCd+C9q1qJggZjVnwcC0IH7qHp4zZHi/aenwNb0Hn4tE2kNSjVKTS5/OY9yJq
wV5GQfDuXC0Fc8AQBfSdRQYW2k/KRs9tHLH/CO81gsRM4tG5A67VVCaenEece8rW
/4OR8R994JlWD/NIOnI3qW88Va3X9L/f1VJYhmmuLpVXALDV7QWVl12xDaa4snHT
wQ/EzNAhmgmOQ+DpT+0SBpttb/lMe1fPAvVSADQBn0fYTxD09ybhR2QgdzLibnhz
piwuS8nd30GQc0hp+ecVNVG1CighFBbF7+m66af+v1yIRW6R7WTS9jHZygQVEn+5
SxD8C8W/Q+3fLvhb3j9rDciiKS3q2aDQ01JjDCEOdqvGLapDDXLNu+YBTuNbu5WD
YY8yAeX/R+myLmI1t89zY3V9ytV2cj/h9gU8pcdjrDAIToeu+W4GMzlNTiB2xYSW
F0ItsIzKOlO8JKsZfY6VtYBA0xBqMf6xJQy1Ze7sUS44gepZt7seUUettOV+yON4
tGD5m7N17F/hT6NkSyHTGhOB5AQ6Vu7h2UnwNVIFLySimWN1Uq96FUHHGeGX3Mkd
rXXUBCXsbe/r/cpTJgbjv2FFfL19wJxIqr6Ayjf0uKaSngvyOdZgro+C1K+E6mfP
lhD+UFbNnN/pkZWKObSN6oAFeRGpQhZIM6wy1my/1WxoaqUjax8LhYAsk3T6NiXl
7kTlezvdSM6PNloBIuDkAwwNzp7DQpb5OWeJr56zWKL4Kf+XJLoYDdNZZbSYxGzK
93P12b28ienq00fK5eZf1EXWQ2Pl9MQXj67kr7lTtbQeiE3rTPbo+FHi5tOAs0xi
absU39M90Wf5lRlMgZ5ryUgjjIHwL17y5z71QtoAntnva6Sa4PjWLwBWANmogKOB
cp14VLlntqQV68WiIZ91kI+KwaQ9CbaUVxoj9Mz20zakoYhgBBYkRecmuHxnXVC5
YxC1BPQZEMV3YWd+G1bNJps3yVu6W1DS4iUKv9CCJIEf05Ir8ZXCWgzt7ovYQyRT
MXzk2mpbcZSR2vBCM8HU/0cxGWBUoL6MlXinK1V5gXoSTmGsyYdg6JKtagjxiP0C
5wBegvHxxsUTDO4dXfQMnjccB88/UXaJQtK0K85i60/JnH36FJK+5iestQpx0qBb
B3/iq8UTlVZAq1YBfDWbbif286MLE2Xaq9zjsaCfnL7mH0iCbOzphqFQdTa2Ly20
UoYL2ye3xHj4KZ+5WuN8i01CklN9OPD91bcgvTPuuSojKVkLaV1pbl3kiGS9JUlo
GtqWmOpBcY+PWPV5NAAnSkjSUgmQXTyKJACaljHP6rmX9HQ3vPWGdYN47nlE4ftl
Z6DimzryoONaGONHjDlbMG5wvuoLmQIcM3m2vtdvRHiPkkfRFIR0PUxe5pR3BtRA
+lBXs7Ctbt5JGvDxQ8UMYBcYNbIe7QNiaXTcS7F0P9AUdIemL+rl/TaNhwmYT1PY
JCzG2sk8SeUK1rtvyoa7i2rmW7dbtV1Lgh4dTjXj16qrNt+NwrpJB4fGoFm460gY
JMKHi+JaRU5kYwQnnPDIssP2sElpGhQAuO46eoVmHzQULbcBn1WeL+JrFN1AQOoT
Qcn5CuaZNjh0EJTl/RURVE47Nd9BUmy7I27ZfPGmr/UkUVuTtP+vJbysVbVNhbVQ
IWrsOyDQ9okIMXZ/y+Xej/eXcTOgYNVsJUbEZ52QNNIho3GUIi4ubf3X0TW8pjtZ
yPlIcHhvz72l2ab/SJr1pJ4YFzSntaEu7VIqTvFN7Y+DLQFM+W220AWp/G9Gjdy3
ugRmabi85zUrbvOS60a4zJFM+Zf/is2zB0bhtRyMyt3C2w3OK1JgE29k9U4L0jR4
XCbck0RlEexPRXRVyIyGX1fkRdD70ECO3XGDawbiqkWcH+fMVFJrRvJHed/i0KXD
yy67xie9sHg1+Lu2jd00In4onI23xRTNoq2sjMhsHUpQjSZ+uS3eTduM4bmYgmdO
D0Wz/rFWELmImW5udY/t/KM59Y38/vKJkuK2VKVtTwrNtb5ahQctYNvTtFbktJ7E
zYw2HvkT8kWb1kfIbWu03HKHZ9suErdVpQihRGGwwrqiqQhd6dIRffLnDtk9f5jZ
v3EEn+VuxTFlieF2Jr6eR+UqoVpLb8Ws5A9Mio77YTPfn3WsG4Pd7s+q/FXxw9HW
G7RfM5cS47PN7v9d3l4nimfwSfKMKTha4mi3LwEsD30m/npoGF0MhyU2Xoy6XdVe
0sA2lPIQK936BmkPIEUnC+dESJWXjuhD6iolLD0M4x7QHsksK444k+Q3QfMopNT/
dPsQ1bXumG4RO5jcU4mFUpjT6ON9QSgsVzlyZzvsUPTf5m5m9U2ob3oUkqgD0TlB
vnCh0hOcF6SrSKIFYnzk4GIYMikC3+DsilqPBjPPbXzIs+3vMOVVoPWUKo0kd+VH
AOxyuMdvGvn9BSRipdUmDxcvvKYHLMoSkn8BAK+qQDwikaeD2EaaAioyP1Cqf4vF
zMQOk1T3yu3rLXWe0WvRb0+SDCf9yZ3aMktqAp0V/xbBLkTLrtrhNNqx3C+FYM6S
jsIMUdl6JJMoAsCD1nGsrLIp+FzHy1mwckoBGvqYcFOoYhIoeZ4lx/ROb9kA/uIH
jIzUM715jiIpe27UFL/J0C+1Np4gYeSgkZz3sHZQ2tmHvmaXxoJU2Ks+NZnOG+T4
PgAS14ea9Nt7SkBV4x0qLjJckDrfA5MsFmAj5Nj58ujGyKWyu/P+aRDZccLqUfNF
fPsjSkk6OeleldcLQWkpc8xKWt8aNQi50sDOi3zS5g8B43TwAw0BrfvdUaqy4J0R
OsbBeC7RRHIpc+WZk/kQd84Ci/fwzWEAT4o2nfpsK5Fj+vkYmUNYvTjObMbFFtlE
eTUy9mdKEGewjc66FsKWxDg6AXf+s3Ba0ydB80oZqjrqqPfWC9nnzEcEYXekGFYq
C3ez5N1f/j4QT/CYG7/DQww+MFhEIwbyaBgRZUSCp3X9vO6Ti4pNH/D5/b+6wh9I
8StEIYzZYAYq2B+lPeCkkI67bxgxZFrS9yLZfNO16hP7bUu/9NLKPf94336Jshrz
QfN8toRhxj21baPABOcRSj/5hVV8hBL+gmJ9tZSbKYBisgkRVF4w9pKo9pEjK4W/
iOrnHPTeaXZ9hUJi5CXsOqnD40rmrp2BnnXfrSEVAvc3/4Y8xp2TYwkLV117XPGg
Y8/OsLrYIKF9F3+g9Bt/VHd3YUVf0J8fxu57oB/iCZLggERSmsnIppFSK79mI4hC
XxHEMcRGtk1i/JDbLDHY7yncxhZYyQtTjlCOwhetIa6vgCk2k/Lejr/lASYTOftr
h4ojgt4FTRESF2YV4U0FGi/HsNanAOdOOfnf1RmLvl1esz+UgDnMBiq0S9TiOISS
k9N+OrIQOWFNCPkUlUEiOoEkkS8dsCK1QzCJ9Opz8MKr3g0PW8eZ7/VHSN5CQ83L
Y9xzQEX9fIMbx2q0/c3E/S9GE/r092psuXaDltvfAG5VcjmQdEPxhOxAmgApAcLa
SrugdX1PxQdEoJnSANLJ67z1THa/sWaCfPTe2DoiT3L/caSMrIAfKE51+FS59xBW
rupE+M5c+Fzuwd+NxkaSKOth5xv8KzCgwZcrTtU7tuenDbU5YCjhYw+qTrD+UnGR
D731UJDjMjvCgzMDR5otnvd+60k46Vwt3Yxed41B7VoI1lyeDEZOeUOUPkIKIOB2
yvOCTkTkkC0qP6rOi4AeqBeZUmCuoT8vMyDF549y+ES2DWLrCMeFuyOC+1Fkp31X
q16WWT2iB/TCN5W5f981lJedcT58ncfO8S/0Fp6n2kgIMN+w5ZjfhvsDaw0Lv88e
K3n2bFfj9V5OFEW/5wBQd3KrnfXb7zr6soTcJ6oPoGJxpibXbyYUUYFr0ROZx405
hpGHgQ04820j7+2Iu+Hwc9Rn045m/hHLG43EVAGeSYJAAbdhyLcmXm6yFel4VyQR
hnMcIzjhBL66gMIpTmRBbUuCAgNLZrOfbNqF4JUJCFJDwjV211Jmse20jXhF9Ah2
LXJPnCnrSvDROVWX90Du9T0vqm2/b7Fu4tl4vu1Y0PNFL12tKyjer2cTLT9Ox5Bt
SZSjWIOy+MjIcHqkKY/OaCAwB+/Ev85+pHUWFn6pYKSAVuVzWE3XsB0lrvMAuWVp
722yJXJuhEwc8OUVtLq3+hDebHjiXUVVpQpx8k1/hHHM1C+ob5/tiQSnqLb3dD16
LdJvef2DFzHcypk+0018q6rxm0PMkcLmDa/0+kwWMho5B2gAdW1rDaV4NkNHc14r
wsYlcZeDT/wnIufu2CeVSjORASWOXbMUirXqpoIYBfiUC1MJw/vkY56F0O5axtxW
mkLCAr5/wHP3YfCA7+HuXzNWH9Mbt/+bjo3CzqRlCkBNHXYas2U9xwaQdN1Wpyoh
ldDEjATpPoiXS/XoUDraxc4jxFkL7ihmM5WjkgRaSq0ft+gLKrVV/u69iWYE2eeO
dPeQUVS2lwc5Nsd5KhUYjrrmUvZ4HG/CjqbhrQ00SVjS1Xu+C3ah4+W57a3HJSDH
DtWCI0mp0SOJLjw3gt8Zdb3JooZ2z6lLRNagluVs0V1dXqlFZyajdeFp/t8zAPep
ccuTiSmO8f1bUwgh+WDYl7CXOc9xtTGkH+UTbkT3eRTEPEZYGHXSCbEz41cFtDv/
ZheNOBL3AVm113QAFlvinlGm6Tucs7kq0bsNLO6eRXtbkTqtgj8S9IpsmXij8Ekk
KGCF0mMyjlpkHZhPexoO/mXxoTvMRqS7p6D6TEJadNrCDlimAgJyNyncFtPQjiED
fdrlEH3x1uTBVEG5cYztpGwcs8kCtod902wiRsrPJHELUnFMI5qclvFwX3zLZOKW
PPL5aPSC4XtUqoRJGZFav6MFORubJcqpSCLFRys7VVrrvihvmrHyLgka8wnjS7d6
37Pok+ym6sPZ0RUqwRRxT1IJ5fu+1SLGP327Y3i2ljNkyclo8x8vxO5BD2EuJuji
jmHE+R4qrm35sf66RkldrcWgofx15V6ehcV+B5iZzcZvoeSam8706X4yyesTbF52
bg71qNeA1hxuMMcsmP3kJdksL1iknt1/iU2a4tKU4F8T8yLdSGWUXW7WevfaH3LD
QFvYMXs9RQeg/z+Efd5kNcvOsVDuMiA5nnNPxg0d3/6GZJmv+2QZl0OLx8ZyAEkC
jmLlfmZ6wPxsvPXyQ1rq1eYeqKZMqhHQ740OeXuHohTbZKwR+cxY/Qi1j5ZWHO0r
96y1h5HKBizjMJ+ZIDGA3nibOgaBUGtzt7cVmdE/7epIqmY3wjkjADjo0h56paOB
mLbmPE/YJTL34DCXj+FPdmAHNbqy8pRV4XfcTKRpXmnkfhu8CkDIbXDzqP+tcLlC
pWbzw1MDyen8mt9kJZVXOGpT4C4Gx/4dY3OyEyUzAsSqzEid7I9uALHsechc2Osa
FxDLnGCKy6ipmns3nIwU7IpaBSQ/gG1oMWpTx1iPgEtH5c5dJgKZy2a7p5G2Ec4o
bMx6HunCt9eXcie4mftdtt43zSkDt3MIPUregdfevQ1dzRLfBicyvPHTiTzP2wKe
rGwuZ4MO7kqsBAfFaEna6WnHrlpV+w+9k8eVGDjdOGk34w/zodycG5Y/khVR2P7m
ABA1AtlRbvF7bRefQQ4Jd90bQwDIzo+1ss3PPVYGmoHVkhLdLrDAVNzk6CbaoZVD
/zXQCIUqv21jvznv1ZtHdugziPrGqY1LZfmFKuNdRU8eBhoq9NEKNrcBupodQTE7
8uo3ZTu+d8IyzrqNqJ0jVZY/vx8aEJztVO6Rdda6IWUvXCgiJ58BUfDQg1PmEWJF
dkQgblpFhGTh4ZcmeGC8vFQ7ZrwFintOfOcrtqCF40GdAz2I8vzEO9kby8GiLTDp
qUoOYum8gYLlw1mzLHqH/QbKY/y1soDg2pkY65XHfeffx8P3X0YytnmB261MnQ4h
nBcjHJeceSJ2wdj86rYKmM0GhExpe5W6mxIXnIVTTHVWbO5wizGSFACbMzFyZRcW
XKPueSw/qzwhfPFLsnNBBCV0C/vls/gkgQCRa37YJsjDPiF45S7DT2F6z999eGS8
YS4mDY0B3nP694cl7bXECq+Lfpou11yE6OU7wAcCKpFyD+ul0eBWU5e3KLp4uEJq
7E83Z02fiPofDt/ICANXdsnIbmTqAKcDiyy19O3Ae3kiuPUMhTz2fv1vlm3Mch89
IqtaPCkIzJ4OjbBMTnYXa17rMQ0Q87HAINVd8hWvgylHSAk9Y4lSpyCWvqAWwg1t
rlpwDZKPGtQTzwpkvmKVERawgYFEBx3XHZjrgWJaDFztaoO24E1DioR2lnAePDsC
Qg7N4yaqiKiJk8TcIpqBXTspnVFxPtDvQUL+e53eQSrYApfnDs1SQ7EHkREhdi+y
LL8KC5B53lrdZNl4RG8Mt/1Vwqx+9givSfCEzh6HUk8ONXpOOCfElBdCpi44Ghrh
Uu2H4W3epuXJuNOQhq13sxhvjZekDpA4bvPFx5eI1xeGTeCW/t5cgi/P8FCV1v6o
79ng55vBrDaOMXCcWYJ+E7ggj0CIeKd3knCLZL6tV2GrInKowLYrOTvU4u8DHDTI
zFN1rQn+U8T1EUWUWYUVOebo0yuK5vPnarpMqS15948YRwonOSUs3Lt/dykoT2Y1
6E4qDVOiVLKIHmSItPgNREA1icww1kq7jlGKgCrM3GR/QQ9D/jChFJm3RClx8FC0
6CEH23ZGBARzrWkVTVKCQsLmyjX7NK0umfJZt3jMtlLbjEjfBpxCdm3nMJ+LlXC7
U8IlsquMlkd1rjsnahVOSpee4QzK3w7p9HPEUIDjJTDpk8ZpuidBkuLNZXMJFQYr
yRMJdN8X6lGzbm3u4Zr7q+kFx5mJ0fnNLeEQN9x0pCD9Yy+iUHgMrinZnnUf46rS
AOK5teydobpn7Ou6Ce0akO4atlAsdgE/hdsFfYOL5mzR5fcfefVH2mzYY7cMbbId
vWagLhKSEq5anTRGz4cQsd2twizIlylKtTEcJ7vL6M18VmmDGfjzeGwhEy15+pLS
Wz4yXK5At7gMZi+OJksv9w/cubqeKqMrit8PBbfY2P4nQYBKodDhJEtmkSWQW6S2
d9bZl19uchb37m6N+pFQEwFpQwXNMfS+jMdUalAiIUOnntwbf4FqHILYcim7E30Z
xCGhnCFJxnPEKAApNIowyW9nOcSUbOKr5qLjbTzAJVkmpVsX5X6HBTaCPTrHZRiX
L6sIZZHcGfYzSZmgVeS3WnX4tgHJ6CDtdTagG6eFbHpmll2OmRujAdqEqyR/Oll4
7pB3pJSq70LEVwSHL1d4kXcOhzJ3CGYrVK7Z2AbpvWH5QNoyZExSO29/dpTqgtIO
JsJF3TKk+mO0QhuqQ6rRQgeutd9HeGNfgu/7lLJufiNDyGgNkRXr70vhcyUcMWic
0/lumLRNxyyHajYhvzLOPX7Afj14rGqudgI/deKL7czTxMY18w/Eg3Yne+JpRx6p
5br48rLquuhUrn8VG1rwhidtCHwaQiabjsl0F/4Ep2H1nWpQXmcxN70vG3aISLTh
jSD8hnh0uVWbsLIqns6kIfmZ8NS+3fH9tY9/r2m3XpUvXAFGWLwqyStWzh899mad
YyO8K4LeRaEkPaxuu6hKq3ySBoyV0lUxm/dyZ5FFBcTeWLCxv3Pvo4ca9oAnlcRo
PuKB8ILgcxeoKi7u9TV2J9d0O0n67XlSkY4mqhZFIhtIi+4CQJEAgI27/moFMyZj
egNteIsVd7OH4lGrmKkWQUHHrkrbhbwEUZ8vEojqjiSBTKu9VqeOCoqyvXGvs25p
UwvQzXpe9oA4H2v67UBqhlct7fed/suBODgMj2c3YMGj2mFcRwOGVTG1/l/Tor13
Jphtj4e3viGq/VDd2UnVgQNV7wFt1K3Bb3feXlA+QNiNA4qt1rD/H1ZteBC92oTJ
rhC2KRpVCJ80HfeVQ76OWDUn9TbV0aFDEUbe1WEU4T2C+aX1GPeoi97+EBUeGEP+
neDqNtKuhbXWLGcotfai4/mOeiiCdbDvXuvqIgoS0FtHmm8ZHp5qktDG75E648Vt
1pYKxA7WwA/JpSw/gCoiwvFpbevzC3fG8B8VhA/qWJykEgKCoGIPB2bHYWuysRkh
9edBYRBPEL9moTQ4sA/EZj2BAIElR8r3K8TLT6Uzf/Sr54fVGgzSH7wHeWfLRgow
/4AW/6V4WlMZeBrsadj/CQATyo/ZZIenRLEXIhpSX0AyR/LFbzo8PEIfB2maSBPS
HGtRSW/+N1iwd16DxzN3x5sutTMpZ9MMJzBcbmZ4cK9BaP+RnZMb7cSPQwp0tZW5
YbY2x/hIfbVLmO3+Lircy7L+TjoQnFz97q1NZ6A57qJc5X3mScc0cYJkS0IuVNy3
kWlfNNO5NtVV6ZiBSe3yZ/JHCQdti+fK5Cic4cQZjFOb9O7Mo4tzfczqQRcpzLmU
ev6hJaaIirY5iD79aXFvXuT+xtdW/53wr/Q8NQwNWsV7c4co026lDaKcSGs1crG4
/7iAiJm2DraGZ9jNVpNXU4Dj7eVk9YBPYMeq+TliMkWvpoGOEejYH5pECyC+R7TU
VjIhPodBaFS6VJ5bXKDVlFUIcjtbU+yFnzKW64XgFX1Q/h4iPaZuT8bxpL4ye3k2
5+ytR2HdD9n2ZmCWtyHrs8LmmynzbcMFPySIHkgz7YPx1Mx8rGNhP8+AK2iJgvEm
44bxdK9EeZ5K6gD7aGAfvUpBzwRIg5SJ3zXXsu6YXLzUWamcd/ij7kuHSY1kky77
qcMMKz7NrZfkAtF9GE4utOr+WZSWXfigkGM9tjDKjnUoLSRhhYV/VJT+biqhbm2i
KJZ8uaLAh57sfGq2YW6E8o9WcTlO8KHGr6hiVkpLDmtgwejYtQstG3kz8HjHQfy3
9v9rrNefwJyE/xOeQCYHzQRneuNdQhTsCqyu92bNXcfPU48AcUEFOLo0MveH1TvS
Aw6So6vPhVRe+kt+mc/RasiJnktFcyLeEq+VrETbQ6GZPrsH+i1mTUhoQzwbjQQE
WRSLClrnpLmJUL/Z5/qIQZVq5Z6+Isdf3GTwQ/wy4UnrBPni3CeOLF2a6dF3Wlgl
UknYDZ9msTOZEokMIdQt2n8jRlKNaFvmlR2oOF/J0BpuBSHcbJEpgz9IZqbrAyO+
C7hhNiy1oEJuCl+gdG1uc75hlyLf2GY1zWXFP7bPy+jXWjKVzbpNgbP4cgiLbYkO
anyK/u1+HuEBdsqGGUByQ8s8y2pLZMj2peMI/U7l+mNQNejyD1i0+A+wbD1HxfgW
hzczJL7E697m3U0cE1JYSYLEgfIQBaHbBFP/x8ure4rT3QNuozfR4TDY21LcjsK6
QPsvIAHwz+r9V80C1+7mwFy+rL/NgdyGXOn4N+xcvGnZFxCVfSaWLKktfdLCHunp
t94Jl4rJnKIR5nnlaziOOL3E+i3OweuRGn8XeCAC8dWIjGg9OqK5Tuz+zXDSFFMs
s8I03dM+H41NLp2hM3vvfaBRo1+kaTXQBOb31fs2+LgXW5qZkPp7kstAtiGNTpG2
op9EEVjmKpKC5G7YMD11vtmFhTH9RYSrykeA7RdqXAqY9mm+yCRBj66ZEEO0xX6R
VPzPSr4l09jrVrmxc9PiS3ywaw/3jG8GPFklaIlfM6EdFSa+lWyqxZaBPsZc+TD/
hGWE/SUhupi53r+2IitcTJkaaDhPy/yoPV7B93aXzj5KrGORGvrFYAhoNisMIaKT
WnO5dIhHC5KTwvA9ARy1U9DceFVfHTw/y+tQrSyREGfSUqg0OMWvwpZNtUIsYaCq
ZpxSoARHQSLdQqKt0kz7FtvukaZ0RzGJAHFFeUl41n1IcdEbWu7CemPobft+bsNj
3GzDtzyVrkRnpEiaylbrttRv7vCZmxXxGBJB/SfUsTVxC+LSPJIS62uRgAaxnuQQ
7BybK//6/ZRNkNF5oeVywN6hVK8cUbZTR7SZ5/tSC2Os+l7Unpmau2Wb07n4UdUZ
`pragma protect end_protected
