
module eth_clk_ctrl (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
