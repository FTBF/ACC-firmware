// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 03:56:42 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OdzoaPI68VkqUct3gyfi8b6+oCZONklIrQbBTTvsu/nF4volX9FvBTC4DJuFlXB7
Vl5Q0rlpm3PSo35BRyI34oDf8goqF7MHRnI9Wzi5x5ul3pKe1kXa6vL2PWCVWQFV
3bc9oF2Er1TOzUoph9pfFZcvB1raYqgGTrLayQWaaPc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7696)
7atV5/PiRG6BjTgHh2cFk7OI1vrDF8/uACcc0+7IBixA0eBoXpM5zKlvSsjPObaz
gYksc8f2jhWZ9+LCt8jzKtKvmL6FkpGiqWa4XS2Q7VeaVCVIAA6ZeVenw9LplqCL
le0YMO+JjdJykt5mmU+GDQa2vsx1ggcp6w1BBQ4G924tfqpSRdxTIoWnhDRE3vQ6
esYTZR2TJzVdyYRK2o82sEg7kQPGHTfK4FHLzc8NcNY+xcMNQfxciQIGWYdxZ2UE
ihEH07RjX7y1+HHSQcvgzFDLYBExNHXPQrd2RVHiKonVO4E6otoArCKjjN/iasKT
ZeVaBnYaGXafhoc+G8GL4xElM5aSxBPu2fFePQEzczk9lGGLl12pE5InKauvfzUl
HuyHSyKOhGkyG9jxAa4d+Vonv6sV1y+Hg57a15tb7lAdkJUdrObRu/FPmM/BoFVB
ce3wMIi62JmKHxx6COk2ovgp2dYvzAxH7ZsTfA1ppkB18s1s2YlrSREu9c7iz0v7
EhotfqN9lzE3paYSReOI7ML0vapVYqAmFnocnvE8GYEpgHn0EvOMy4Fa8e1cCokk
P1wlSaoDKIbjBdbun5ToK5d46CGD+/5ta3al4wSgWmbmxizSOodYYDcK4joparhM
LOAWuKwxNE8QBnUm0xK0cLmyVWw5pDkxTNXSncGh6dc6eS2n1odTCbCHT0XzGIvE
9XGNF/8oeH4KLOadv2jFx8pn2xa40QEIHmeGtGgpfp7Cb0t+zbzlOne8hzd+200V
9cONcmbVAUBtWF9aHNrrr1u5ihtZSCnNfCexHjDlzYLzEd/JLM0sVcwiV3Tn9OTI
fyjyE8c80Q80PXLXQj6rU+fio01Hk5XmPJZJc7hyz3QfdEUgXCLzNnsrqEanIWTS
02SHvyOs3xJBkVnui3Djj++nrmaDB+Kz7wmL84XwSvTBIuS+4lQuP2T8Uto7sF37
uDYaIihDi12ceQV4yI8pBlN45fRCLgyNHJEHS4oWen3MM0Q6boi1TvGEgLWC5HHA
MYzuLPmjkphLWUqSxi/lLrxi7La0+IsYFxXaBJKjrpC34vRh9McaXTr8gW8GDzpQ
LsD7BbWLvfR4aZPfIBl2CiJYtxeTf/4RLahso/bRjpv2ShIHT2dg7yCRKP3d6JCH
ByH+QDC4aszjKOHV4cWKFFss+kQYsRxTMe2KLZ4jq0xNF/4zygZz6mNHMFuj8ziU
dTE+lct9di4ecTwc8cDmfOEK4iamArzPHCmksvUSX/CDYlEoxRkcMuKY+L4J/fts
4nEC3uSTQxNLDYgIi9DL2aI1Tcl8AEoTLSQJW2KELSPmxDP/16laF6iyV9FyepSV
lpaAGRztvXZYaUUKgHN32ta1axkclXR5+JpwTYTg7Fz1pCUnRYXBUJul0jSGyYNf
AfxTnzdF7Ou4v4qC4ix/NkfURt3mQ+XM5gWg7Xg6I4lLLbqmltapqSAKpquAUo4x
+HSeUJ2i0mdTYcnQ7OIIaRHW5GXWDKZlzQ2VqHXfXaNAACufY95ssg6Fj3blp1i3
fOi4+QKOc+jU5E+SA58ODrXhQ+iu6Ykkg/+1BYo2SFAwMnwiNzmyOKPSQyydkA7Q
m+XxwSgOzs4Oxf9debpqUeER1letIlJQls/BRB2bJeT/zaj848MfiNibFgYrMOii
RIr7+YsVu5sgi0REN5l8Kf5LulBA+zKY1oKs9PnGhEJwKm9XiiowT2Oz30AfWJN3
cOlcQhBN5i29dcbGIplrvSf3P0Tol29TW/1E8t8dipbDv5vEDRre/Tnf8vehkMUc
WsfZ+Fd4wK7gfD3G8A/UUyGWP6fbgeUxe18gTE38q6UcAQw6XBZzsJXue+PZ9x4J
QKfwT4sXLs86CkvXJAvja/EVMlrmoefS6GmHC8AKkfSeWbEtuy+9qIKgfzkx58Iu
Ocds/B70WSIeFGU4+kQFTl9OhMCCLZr+z0aRZctgDkFOTm+p4lLa4deW1OMMeBTn
kUUPsxYQxNND1y/CJNIRMvsUTzSMKIPcT6lR7TFEV+DP+9Yj9ubRD8aJysvvV+Ur
4EZX2csueJAgopPDE9/EyFMRO074A3bSzfh2JGZNF4IC2xIvXYhO70aFn5p6LQ+z
0wimJfva7ZRjYUuIXyFfzQ2gKkWdR3xQyj5ZXtqmrm2nSx0GdrypwpD7Wi+Yi3+H
t1SFFZgiZ3+gwpzHH8Ou2oupprVYqQYh80yV/wPHGNLOtYUTstOUc91ZJpQr7rrq
CBLXVEesYgr+WqKdj8+JlDQ85eN4GrV7JXBg+WKAroEJWjUpfkZrvGbbp65QwXlU
dmTg4ABmOr1Bz4fTA3iCWd5ppIFY/DEq6GtMqpCroJWFKetg7qKUdAz0f5sJPzE1
rlnU4CAugXFMz8u8PcYOiq+6sA9vdlErkuR1lZojdD45ea6YtbCa9HSxNKFfuEmV
jG4sVz/dfkU1iNJaxgucW/Z3Q70HbkIuXhpYUaXyAlvvM/Cj1DWJ8k60/murVBu4
cvelc7mNMFxGdxN/8BWpnqa8BnVZ3nb4dAZDIS7c3y4vxGY+oOnT8Wt5YAwP9fY1
ASaLwU73qFyAd3heVT2q7PETmXeEElKKpuBwIDHDqlxLQzKUGHPnyYptN7T/LseB
Fi4SVj7bVdFrZg8nqTw+Bv/O7kjqJ0iKBZGueZNICmzj4tYw/NOMubqQUiQ8fszr
PW1S3/EJsdo3D0VvphJPaxryYMO2r4LU19pdDWJ2eSEF/+IIW2KpvJ/Ezz+T1S34
7ffglQ89MJcP/xQdgGSvJMH3kDTUEtpQ9T3kaviAdfHBPm8MZ22KRDVllDdo6Wxk
F5zqeIzf/cwHTv1h/i1BSj7R6oa56dfXdEfv64UhJ+/q4rjRdF22D2uWv8IT5F6B
USvAaMcY0RHf++imw7YiMdUMguk0raPx27TCFbE6vUayPNHRbxj7Tc0bCQ9mnDig
3p2S0EzvvGrHmapsr+TFNuKgZJLkcpcwnihKas3j3DGYyqqzGKWWZIX+xclqd1qA
MlgZKSn2gazD8lAICt1ErIDrTrnmfcsLI/yfjt/zpYp2QWdGlScb9N5MWsD9zpI8
vQKWHUnEWZlCGLWp+K6+2QKUE24/KvBZy9NEYyXCOfjoCOyzJivbfQ9g6aNMoMtk
VQkwE42wDR3euUi9/rGsAy8f+Akeswa39Ejlwhmz+t2XWK0M5bdiQ0fR8RZqvWUV
PqKt7mC8i/R4xX6aFZEcYJEK+uM6PnfkQ4QcUVsJ3AVmslqFu3y4eaQ84RG9p/Mn
s1RKy0qXKEDp3ZkFZ3D7HV+oFpwdaKF3SlqwMChatauFkQZthNjO681myT/KvsBs
AX5jqeeeTO+gkCEH5U8+moB5v0NuFnAgNMp1waZEprIDMENoBhc3hO4BsThvG6+c
Z0wG2QinVwFYu8nT6LZ9fpqvQp6OL/xxvPhGxxpyDSS4rGCZGQ0lN3DNhaoYrxe6
AYzyhQT4RNHDeBKBGoOC6uL4vKURv4jmQ12XELH+lUxc938A4rhdK2fxwG41RsyN
BMifOB1qQM10PvvgvJlJJTrdH6FqlYgnC7kdi2l37zKb5RlseSQZWfC+WITq9Ahr
setfSVK16LSuTiGwtAFCB9x+IFUbjIoNgiH7URGnJxYZ85I1N9gicMiHxvDedKxY
DPKkVpZaEZGadIF8qGsoA8fIAvVo9+jjjdoypriXtw6FKXoVeY2gb/OChbZlHAtv
qaCdRrkeTWACN6cDJOYB9P/Gg/HhFc8+7ZVhblQ5sXmzdHPDt1voFaSSZ3IGk2ha
dLeO8X2eZ47uUr1cznITTCsgj7liJsyuwaEoZf1Wa8eOz/KvGIhreU+WIMb8cUCY
afPKsPtNoXdcWhVS4/+w/xDM/Mdpg7/aivJ6vRV3/gGOI2z46aN2aBl9QLLxIgKC
iFlgl8jtJ3LepZCPtPob608ja9MCgolVEVGr/JKfdkUEWLweKPjR0CMvBDDeBNLt
RshAiFrZvAdMESfMEpbEv77q0lE4rIkE3zmtBYWxqHc0ZZp0dDo/iJ7aY6vL2fU2
rFXeGbxYW38kfUj/wY1uM+75ytU76vxoAOIaRZYO0hfPLBWkhzNhq2a2heuqrGQc
jqpAhg3/m3xKWubH1vjZBI5pXWokJMswWeancBDloAzUWWyxqSHj3TntEraKWjC1
BQBRWNUjyCkVXhO+FvGw4VO2f0ZRdWhR65/1S2mD1StkJPvkgQ5OBMq2UgRBGzcV
0RBa8+rPP5JDL0ipI/1CZCRUKQNw/Evd98yRT8SfzWKtOIGYcrrdlR4ZRncEouQv
pgpcaHh8ZsZ1+oNNDAYQGJLCu7a2V80cyEcHIZm+4XMtqmtuSPHZyNTxG1Utp64u
O/GlWwuMTAwcJjlKQwHJrbRk1K4SNggeyGlLEJyY3knPpaMq7V87t/10ozibPiWc
ckXIRFWx18m99OkqXUKUdJGe96F4OZjWSprd3qd6i1TcGamss5tbXpK6y7Yx2+jL
iVyQ4UmX/jAvS3bP1cruG0QwQa2xlTe39Df0Lsgzdf7X3Qvb7z1PZrzjuQ868fxj
cVvDfQByalrf2B9V6aG4w5+EOTYJNB1rx2glrmxbBnZKE3SWr4EqMgMyR1QyJOK9
U+AWeVVwrX6kBLKa3N7C4TuLmr01D2ZXaNWrE8XhAdZ0EmGDu9JJsmaZGGl6N9m5
fpR+moiIr2EzHEOBr9g7u+hHdtcA7i4e2I4hd7Vgyv5w9JKmvOFJ5asfxAAsGArr
11y6wFaGee3YcgcCFXWfD9S8T9GC6B+KJZTz6vrOQrUYGrvtk8my1dQQGHFB9nnO
e39OyUt5tQKprEmgsdrxaO2OV3NeN5me84UlFu5+pDRfrOOrWnBFJl1xgNcRrrRo
q7yADPlQHK9OJyoU2mqpGLWKYd5DydMnOCiBqnU2zGKCPz4F56il7K8ToZMxA9Xc
bsAoAseR71lcLRLx6G/0jZ8nxQ9ukSYfoEcz49zdqV7fpt81LZ/+2GYtOw1FsWrZ
mu7uApaLhBFqGREAFrXKEgQwUmsUNrbuBDaiiW6zT2Fpy91/t61IJXOGPdwfq2ML
QOzuST8Qvaap266VEz83hrmDVO4HqLnIqg70kvBdlQnFWU3NJJmpRX8AxBRnoWXo
aLHAV7s+o2lzBn1lavA4LFu/WTKixZjPmGD4C4NvjQMvvPmwQ9+l/9wlwcxrXto/
vFhPMxo/FLVg3vpjqnx0D9fWWGtAckqQKPOpLX5kQmEElTA/q3w+U4kj66PtosME
5dxak3z9879plp90ACvE2LyN7JMUYHMcgf0J0mHuTdZrZJdtpfS4wAP/8Ba3kuwQ
yed/8CoHG5w/QUlcpN1ntdtk696yzjA4wFv+hq+f1XHDveTOOlAyTB6TdkqG/UN9
jSLuEmpJxIwrbDuKRyFcJo+0JxYX+MOzBrMg7b78iHuGoyfoVH/oa+YCkqEObsJM
JhmarWCD6JsDN8lGE71QnShPKD8aTVTNVRJUKfs8lHCT35YJiOs6zAybkrQXZg8k
5mjK9mu4yBZRk6cwHAOOAh/gLUHexzh2YL4Y1FKU36rtzXOnguOtk4Yj1IFs3fWQ
8OQIUi6I1jVJ3qGseoCuD29cECtWouXLpoXwH2Zo8EMbvVePfE/ZbnFRBK7tYKdb
zR1WWJpwC8TrulxUHXrqTrRsBesyZhkDDYdgUyzuS4fp5Jn/tCrvLD8yN9aBXK0B
wmjb48PuFXi0gyUJnSozB24oRDUEAcyGidAAjDXDB86YMyH9G4Nsr7qMTH48Y87J
PTklngYttwaQ5tzFFErFBWIdHNNQ2NZhF0BD+T6unydBdVxGvHHOvcPvFWKp9MjB
psYrQZ9I29KJlR1cH0url4ugtarzlsAed2zOnjqp8mYJQ9T5WEHBjnFWuOEHCJkg
t8UIpBGxU182pRpszrEYBXlaQybB+i6uwXmG6syDE7ok9S+t+JT5FTsunNGOBTpM
/uMgVEvuQ5DqXi1iwi+48zKE5Vj/zvzGVXJnJXmgy9N4CDIYd5lja3uT2VUuZdOu
mueunY/Eo9vkdMWPDPjof8omEFXZANY7Ts29Au3QsgHqHttFtCWFA0x9lTI54RvC
d70dH/yl6pa73OaE+WUSqq5aokSXeBHoWS3+36btGSyrHvnU4oy2S1Hp4PPo/Pnc
rnVV3bTks9LPhy1R98XegTch58Wx2yOGQrnHayTKOp8QG5QuaU2tpGU+XdPKLgmN
TRb0ZsHrgMSy/Cn/qPdi0ZfWdSH51hKjDAU0nLhxHT1kFmj8l14GdytWJ75V6K1w
Tk3im4gLA6iAs2UYzvdCGxA8IvQnYdWsR1BU7vMS2EKaNaOi7ew9TDfstqz6xbsu
NrxLofOcCIBPVR1MRa2L5PnfV8YGW17P36gPbKFJq4qxt4tQpZc5lVwf75mVxiIe
iwFcma25l2sv80yDZIMSUdmarLpV6bOtU4oF1eM/CB+CZDgMON/3DFKi4s4M0TIS
O8wFUg+h3M7lFKRYF7tbSfGcXUH13teL+cPlN6uq7+jHzbJm6TyiEJL+aYB80OYu
fUio4WSrRXNZ6AEIm/MFhhsx6IjCnqtqc2WsZGNja3B6RiZbaVJGAIIJaPy5xQg3
FPuZoBDHlqCHC/GW05Fx3gKbQOItksrmGnDZe4K+XhczFZxMEErGOiVfxUKRkwjV
5i2fcDBG1734cQepo4td3/Hlp/q0qEnb5Jifj1uspoMtl3mEVJew3RiOICwOL+ot
2Z0gkEMQ5V4eMjB4e5/ew8V6KS+VKNssQD3tp/pLb4Q14yZn6SeZAJpbX24KPHli
Zc5Smvb8UhjNnHhPm6THQjo2xsZWO+qpDo9eO34p/oEp6QhB1bvzmQVyGUrVKr5g
kIPNDS98b35egP8geqo5iobSxhKXMaX7q71GRt8yv8XejTs4mVkILHnAuM2sE5E2
e3d2MoCJDx9JpG9AO7fMGThGunwQwTlyIRMaAqtvwPNEm+pOi6QXFE4izF1KZEYF
JtXa0dIOKizz1sQwpMgB8UFHYxr7DFqd7kDjXDlJgmiaJi8RXSpjBpPibTbMyNJ1
mnR3hjDpFc6NosSCIV4mnjThVvAKPMc4DVzuFtLhgKUvqbFPuquxW4/9RqZf+Gdv
ncH4C74+PEyzNCH57n+bIEUTXwbiYqpYJw+SMbtVyhhBHzSPPy8i/nM65AAMPA0P
VLYHbjfgaPrb4WWMUUrXQyMgBa9Erl0BCMQssvKSrHCLy532L05c/sF+NsSnZmRy
RC8la59zjYxJhwdLBVLXc0UXc0erj/U9ot/wxG0QNja865aWJKO8BBkdfYPFvWJh
UuebbQiRuoidtpO7vJTnRYa3xDLjebrnJZcH4UuxUa1557+1FAbv2bmhSKy+r7L0
T0cGknHdLh6o+YlXtbWONGwSrZ3nHqBoozfaY494ZKOwfpttt+sbr6tNb/9fBKgm
7g3H1JMZrURnV3DNYbLYt2Hbj2Zv+5zcKFqn5fsN7B1y+ZB8p2Wc2uofFPDhrT4f
N99HSuDXzY7Wm5rTlv/dieRWAETuX+FrK5gllayvmag9FLC4F8o29QHLaiE17qU1
mdQndcrUo9F3LjJkh/0R18btS3ECgfEMBwWG/duZLAfHnToRIOGy6O6Eoo82RH5h
EVHJqXhkreBJPsfg60KhQlenFaE0t0EDuJF156ZJvpspm4KaViuyXpWm3H0KZeka
AkChJE27HJgTdhWnAejuhMXcU9IWw7w8qhGlFNSG1PV7VAdpvrriEHeEP+PHUzGh
DsfZ2qnBgTzfVUo31GyO6R1iI+2bx0a4PP6hhACVOvZ1Ykg0wOUHnuPmEFDrDH/Y
9iBEDCFJ5GumilKbIvkWKdACR303Fnw933w1T20FFUKwH7sH59fFkfPTyThKZ9xP
atUN8eNihybO/n7v4yvZP/U/8A6DNHqqn3nxpZimWawYklhtlcZPbNZke1BUVt8x
3LiG147YBAW2m19wmoe6B1tHmOIaIhXlHHrCUSIL6PvZn/9Dp+6KE6MPo6yZX+rg
kmwp3uDLgF4a0IXbBpKBkUnf72m8G31N9tGaPUSg3jwlNmV6lZ0oZiulf2WlRkmI
iTq2TqOawlPOutBtNhF6AYPltrO/1HR/c7MnrQcmQcOpTczjoUzyS16+Vt+SvgSv
8w9vLhSBJDTppM6tNKq2iXvy+UDvPJHZ4hurnBpuJLS/gxHNZ/F0hoJ+1i5M2Flt
Zt3ldWW8fPswsfJt26Asu3nGQhXOkvrldOlRRENivRpiiN3QZEqbdVlXf2EhIQq1
fMfxbi/7FpNv/7jY6fvM1rH28ZZvyU54LQbk+Ubzg3bGx2FU9YI5+tzi3isGZwYC
o8idp+A14rImdR5XEteUmKGp8hyN2z83gwaDIXxvkhtUEFWIjSPVWpaBr2/tWsvW
ggOvbPK3YmrcHeW4AgaPUOJA5hcNLN/CSomKlkgIK9ZTHsw0cvaEiUowps88nZAS
Eowtjv7WNUf9xN5fIxvz7OiFozL5ppPK6dhk8v0rKfNj8KpnsSHwp5CKI2XksVyW
TSttruDVab1TICt8bLfNr5q0u3OPnY9O2V6jlVT4eWhkAsmaSLBEZGXTYApzxu51
UebwFemRuqwmEtRTswq36IbvBl1eH1Pa7qqC8peCLZ1UIyOIBKJXqAlxSlKTE1x4
vmnaPIlcRLq9hrI9H91rnhtDeBeXf0473ee6E3V1pUoP4zF9VfQCyXwSIBr15K1z
9XRt6nrxE8fmTTVz4bBHpaC6KfUawzngtvVyk/DT0n1qLCY5YSUcOiCf+p4pBX1m
3pYXa7Ag44y0cA9+Q6s7JKTPPmDvlXm9mC9rBwG18soqoiy1LqYeYFl9hS7fOcte
Fjzcms7puZBUevZgLbAjzYq9wIkigauM17YtdV5CFcWJD/VqiuvG2qLQ+aDSKhqs
VCy1Vk6MG9VVBJgp4ZTy4YA9OTxwc28tJ3ZstEIk5rLquH+5tczSV1wvnt1Hg06g
35aYO/s13v1cDbvaovIAOTnZ2mGwjMIDKZ8nTmsolG8rrJEo/YqNlxls87zKPMeL
isvHVKhL3X9mFD7sBRgJMbvrdmS2qFsv3BtjjebgWm7BvoLUrxhLJqB9nGn22dWR
lnLrJ31mb2U7P6sGNEUcoC9ISpJwVooG0YSDg/dMG01F3GKC2/1zwZDHz/W7bbLw
mP2rX0cib142zFKrhjdxiHA18Ez/gCWQvk6DLQSiF+ASJ/UINfSNl3Tgt3pGbI6A
rKPtGEkK+h/7LyTtVwlQ5JWkHGaJE7rTCOsQMl3zglDI69Sc2L63Xf6t/AShf/71
UujgM9Ym+2BqD3r9ashJShD5eGYlrEb0MuEmn89DsNSahjFBEQz37/jaPDGFnmWD
ED96sGK35onRG0OM+Hu3COPv2aUM2RP2Bql4yfKjcYZofByJTkYIf/wK1aFqrhI6
dvmDhIQvfyICRipNxbIKR01hxscjVZoY2AG5Y7Dcfey48ugkMZAa3QYTAt5OZwh/
20QgdJcLxxAG9tdmOevhtq16ad/peQyKCbapFudVHYvtOvWpLMRcCRSyvcLm7jMv
5wsh3RxESMj14p+jRF817YVE5vFfqXBsftiVk9P6Enic79+noh4tbUx+dgTWn8RZ
O/CQCjgnZA5Zi8jIbdK/f1zlK/tOA1dWpuLNGghGWc8Z+Ov947SLXxUtqk1L0SMh
JkCSMgZZH6kCf2u+saSXXo31BSJltz1l/ZojbHHImJENZPsZ3MlDT880UFTej6a7
LUFvybt9mpT5b0PPELDBb8V/dVjuGIRqc71139sLLazDxdCGCxP6sh/TY2xOcU/D
GNRTU50NJGIRXkA3oLr9vWGGTC8bWLWspoKFxQS6wBRXUrm8gPZrdf8NVgbsSVQa
ZZEG1+55b1qnnBoJjCjs/SvLEYge0SXDneccclKj1NsfJGRbyttsax1m8BCrqSMP
sOC7ygu+UjGgqNOHlEiYIraT8xTbozSj1SyrxIVYTwuP16N23xnpUy5aHTTA+EMB
FJDBbt0HoeY4R/Q5SFtPuXq8tIgqaUIzyaCmUZnWIhmhszjp8E4KiQ8F+0Z4eTKq
dC+7PnEW5hT2bP3C9XKgK2AKymX7CNJsS9aLSfCw/pVrCcFysygCg6u3OOCe3787
UdaAmRUE+51kEmUSRAppCYYf1JOvuQt1P3eXYV1NJFnDdTtl0/PbEM8n5i9Xvuoa
FryO7s6iS51WoFc3qMej8eJJlycUG4iC7hbi8ByzWM43kt1D8DhQXTY7QeojSKiF
5zGwdzgayouajwXVWZc29w==
`pragma protect end_protected
