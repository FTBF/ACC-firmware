// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 03:56:40 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Nntb9dryEx8ST5D+7oZX2HjIcT0bHi+F46/WfG5ULdjG/i4K4I4yWmxymZhvGyEa
zDe+eElTTihbi/iniNrSt5ExudUwdvm9Z4eq7+3fTHVxZHvqdAl49vHqQ8SA2FOo
HFCcSf5Y+7EDSsa0DdkMAAN48sz5YJnPyzyY9xQkkVo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28208)
uz3OnNSMpbTdsr9uxET0ib6ttvr2j4xYdr3kXVmeUB4ae2EvcaRx9rZBkyKimZiZ
BPG4gIzfYDajqkSQdfi0d2s75U0c7BVj+wpaYeQIQXpF7F0CHRORI+sf0ry1oH9r
GOly3N4uDddKgvpT+dmVTzqbN925dqYeyTuzp7m4VUwehC21EaFKFE3RXSMGPMQc
FG5uD4AkZ9aCJMpNjpw9XhIZGHhtGDp//qK1qbm800VcAJqPJpfCw0qZY6jZnMUD
PqRFYWsAbHFp9o6uQT214vu7LaKwN9kbDGlYDDy3moCPN7pdJMw0Ao3L2l7tBZel
hUTJxKg9NoW714JvzPj0syAqNPeQxxUiENTBrvmy8Jldk69JA6nzG8V7DWLdnJgi
X6M/nJOLcQ7twWIkF7L9M7cnxrb7QqYXhOidduSowHW7sX2KYXFUiCFGIxW0GIZ1
kAV3bnp+hwc44oP/t1pKYPBUrft7hwVg/VMwajIkfIPzayJHT/e3MblNhvhFdPuE
i/etFgx5JXYg40FfVTo4ssiRQFaRAcduKIwyWTqDM/3kiAVCCe8Dp+RGz5yAXJJL
IrmZCKxn6JiUCbmMKTP9BO+jstkYqE3VSK2JQ6pSDjV6TjOUXdmLXa9o1CTCic7y
NaepXSvV4KJPBWXvQI2XPgfP9BfAAZm5Kts+/FUjJIhi4XuBVKwTNGq23TEGP2vh
+PinVeyfmFcrVwYWgI1sMVzo8QDfoFIwphra31ST4pxt+EpwR1mQNQJlj/osKc/x
uyHHv75laBbKIlVKdVMcIEvKQV34jLoM3HjLGolz9VDkPBQPCvbZ49WO+V8APPfI
c0Mov1GHJPsf+s9TbeON9jZBPP5vCOmmLXwodvTMJZp9Ph7HQlJNsA/BIM9xdPdC
6Q4QWurP/17g5OfWhNMmpZB41mmzFQ4JKZ0CuMGfw0NqMHYlyqex+8EO0rmCpVEn
RM30IBM75SaCRXM6VIZJ1ONGsh2xjTn7uR/GxtKj1a5nj/2LgCD+zxK4TqNlKTmP
bsDC0p+/r8ecUv4UxLmkrPPTddbgBEQI59JIap5ZqXWACTYnuQSf9zSxG9AjBak2
WPCQHAHQS5C7OQXpJ1V1CBprOybkGL0N1ZSfTCnrabN6sy1j7VmfKWhDiBeOt0/V
Ymkj6kdZZhWQVkfSvOKu99+sRMgbP5Wh35uatGh6VqJqfRhUafnREC9GzdT7btwy
bxpURPQJk07lOvber19Qc97sZCdqp30zyyfDZToqjuUB0zeTC+aJgpWdDwfzj7K2
BsMUh2irY7o9I5UpThQSFtb31yQ42yJs2us2vA+hvdenbE9MEUeURWaS3hqbj2Ae
OWRmlOctw13Qi89VzbcpHqBAlYS9wVls0ZEdqVWD4tnay5qpfCnePfwlE7Di7GhH
aiKmD+eb6lCOzrs8w44huLfutboWP6qjznPchxtLWwTpgGvxT68EmL83u66/rUEC
HDC6IZFT6wcs51CeeddpxbbMVVrie58TJLPf4dTTG831n0FY5bn2JpK9LLE5+Cqp
75JnRgktT+Qd3tvjxamjBEgWVkHkBUJyxBlobL9nFeZnN4Gzt9OgFqhjIM5s5U3q
Uhe099phPygaQxGP+Iqr/zsvGAn9EnDO26A++YJMEcwX8y6dSVsOYdmT0JYQFD0q
9vuzJAWKBCysoTZYlMSu1e8F3khBTHceXLEA4dNR56/VvzYLkncFvch1xwY+cKNk
iICqUBZVVTG1DTHTWUdpexfuK5R8N5hDyiGFcA6zUfQV/UMhtVHZQ0qxRLWgAzko
Faxo5NoLIIrCN4bbTv8rpquq0u6DXBYZbyZN3flr0K4+w1lcyC0p7AQk0p7KtOIf
lhs1ofH3bp2M9/KmU6I+8YvkWe91cV7IX2Vjm9hfMmx8UOyZt0+TLZ4Qmdk/GLGH
1//7tg75qSF2R9beKQNVZpGBaKFpkdTbgS6lr9mFwulGx4kJbJpgj5s2XD+dFB1T
ToKcZLn3GnF3iRLHChx1ztUDshj9NMnLuYO8K+vKDoAbEgOa5r+f8CZzDWXBc1EY
bCRRcSCFtYNes4S9zbOqqTeCBBTDsEQ2X6VQytO0wX9Bnta/Udjdx18h/mu4uXAm
KmnCmdlI4/bGhKiRgdFFDWCwr6G+x+hJVeoK0Xmt/yU3yhMtTUeT78WD95ZjZ1td
xqF631mwFxNcPeKbMdGNL6rkC0drUTj5/V+Ld3edauNcYNkkkljZ9rh8ZxLWhvem
MFE+IcGIqfSYFkjzjty9s1hwJiX8BnFgCts/OFVNizWRMbLtKy0fhgK9TVxOIa5h
k6vCPICQMYLDnZP8iT+tCtQWb3ZSTk7pe0rg6TVL/5HX80AarX8hE5higpIGaJHK
BfXM1o/tqTVJ64SIS+M6JdJjYEY329hgOWH0nm8I+76eoYDE9vLxIiqFW9zs3E/2
e/cKDSygvrWczz4eeq1dYuZE8fYjtstWefhkjOHj2SKZGsRAJJPw6VCjigA4BXf2
FkdR2rNPL9BJIBPdzLrExVbPRDL9JjtrJAXxuRcHYMzs+spby/0x4FQvGIJxCpIy
aXUPSiWTjZXhGpFkxeMy35E9phEu6zUm3Th2PXDJmf+RDdM5zhWGFSjbg3IFzZg7
rQ/TMKKqyOloRV4UeNNUrCisvq0/GHg+3cnvTsnntWxH+zI5eXfr3ZJ3wgZUCRMJ
6vGNzi0znxwtWAZkCAtCm8ZldLLbaq0jRNcYA+qZEkF8ipGX+8ZrJnHKfr4jqJrK
gb5ctR8J2LfgHhj1kIg6rFQQqjy7jV1zItF66KLDL8LkRHJjONjRl+6/6yI3eUz4
Wo7uAHa7DHmILmNBArTedZQxo2BV47LwBKOMFslMV70GQw88ALCeI6YYbBuiXG5s
hcpzOoUs9izdFNopYn8jtDJHPnceH+k5CymjqSZN0S9IYZvLgX5YJLF8OHJWpMS/
D18IZt5Q6Rk2zw6T4u5xQ/j41X/SmLoV8qsHpZ3eGNqr3mdApUDL237P+6DyOO7T
CakH8RV08XU+aeOWas5OzsfCAshUW8vcWwYdNoVAKrfSkOzMTd3XzLbk8t3HthWQ
9cM26eaOirRh2TMcyDAtJQxo5rUgGCZtgraKOd9CEDWWpEw2xp/gn9N6+0Kj/U/G
KoiftwiFo8ShE3jS66VjGStOXkxEBQjQyzARFqUDYL0nYpC/+qj+IPk1lks5Pc4t
R1wZ+iWw7w3zlC1/Aufte3t3Ym1+xu20QpgeEQlxJbSp/UY7L0vtGLAjeB6z4QRc
iswqtQEyhwcIfU+989l41HrShIUoeVJPxLkoOFmbL4KlX+HMJERSQ+xJVlXLBrKg
Hfn/kVpRoB1pt+9lkJfyUf9PXEOjoBsMg9pAEvsy0xQpZrWr0iFa9zAfUK/iCkEv
JrFf2L4EHMjSfeRm+eqULx7F5YFi7v6aelvM6cRbn+ZPAWag+y8m1JGmnVJDWUwt
UnKgUuaZNzyGrXCKmbpb2W8QHaxkKILeFvBO5uANlWDf7qPtveDI19VnRgVCYXSJ
+5bXFkR2EB45tc/ut09O8nfiMKTuNEmrq8FtbTvbWhgb1dO5VbyPaClCqq78v1eZ
g7+ofuqbuO39mHUEdkd8uYYp4AjKire1loE1kZAcM5GV3/vXRHZv7A3zwOtEKktE
I/Yg6TM06Yuj/oV0edGd26JbA74QHoA/l9g+JMM4mo2KNtEx2xlSxuDXLx1FdRAX
IyE2j1lxFe7iHZ1ix0NyYaYa5Q6j663ePr3+9Lyt0qjg7QCLTqcCnV/OXOU7DLjy
JxdTLfkX6vwDTU+jT39xk4vMmOXSOPBc58PDUnnuPTrT/C6eTllkLaIEecxP8bs+
0UkgBM0oBrwghXBk1v/qs+rJO63UPogeH5Yt1yg5LwJbVj/Cjna5A7vra+9khzoY
0QjFR1zaO4DeS9llnDJxoiSSmaYnJNOmGsAoUYWBmh57eUGuooTYZiewqzfissc7
4BBg3QMe10qhLxKkt6zY0lrXW8xZTTlwa5xiMXIMH9B80vCBCqzplf+SVqptLW+2
p6HmuRpalmZzpUpQ0/UYGRsDEOk+7R2XJDqGuTZJvkak7UBAX5FeUM3I8Ye83SV5
ghhzt56Jakn8eeXDByWhHnV7RUAhO7cgkcaOgJPtCGMZDm5gdANRV3sO3+IcEdSv
tG12JL9I05hBZWpj1ZtTAPFUWgXoTkCIELwjI+p1Yp0zXj8+8tuWAaePdQy7ZR58
76gVqgbWppgsT5/iqFedPSdQBJEz+WUJRV1oHprcrbiTLHjoWa0r44sbvdY3l8BU
sCcy0+N82jeLT3QvTl0XWvzqbr3n2MXvPtVJdQCHCVMa4tr6asIuDThHXNdZ9WPD
vluTWW4TfTQdXKYJzvklc1sVnYpLmyquUrQ7G+oG/cdbknOi6E/ngRH27P44J8U/
DhxImnPjLjgwIHW1fWcGzgr9HMsSJ8onOTKKvqaj94uBDZnIR0lYehR6crx9ITvV
QNn3vcO0WSMItd0eeIBS07ycNjR365PTGA6otu3vBKOiveErxYkK9Ff6dFiEr4Lc
b01f/drdnOBCXaJSd7nr4xAe0GlGJIucW1Ly4B7KrtEYAVyl16yuI7TCtXMeThuv
DBYPWHcT2voPPpribWNKkskdDVN812fbmhOBe/bfpwwwiubPZe4YbNPB6U3H7sDf
94ESYCiBDXYi2tM7AB0Kn98GSQAqNGUkCRaJp4UrggUkFXmiD0VtSsP+Y9TFRo+y
7xVCbEKll1RhWDBSigNJJV2wSoiEHkRsb5cZqnoEwGhuZDUWe+hh2FP2t3TQGZqW
/362OVXfhAhfa0x+evbapEUQR/Wg867lVsDopw9sZQfeZ6z+h5PgGilsKDGn2bbs
gtnQ7ntjGoTWVR6pp8Hy9Po2wTBkxvN+GAIvR5kSzHWyYjtuvnpTPLut8ibfu0Zx
fVBvC9vP+G2B3ftBNBXH34K3cgfCHA7PVX9iBP3Jr/3IMVxugwS1Qv+3ZVYCM90T
SdjigZCaIe7RJ9sgrxYgqlzGaLDShDGHkvxr925MMlH8NcA8BoNUAD5mITy15cC5
Sdm6+5tLgit4fkC9qPPSwuPWVbVmT6NKLVnZwJsjZ+M1IJxVOG1lbMfPUUB2sEUE
SMi2dzukZPMUAs9JdiP2qDM/VPKJTMzweWGYjYd/FlWzk9PXKd06Rvg/NavgPae4
+IIV3qKOq2iiiSezLls2Pz5EfehTACr9/VVBa0AwOrSPYeDmQ+ksH8vZj4YZE8+b
YOVpoIhB0VnNuM47GT1oX2Ja0m757kQSFEi++3Wu0hdN2PWHbpXT5VzjkJafceDG
okgU21FLGSZDdqBLlQxNBzNq+oaxLTLRWx74RXn++htxmNxb/mHtjBXOYYo1TmKx
dcJQq2VZeEpPmwcP3rV4hsF44lMQIQj0r/TPWL+1sLTLGZCISpxIrqsvvjqioF8o
uCN/OVAuQuchbdHb1hrLrfvDHLPCNDI0vcTA40YjX0CR3kQjMfO3ASx3O6eAJQD1
bVQJONP7bADUevQtcC3XQ2ns5U1/NsgyxYPkWxnhXf/SDopyx3vabHPlqU44U0Ag
smmjK0Rf09II+JOhIxNVFC0VR5SxKWI9F20yw3KVmo51gI5JmpQkpuBMrHkCjGe2
VvI10pfk5A/TOHXvzlWMXIFUxECKGvn2cutBs+4t9TXERIcW6cK2bE8s4m7SavRF
y3ytBF9oMhyxmuiu3iAZlp+FONXrRjwZwQ60NwyBSmgJDxbf4d+/Fjx9eK6lht3M
F3Kf1LMmdmNUO4BLZ3hrBvDFOSiaiMhOjT8M2KovmHEOo8J82GdFOZmt31xEgaZW
Dq3/uN4pFhS/Zq3Nd6L+Tm4PnGBCvAgu5yxEndtnJw+uaShfHrEAEWdcGR2/Py4y
hk2dYHCqiGPAU4lRj3a52lFHxX0PamBkJfKU2g1LWyPmHuiQFW+SKb2ybWMxkXma
4di78id/UQ4QZ4IC0iyLoTrrhLaD3Y20HG6zJpIPHP+WVVICjdC9xIyDSe589yNL
6rKbL5FCYO46JaDmV7eRuhGmb8DKSZBvuFn5OHtojplGK6Aa3IWtNfMLbaQgfaBU
9J2B68+ZkHtnkMBOU3273kBDEW66mKNjBHBbww5Vphx4UFkABKUH1CUNDLtwY8is
NOQpANQC9qCHObVtEuJJDR6z427DtViTGCHyV1wxOE1q5cmKywcn+JchGyA+UEcY
7tFSZ/tzB+7WCMoNJVGetNoWDpsWDGNVPriNOMkgeMKzAzsxnjLVxXv2Ns5GC2MM
X+4Aq7wO8XAkxruyS2V+63SUlg3eHIoXAqRbHXv6KGltNVD5NTbdOPg9wO+glpnR
eq3TLoi1eTqgj5+DpIMMNSuDf1+HgAbiWC/I61VZy5wg6F+52AbCoSxoLsMbR0Fz
q2ZgAHUTdCK7dely7jDH+OfuOykDtB9y1lh0sd/SuUDMf0Run+1STosNxw3YP3uM
ItYoYt9N5k4aqtfeKLMS1hz87vIJqAtL0LGeuTxJ3UJ/GCZHQpSuxO4G3GtT2qOP
VzIor2ueqMCKJMwGuvpRAjIHcj/r24sVhlylK3yYob4sfB7aSVZwR3vj/qlWRzMt
moDP8/1rOy5Gaqk6VszVlaNLi/UFyEw5KczFbYbBcnQA3PYCZGzvgdQbg1HdyUKJ
H+YhWbCZKCZzZ3cOlkULhWltk5WADpSwB1CbiSk/ZaPPEfe8flCxScCr1NtrksYt
TBqTtofTyE8vcAfatws7Au7OqUO5VBz6xbaaZpnH6sZuAH8nwiWDX5rzblxklduO
6KFyr2f6n7jx8h/ebCa+GuC9x/GWzCneOqzCSJVUh5sNquFcQK9Jep7iV7dDGIq3
KOJuS7wJKds1qa4A3zOlj/Kq0r63vnz1etAW8WhovPFL2HK5awGkjKKF5rn568xn
U4SvMMFExly0YiH8Emq8qu4gYzWZHJURRB12ATtHyEWU4Ao2+XZOvkwW8Wjv8vi5
ZqjdVLOk1bz7DOxpRPBvY708LgrDHdoyQgkWAzykCyjRRrK6UkemaKGOP26BAR9z
EbZg3zIXD3vTrt13Gqz+2v1nitNPkoALUWfLYt2TaIZtlpWHDety0H8+mmoY7OVp
qh3XLu94QPp6OnpxC1XfVbdFKp9hpIyvWomCBplZaz005noADqo24olpT3bkDIdc
P+pbx46Rk4Z0jGs3H5tHv0C5xIS2VfiqLZldu7O5TbXZA08wU5/uNbw03TpQb86/
eSeTQxSUnEFWt/lLmEEmvi6kQC4jLigwyQzjYwaVVWXmnU5xFbg+68zbAhcDgFnP
T2N3eENKq4+N8Vv6QevI1IK6uIt4SI+FvnqxljrWiCwQvBjJCVGeebeHeXXt9d9f
yl7yE3pAPjQryMkFzeLBjzOzcAOOWfH2lDdRkXCutu4enu4jM16MMpLLEkms1iOe
MiM3FpIdmp4s3suS6Z3slj4E7JIe7AUKp89/d1q/15eV9z3o0sJMUQYr4EPNiH5+
xD3hGSKhQbRFAJklZrq2RYsVqFC/F7axclJroSgeezI6/AbYCxP9ZvnLt80pjaVe
+q9q5jMWqT3mQn92oUe1ieRE3/PFThHZNH4jwuHUFKXkMmU4NG6wabZJuCOdI3cD
LgGHLmDPQ2aUqvo1vMP5Vz4XelF+DSDzI/z7pp3vZYISiPJ0IBVU2U5kZdLXbZ/p
eB9+Z8TabuTcJ3ZUVaxeuxTmdw8nyBSuBR6PpHKZ465ICeOL/z9+d24TfXAcIDbv
Y94uFNCnHlPp82pcnG0pL3ysj0OlQnkfg6eZ3ZJgMFpsl0t+3WCfulE7+jeE1W6k
7tJ/82wWoXdmR+ka2jj7vixNccuEmTHBgNeyLK0Pi4/DcvLquXUXfeaVG5nK+9pl
9exX0ET/nB6CLbJjSSO3Y31Z3Eeix2XCIluf+vBAtOzo3UJRk6BEgIeD5c64qS+f
IofdJLi33YEOF53b/b9ukyq/Btha9Hma8AXvwkSH504suVO4haPpwXQYQtIAV9an
nXJ8pT9HcSh5MX7taHni13zFNZ5mxTv8aSd9g0v72+Z27z3wevX7wSj8z0X3okTn
6Y4c5vs00GdJsFBpH+ObEeu0khqjkXribrFKYaCKwyzr2WAOmVTU/jMB5B8wSyXr
FWUC+vIzxMHDbPOuc0R5kya3wcwDXJgLgIKom4ir0x1Wn9iQNUNy5Od0N7V0r/OM
67NcRpfqR/XqECjny3Mv50NctPVYoV4i3Q9ejyedFrKQ37EdWNiA6XNEhQYtIpYn
DP3DGPaQCBz9CC9YT4y8j/YewWdRsb/4Hc8YpLczPNYY3LgY0K5GpC/2aLiWLH9g
DyNGAYhVeA18+sqo86UEIcjtPEbi5ORZJDO/NUjtedO+0WKwPAiidoRF0YKXalZ1
DaBiPIDBtuYunu0ie4LDU7jUEdTHn4mDefvZ0EdfSfgBOgqk86cjd711hibAGCD5
ntnAoGzNT/3OZjgVK1Uc+z58Nc98feXDLYTbW4g0Dca56amuV1I/r5v5g80OQ2Ur
Tn2x0iWD/iNJJV6oBmhxLQn2k+/AHHawG0X7g06xztCJuSuKFA7LsMJBHiHMOmi5
FiOuu4jSg8ypuS63NMciyPGG7Cn93KMYKgAqivpkvMmGIZltl6f0qvY5fvo1Tb5T
LWoHJVPWdIMwiTB3NmSH/2+9gRFQSOMfL1ypVN9vaSfwnGOgxn/kEaLatp19VLud
ad8XaA6Vh8Q1tllmvafs3o+aEV9n0L33eCoSikndGDNQoUdJzoE63yKVvVLQAcC3
WD7NQi/0Tmj6OX4NQ4GqtR1c6yEzBJTU90pumqH5HXh+Olz5si8cF7a8yx00OVt2
msP2S3c5AxOLcsIXoaDwulPOhnplB3RUL3Vw/zLEZyn0bt/tbgiUIsIfaXnH4eSH
vzhcgniRCIzploH+CprVRXSCIy/hTCRScv5njiIpjXoJUEDqdxC3h8Yy6Iz27Nn0
lz+dojQDkat9u+ywVs7K36JeJnMWebtHfLmlgDwnLnxN3E3MCWCqwHEPJWRRHMZI
5DFJP4wBABVHYM5NWKb534wwHYjPQyLoI+5gj+qSAQKurHI4EhWIf8z2PvBmb3bk
hSBRsVD9gFOte7v3V/17nRNJA0UgFCEcz+siggSuGfbprWILKS6oSjhJJfOoyUd2
/VKvjuaaKjntX64hSMRhn8kaXMmbbLY2fSvPx7sEnTRNDnBuqeDSRhzsZy9Zly6h
2rMACgz4jJSgCcc19bmr0nobpSaJRn82pZwzy2SC2g8RMoZy5TgVQLlAJd1YAICq
jSO8UEcJKt2zev13TIQPc2sICShXAfDQ1O6yr1ElUPCXLP4MUXti9txL0oxlhjpr
ERCxuS06zm8H7wn83oM+fwU7mvzyP85oy4Wi3vkpgo4tyqVdlmObW700NSI5GbCd
HvdKZGQjpBWChbyYULe/PhPz3HYa709IS3fhLuh66Rrr1T6SZAMy2DWLJlyeJnD5
AZ5CYOgkIPTKIEzp5Vj3Qk596YicgyUWkmcjF2s4isAtcpYtienrssTrHN/6rLKd
ZguWtvpRWYL7KxQdis3/sN29KBd6MP+h3nGHuLUBGGwmJ8tHigKkCIrWC5i51lpB
L9kO7zPqRp8cbq32znBoXzJ2UIibaodC2afLqr5QIYmnhkEMzaTkdep8n/KmatMK
DXzdtC19ryi7OwPV5NMhYY7F6rlMAto/zYtsnQHAq1ReRmEC4M74rFMV800+jm6f
nzrPt5xtx3tnZjDLTXqhGEmwnIMkGwQNN7gRzsLOnREDvlRxXyN1E9U8Fyk/wiHG
cZo10IC66jCVhQgnyJRQrts4V6caAt9kN18DedAT+p9qF+fmM6qXQvEw4UUgDaXC
cr9IxlQ3YiwfnyxJHN2ArHFUQyIpBlvfvKesD/rZRTZ4vaRqivlBD3RLOlCmvRGi
mFRZcfocwN8DSB+/MrukS9YZnWXmgQUe5bapUwBz06ZC+gaSdXEuDVPkaszEsUnT
xoNuiSCIkS0iu18wBiEWYA+nGT2QLSfcft8h+bVxa4FI6ULUWRQPePNCcLgCKl+r
xj5ZkFnDkcrsW+PUPZ7TKHoK+3utFcUXYKJqtfxtQz0ON5EYuzviLrOyV+zX0yE4
nF5V1Zd+KO2AYTJR1xDV534uLwTtJf61WmOfTKeZjZbLMeQyOCj/iCScuvcXryar
XK3I4UWvNxljLzJ7wnZgeZD0HLfBnnoUDYlvSu9hjXPaUZ8nyu5TEp+ud3osACqf
y3J+9V44d7tliPHlVrKsEftMudJCSyrkopSXeRP+Q+nzerOLKkY5kUkAL7d2Mn8H
3WnKTFGc+IFQ2is6m3BjSN3wN2fUTSVlRHs4gmiqha6dLh9Xbwg08Ax7707Ekh7A
hiufHMp4C4lYnfE/PMKZjn3HvOuRK1L1GrrK4E4icbxnxKqP8+Jy7PkegC85LPdy
gi5vYt4507rC8JI1NZCTpGFqX8VImPtCSX0kY6AFhrbstd2yGqZbDxErhbArPx8j
vfIrZtKsqk3ivFlfvLs+r3mOpCW+aHDZ09Yv0R2MzTmvoSahJybyxMq+30LA7QsV
Ivrurh78DirDIRNWc/d86jG0lHerfyz/ExHji90tsqY3I9orfYGPUaAeT8RSR2bw
llYbACwMr7U+D1c/H/9GbpQTCJ1AZJmyyWEEJtCSFnadPrjf0VN2OjKBOS5Cmfyp
gkFDcirKoIxWdYeAue5gsGA/MSbrOuPpOUunIaCKXohrC+35b900K1puejBi45S+
EPEChUd5z1vVQUbZ1Ee3qJy4dQKM+HvtR0fTjB0inu6z7AmXmcBEQbBA/t+70Pip
bJZ9DARlfyJkHrLHkK7mU+3aPu3CSqmIgnYWyJhK2IxqZtMYzbSr05YkkgRhWSx6
ejulk/FK5pyRH2FYM6fb/VaIZulhmFgr26dJUAjnAOlAnnoWrJAV9lR4ZNdpBiFh
9VyEQ66k0CAUB3YYVFBJ96UMN2WxzcA9lAD7ox6OyDjFjK2mk1G9Ny/k+vQpTH2Z
EAYpCTfpugQFXFz6F0/RMPJVqdlFO83Sb+GPeq1ewwKtqV7UBccRqoxuyOAHOGy/
6hDxsIJRc2OxS8BK6tGz51jJN39acVQM2u4Trz7Yj3Bmy4qu5Tvk6Szg1IxPfAES
e1VecQdwOFdYpQZPO3jTtd+QsmFXPl+huomTq8oUSF5NxN/M97qQNkhyC5nkOem1
9Bl1hanmoA/DdVq3CVolBa9L6N8hbNFKvzeR5w2YRLOyVLbbFbK2OU0uxv4Fwr6s
ftXzfk/+PnMvx4GjdCS3npSYaVc+nqzC2420gjU/Gauj1AlIDPmO70GlvxSeQHat
9GU4ZT5NTxPtgUo7CHA7KaGkz+9ee0FsEB35xduKhFbNL2IL5tEiJjwlp3/con0P
aMVCGlC+7DIuHVa2YTHaHxxP4F4Stfdug867hl/JRdZUYqgGab0v+9y+nlGR2KAd
WrWR0p2XVslc1uI9FOdsdJYx5F4psjB0hsjYqHD1jfgDIsXmQiS6gk4lR1nbiRme
zekm1yU625hHeIVE1QvmzWTC2lIQc0A1XrN/vQ0GpK6RzZJZbWGYYHqXKYxvogv9
hkLGIWhwiudkUATGTpCaM2aiDJfKJx3q45UeuwJDEAJntdKKb8pd0fvBPsr0OGq3
+FwxZ+5d2i9y8AZ/9MXoxIOOSEOaYyCzad009Om03ME1vMr1t0ebkqM17B+Q7xrS
lPBdNN3qMCkvDwDeN4xajdUXRGE7SigNDZ+M9l6kJ+0eVZd6IxY9009LBtNZcxWe
nz+MqQEE3/sfwQHtsSST8jNsAmKBUwQ8jMKk4CdQc6P1l7Gwifn4uLiGLXyV7ump
VC91phTIw0GGEmCi6+F7dyBWcncAKbBLg4F9tlgxPH+XFJ6rcUA1e/qdyPavIswk
DLVE+Ng04BAcsXtP6Yl7lmXtqtW2ngy9hKNE7fkQKlbZzLqkkiv3wiY0+hwUMQhT
sODIan+LHt+gkCAsKWwxwuf7A6EAVr1yBB9dBssaDrKd6fKMSLtDioX0hvf1FtsN
YZ1cock9+JG2A2TLKr7zxwhrlJ67wgHxE+b/oQlWkDm73sB2ijbPsjvePiy7bL3X
k+PWAyMciEwrvvAy5rTli2KdvRHWbxmueCn9AEd2WGbnnec7rlI4O7hPnhwZ5DSH
wlA7+bJaCu9UdPTzg1A78UKKbfQ3VMGMJeuTnGILR3swPvZAXSFR3zG1yLSCAGwO
MfpZikfsK0feuwOGiYOzwFG/R2bfbUFeYAygVLSzmQR/cLDYENEMCJNXx5x4LERC
e3wnR7e0enJB5nTk0VDMsDDwKH8PZOAssgb/Db4DiB+Y77NT8quR1dSF6QgcC6KJ
YsU+j2KLAhUzZbVcRTDeqPh7Y9cENXHXg3LeiVvsBAEaYDTIhYkP7TWqaC4SdYA7
6+6t9Aaz1Rxb2NqOylyrQbr8kZDfvK/1AhiK5+wtxjSvCyeEdYzUglNdtEcqUsB2
K3abpx0msTgGCQt5ypoC3qemotEwqEgT0/fnGmmrcWIB0TG9BG5D68b1Y/50KMV4
bClQTO0/0fS4gmsRbHgQdZ+ZDZWjogl3Oud0gPEVI3VwLVgQhnqSz71FNUBN6Yah
cboWDs6YxOov5fJ8sth5pQwNwK34dYNYSva6vSMEgI7IB0Zn2v82BdgkqYKWJ9Xa
5BWbmiF5GLK7rZFNs6rpcP8KnscbwpVgAuX2xkelQTL8NVZHvkV5zht+HlIZwVBH
EIy1Zpg2FZJc7XX7+K7lTbCxqEVWFDkLB0mQ/ZfmJtM3axMJ8f2gHE0GGq9B1vjj
LcbK7wVlKVjdbedGiKJsV4f525slwkAjv/DD7b5KbzHhoEyv8yCor4Ve3dAzx0MV
MEoRp2U4jiVa5A2zI5apCiNR+y62HaGZB/BFBF7ieWjlB3YHCJaVeAP4NAEqNnu4
nvKfHJfT2/8I63ItuwNEXn2Wov8iFUmYPefy1aLMNPnnaTrud0ghL4vuFHw9x4fz
tkt6AmCVM86UuqGA3zpocSil6CU5heInVNDWhabMIraSgB2It5nRILlR3uOP5i/X
uZqeht4Rw2KuPoA4AQN3a81rxhrN3RROC8NkyEkxOL+iCeDckVOM3P8vgh/MNuU0
Hi1XvrV/NwXmD0+T6jxXLY7HuFnq4AP8jGuFy+K1zmae/emdaV3TgXy7hUp3xbJx
vnLooCvg69uqgLcInGSoT4SgEm17J0F7PU9KOqwgqL36ts1rUzkWenmIQtpxRwhb
Xt7Q8WfcZrNQ86AuBJuQRbsSurBmx+WYAhkdgSuK5NWtqEnfH4TSAN8hdzXxdQsa
WyyzwLOiSAHailHoWATZvZ1XEoNgVpn/NIcQ6CA95IjbpXlN5Czjuz52/ap3miR5
32Os9mVeMFuQ9P97EXWegfzt9X6KtFxmcSh/rlYY4hYQavsBgyhVroPRl6zFd7Hm
gJuSfjgPZSol6t3e17XwRLYF7mqFB4bTf63NJbHt37KaMRgBaPLEBaDN2Vgq4vq3
MKI6lhSLmF0CAv1bMJEGdlWqYkBXMBSdOGPJyu8JnKcj5kU+It6ABgcOpN0zywlM
iAizlaKUI8wl8tNTtfJIGtrxcQOpNP2tUMOVWLzi60Qs/9k+URQDYr/v9xHkSY4/
1IzcYLw8xeC4WwBI2spEHgayRJm+bStCK705N165e8/PZE4W8YOld4cc2MtyIz1H
dNLezkAeDdR2kJgRalZhqRWZ7qzN6Dy6AuxRxqTmfpl2eegt018xqUiQG8Euee8H
s4HUfN6IH9EfUOqhmcGvW53mpqXfQeWbPJYAw0tUHEKDFGT1jmwNiUdKOIquFbui
ymAN1nyCVma34x1cclALIxOAGuPtBvtUSF+eSYFKKrgW9XTyGj55nWTjbi6BVLef
682rBL6+GLgSdcsTcAYL8CH1uHf7huqKow4B0xD+GS/S1fs152+HWCiIQniXja6j
E1DKFMpieCHZh1HvS/PDT+D7wKuSzm7d1bimNOqkkSrnMv4XlOyooH98jiMfTHGz
v70n/+rIH/H5yODC4UPFt0t39CZQiHn07YtKHW2GhyVORyv9svg4n2XwTYu3avOy
5afE+NfP4V+lmp56JeBTamVWuow509NHSw8lSJ+9pMSnqVWdmq6IZz+GRMRSEhGC
90CIsvbzGY5twwfZbv66YmTQxuqs5yarjH/yfBJ3i/co/QHDpzrMqHw75xyHWQk3
bLaWNs20Z0mD0fLqhH/xJXs0xIlzAkICfBBGhkkHX6lMTida8j7njsWO9re9M6fV
16JKGmgKk13r2xjzecdl5lMe7xuLLgg5YyKdcl9BxzgaocXLG4R5QsEgCJHHf7ym
1HG8m+Bv9/YI53+WKcza0BS9mkByPoW3m/ofsUqvodbw6nnbPUTAhag1SbAQN+NY
xY7fQ9UHQVk5w6m64rXzwuv7CxXF5DAYuItrfIv5k+DzUP0h2HOUlsEQsObnaz04
Or576qoQF+i6OqbCLuiNzeDS2PR2dw9K+MVS1OTYFpndsUSdJDZ4FoJzkCHHDQis
11/WQcsHNt+hWB2qasrPdDRuFhuwJmbUpW3Plj54b8wKqOtpvJ7mPT3huTDfesQ5
rB9sgm3+vdpjToYJNanAco+Qo4j/pq0Ys00AoWQQ5riua6YPwuyZah9VnNyK+dmP
K7JykugAQO3+PwWzAmC4ULh1L4IVOfGAnYS7ZJgQeAkvr3wNLxTze/xw7PUryvM5
xVUBXUbd/pTRIGmCj75XoOob+wf92TTPiqBKo8ctpUMQp4ppKiBNKv9MrWkh+z6U
/bUIamjnUxdg++9mUM05rKxnPlj3LqPWwGJ2YF2o9ScFSaGFW+kNU3mu0vcsvVFb
4DkpdtU7H/bVKhVCCANt9I7ofM/KP+ue8fcRv99e5oiq/kE07aORjuGCLWU0P4Gl
NfAXcUcPSj/vqsXs7gepYpHp1wUalCUMHdba74CLjvauKRb2HdJkwTs4zs5x91ak
G7pDP+HbwpEpsNyvXVZxpZdJQSt/1saM02DLkGLRCyhkU+pXCDUsX6ZhukEhvTBw
oLPMAc71PJFWPTPlXpq5WKUZVOgaO4fEQHRQm2kpbAQzEJf04D5IRyxU3I6PMK+b
bUR3lB4bmNXsvVXwx5hjNopPuxoy4HWsdePwxLcFFbEIzk9x1XAvc0UZ9NfhRwPT
vh0GE9rbBS87fipa62j3apJd+B5v/ZCsDMNtml0IfARnxE1bKOPmS917DYaQCO/R
4CMk1c5zaNALyqRtgpT+Pftshy7Xxy7/fHkVuTv4asv3YEDh5PQsdAw+QPSiU3Dj
A8QdYY1e9F1SEd85PJdTB7lD/YfKcWU64sBRXDyMMZFGgEC5KQznscDtbvh9Mnby
aVsYyo9zO8NO/dqcGuoaTl/fbo8s53qH5D6dzsJIYiv4mjd7b+gSEPxwYd4tfIdm
5S4rJi3PHddEqMoQl0dUdfV0afo2bBdnAi8d8EY4cKMkP4+NDIjEcrgmy5kUXZwD
i+O+QaBzzZGryfIFGJSD2ZXrOu5znq0zPq+0YYIQlH99KjW9POPcti34G7uCrynN
n5I5kUQ0G6HnBL1S1XP4YxiqFSPjKmSB+6tim1ql8y5TZ31Gwz+zUravFcoGCcmr
IWj67RuUB+3NDk6iwVfM2YQydMuQodkHq30ogmOmx16HnklcZgjWulkR67fdE4bc
tLpgk/L3W3lsa1Gq1zXcyEptA1KElQszaEuTdf9AClT9kIpcXMrW/u8vBVz2Srl0
UXDI6pg26Lo3x0iq/2nBXw/8jCW31pH3qvjNwz5YokHTJwSwMWT/pjpj9v3FKoRM
qlCJ39CQkKajV748EOZyiltMlLicw3vMowYGD36AxrvzFMVQU7iX8/0349nqRXMh
YqqpEOSt563zgq52CKGFlhHzBVs9ZZdiL/ZYiAMWrorZKR4VDsLEbWQ0xGGse3bx
6G9wXhHa3fCxYX4Vv567pgl6tMp9enNfQwY9KT5XNOgXiXV4D7E5K7TwtxhtVGov
hkF0svR5iCKcVRWGGmz4i74Yf76QRd+rJa4/YcwMWj0POVIx43ZD8V+F1oP+BT56
DlfUQbSYZMvgtWIsBVzBt1LPWUAdboQUZaPaEp9V5sQGOC+ZOt1QcSGhZOfrrlpi
3cjBVewC9/FuQWoGSAhWvykoF1tMMSCn5RvLczfsaVBm0IUN+DxtkGRDpZTNtJJD
2HVQMUHefyIvuAhpTYe5fNMMaooZPshyKCWfiLEc9nm9rDyNjOXjG/9zPDb+4zkd
UKS5Y8vt2k/i9Qd8xZ3MtJaNi5cZ6Cv84EbaJlnyh1meMUITsl8QJaHVlKU6+A04
Q4A9NXfzGAHgDero+Tr4Pkpb9b6M++IHhFpW6G0WDoVnCU/DDS+CGVyduR1C5zpJ
eUC/I2YdtqfVyN8uYeOF06mKsddhcbsHGnPpuxmVeloRYdvAhDhPbvONvAFFuZiX
UUHF+0Ks5c8ebSe2+QzwYx4DLhgF5TENleNH8WhjDCF5Hs3D4QBXWlCeB36fhc9A
siTF+2xj1VI10T2JGnANJ1lxvKtEXU21ujuAwePAOgn+UOWi0V/x/fuQJsWd6zGI
5cHiSLTNYaEOPPWyNAdSfODafbkfs90x3LPMNPNLGs1xCH95wZore30QiVU3BB6h
gunp9WcxBnc2TiPAORM9suDlQNgSRFBNwKkl8m4FEDuh27nK0+vz0WgN4wU5PDe/
kusFWYsWC2Ssx46u/u83oMsZ9Lh9s/KuavFYLyRxVm7XcQzOsizlaAIMB0ZEDIHJ
LxqJ1gy9VC9CV9T0mNs2XNRI6rJF6VlVMMV+Vva8bLaSdhhs06tkieyyg/qUxYPB
aOcytyb5fSKKI6ZQh15yy9WTmTHY9+Yq13SsDj+BouchxOqrx9qSiDjfIOrMCQRV
V1LB35w31kyGGxGJuh+soyG8RkTVmeBPS9agzrefnbAXMJb6scnUag187fWKhb1f
UcEvk1tIwhbdEypffSr3k1spg82Dgbifl8t7BGLq86385cCndLqHKmSnJ76odbcL
qWeq9CnPvDJiQ1eoMj+ciX6h6qA3e24XgvjpXT8Ww9t0bwBDqQcWBAaOUsnLegeE
xYpbd+Ow1HGy6vBq4BdWQx4lr/AHGhmv5gNcGSwyXT6ueNoo5HAx5Dww19zJ9IMK
UXW4ciCT8u/u6wuGGOC1cL5qW4K+IYRpIWkqaFk/rD3S8EePT9alEqCww710pAeJ
QrRHJh44Umh3QZflTvJgAouOm5KZD36BS02NtOQjSfMEGRFf5wzYyhid1Iq6LZk7
06Nfb4ZmyPD/rQqyVoXZthDgDf287Nh+9jM1hVycvwrO0rlm0fZqwgODF2Me/cLv
nLWeJxjnNUOBqiAho9fUotfvzybUaFd51CQJaTV5HniJbfzeg7uRUxTCupps4pCX
xQNSFHCoCtEEiACICI08ltY5Mj9TC9Ren/TQNbmkiXWqpw1aEibX69/sXMUwNJFM
syJ+W4B9VfXOGG2P2IZUrexqm1/aFQxZ9oiBy0iJw5WT2eCtmicoeVGxsueJrTaD
sOvZj7gPe6QQHdlcuaev49Ef/5LK4MhNl4NGDcjXZVUA/pPMSI4wnhF6o3cvq2Om
mkMxOUlZQn6lzZbRNVV1dqV771siyl9MjRIby/wyJ5YS1wnbKSqTpQ9yW5Hb4abV
++cjfBzyhvPAJzBub9hJ1t0ftw0PWrkzdptSscQa1BTng7GEJzWa03c01H8ilp/G
heg/lxF7ZLWb098kvm7OyLbk8UX3xvohaLuVhKk+A5DSoU3Xlh2G6MJCt+d1Q3do
T4R+cgtSv+qiJjsaG+BTidXPuvbUsO7GhC16KFRSbTrzv4RkcNWRViZ+RMTncqnx
g7vQyryCYlLQAV24qXUml+hAwxnhu0RjhUzS/vLs+JKRt/rqo9yJI2plyElOGv5w
ZixvT73ihfWKLdHHs66gJjHr4sndw9yaG5iRIlyoNEe4Vqi5C8DPg1HsXKHhLt7l
FtHZ3Ofn2mGn+NWrj8TM/4ijCR4knYuQG5z8QdzR1fDIDXWhNxlic5N1oxpT5G2u
XLEm5ktX3B2ZophFLk2udTiIS/8/3JfLeijgEBmF52uwYLMvg7NjQQAaF8d7WIDB
CxBCtdEGB4FauGhV1fIz7JSZmYEENdUDEe8arihlxiKIHIbvXXF3pJSgMkUvn6ta
PXtifnV3lv4Yqt2L4xafuuSW0UiPCITGCDjrWvw+AGJvwFnR+MDHA3f0wf7DGYTA
miYAHg+bn7HmS1SPfcOXWqRIF2tlbYLfpATEUb6cQJXhngd7/l8eFT4O/JSXJ4vf
FDs4zgpopbTmmwKszrr5U6K99VoZpCzbkX+sfmLQkeFdT4/WQKz9e0X+DZ6c4n6Y
i4G5o4R71v8M8cbVGXd6GvroCbx1pdqix9XCgUIKzNzbCoORwy7TyWM4AW2Guewf
TiaAZ5mshHzdD+xg5JzdXL8crxX6EOSp6lWTW5lWiGjxuKwx5W+MbPX/IMXIrbcx
x8BU2y0FJd9i6Gvt4YnJknxdP7/tU1e5TEMKVSig6A6LeIwimpveXm5d2iE5K44T
7YArKxGhYWbyIl+mxgIApI9/4EeWaOPjmSZzW1ilPhUdDLCSIjr4e/LGzLJiK8qe
DEXA+Pf6ADSQWTIfuYUoxWeKsGBi3UDzNJUeS6BtOYnDjPNzXrftVdpjux1Ec4cu
sY0kKwUL0omFA9L/BiRL4Jpj3kKJl577TgT1mTqBiM/84aj/9nna6vQ134hRPvKF
jlgiMhcVGgopVZf/aUnnJ4GNS29pFQSbrU2JvRw6o8KHfuSh4IfdGIzT2hwWwU6H
OtQDt9vC/ZaP4BHKMusKFaiLRoI8fhyJ5s1FxKou+G6/CemshlG5NMHRlh2RpAwB
RiMLiPqtAf2H2q6p8v4GogpDrVEK8HOu1lVoCPNXYlAh5o6kYaSAzPymLEZNuAim
c2i+fmQPUSXpS6KJekFIrWeYorhHSLMu0wMU0ZCX8WzivpvIWbNjeqGZeo5GswJ8
meNKDHKMxt3vX9OTC2zfQFNLBl73wpOUjX+72UkBNgIDIrHQpuAnHGu6Tvv78pzl
fVACNABzYPPkehl8gLMmgvRWxkRtsCIFYSNT3cz9Kau8FVfhHnpD362eGE3ECvVe
N7xUEQLHNVc+8Ms5hKnVuGUQ0h19AQiSsWOsubC5d44GloFnSl1KoOnVdaSanQrc
YnoguWmrJBplne6qOpl5OdqQnqZStiW4N94f0jEvcWNZ697F1BrLHtNSDVd/6R8f
JI3denqmflJQXxnnKXGnkAh7NR6LB0NlpWJQNx722ow7X9zV6ZaTYyPJB+XIaoJB
wyk9vv73rvjjwc459rdGbUj17mtQNpv3Rigs+D9NaWZs1fuS8wk+KSuFLHz1g6E5
tMaSuvD6tuRAigPSIFx9e4tc1r9gCMwU4cZC6ewHHb8JCplDUfbYZ3LVw77f+Ooq
BS88OE7wlzROu6g3RIMUboze4dkXKhf4W1gKQ/SRAuKlJhyFmWrwOX1XdzigQ3/+
Iu4XECEloyMNJx3sHJPw3nJpUpTAZVkUlWCslc0sIzQeYgiBtFa3FxzlFgex36ai
gYAHqfh8o0STcNTKCshHs18J/Fqq19Xb+6vB55hxDcHusJbY+gDY410ZmA2doOXr
HFuyu1oUdX2ckoeGphC92QWMf7gHR6hYhgwYgMhspuu7i+lyhHlcJGnZ6j/g/EIA
QxOqvgonFK8+d5VFwVvNGCYgjouObjr2YNG6PMDy9+sa25J9H54LQr4ML1BoHdz4
0SsVXaiz+ejT3cR4mMWtrcp/IdhSJt1HUznetpqmWKpKBZLnoYkoqHdMBK+2wqY5
wIzhHrLFZA4JYkK9bQ2Lqb6WWf7EKYWfhFdRZHzoU5TxvLbQ54EKhYb2UlC7nrf2
dck3QWqX8zKkRrg/IbpEvQmAywFHy2WEe6AgxpZizmWWJ0BM2r98xvLO/oyZMaQ+
HrmNyhUsbprS4pqmxSzmfap1c3w/jA9cHRzwTDeh2v/q1vvWfE3ozKQZEOVbUgDT
2R0nXSP/zF9tJWfK/H70tclFifySqvl5ke9RmKTeBE4nZ+g6s31XxviCIvAMvRpr
ORIpx07mMexCJ0hlGiPe5a60kHugoaZ4jzV+bnRuGZOUxZ7Rmoq8EaV9JEaapHre
2WSGqMMb9NZcu67sg6eTLjxpTkX7amw8snY1PKyqCv6qzDEZ+pM2tPpGslUl+Dh5
HvHXgub4+Hy/Xo7jbqSEdKD4DffpC4ECo8VU+xeagr9MzcTqfEif8bNPdxdVmqKC
92RhWVXoMZwqZTu3xCXEI4m8qbcaTMFcN9cpifM7/VVYSynJxJhSJ2LB4k8CMy6F
nsFkMZXuyGvE1jns7txytY5DvPtnNcrSocN+qNqRyK3D60jY0sA1CRGXNTOu+C7U
h0TgSXs1JyulXnlMTI0cg+nmr4+EwwoMIhajmAOxgIyhvzk2/kDZv2/qwusbAGP2
JSp4SSXUMvauayCn/0H0wRuyNRuovqfltHEYc4qqoaLj0msbac4MCyvlJVnG3haq
bhhTbgQKLeL8dSsQhylYTgcRKPE42mHR9RHGxv5iMqftJdaB9ZPUI660bZmuBELD
vzw/HE/T720NHibXTA5seVA7uFKcYDTE3tNG9N+s5/w8V7pUjjcdw+HK2CcEzPq7
i6WLIMr1wnTFyO3ws2F1cRT5v/3fuENd4mXR/C6Q465F6jBaA4OlG0x4nThWCcOK
aJcqyFr+PuAG33NwgfHSJbcQABpXp4HrsJKa/sI3g0nM+O37iycmj1+L9snIjvlN
68eD2ugj5/8Hau0mXqVyhBcvBR4H0d6YMe5JKoZ3vf3YZ1f+95r9lqA4RbmSa8mi
v9Id+SLZFsmuAEzhVcd5WuTetOJfXQmdkj9XhGvmjNBWjgskkaRFy1QFiecM8qcp
xIcBwOMldVhCmQ4PCcd3Zo6P5SZh5v1AsNPJCrOVQ8uZeQrrcNL3YtwDFyyZDdkU
0P5+sihsyP7eCVru5FBdGzEnM2J8GVYNg009iOgz+zMx7cnK8LDrXnSwvls6yjUj
Zw+D4aEmrgLIvCN0hqmG9m03m8q7/SzGXCneyrKmKJyx4eB5CMMMWIO44FV99GlL
3Nagd60q8WzF4WJS7KqDWYCXC/hls7h4wJzh6PBnc7Q7FhwYipQnhqG5fBKcV+sN
IsRo+HKjZjD2VZsDDt1DNYD8tp16TjGcTt3IGuoxvF52QOmNUlBqgQZUsDwaXKz6
i7d7/XsVja7/WtZwoHPvF+jrREyuimbKvUQi6uYQVUcaSVAnatbgd2qho2sPEOvj
AGtsdbciA08Vk8E+2hZKS/u+rmAqeOjlR0Sv2TLvdPJ0C8vjXJsQsHVMoETs10ed
EJ0pl3ZYFEgX4mZFQ6CZ3BbeHQR1QPbtC8e/so8xnS/nDwmkLZ9xOxl3fpev3jSb
Ri/SBjVvJiVMy0tVPGyonV2h7a7dW+KOfOBVou3d6g2dF/LE0ztdL90bqzfHsCxr
ujZgxan4P/e4hcK7t4fnikd7tQSfNpINmkB3xtTTXz+Z8pPxyTNpkQ6/V4dcKGfC
eLQE96wh0BVY1OLESKLMm2sExCRTQm0hzRtiyIMgCmJSX8mXWYLY9UAiPdtUtHNN
j/1Pw+UhbHZMmURFKuUWSIyNIBDcC57vrp+Qq6xbTyEbuTbFnX+ShZNRsp+odbVJ
OFAnaldCU0GDPSOv/91m4k8hZLhUeTXIshQSlurzhWcG7wKGfHxOU1/nYAZv0LCF
LukbYrLqbns+MEwKeriTFUYbkMjr4TMO3cNyv2ORrkCeUwe3Yam0Ti7O2So3tre0
m1O1sfp8kE+4pD0aXVsxKWyh7LR7zbC3QzyDz6Yc5pppfKQ2kd5K8dsFhC8ANQVf
DOdIxl2lyNvy3fWH4qkcGT7sRpa7ignt5ww39Bk7SnlgtiEytzlj7jWCF00pxR1o
fLsbS7/KyI5aE8hhy3K9rDkspyav5XSY61d44+fkIfZwbHQo6KTLa0wYxA2h5rJM
/Wg5gMcWK/RO/xPlfTxmpkPkzBzn/1FMt6JHBuiJpy3dFX4L4Vb8uVdqi6S1a121
BJSPEyb8nrk0clpvmtmUg6Y5I0Vk1/pCCc2Ubl5+S7VZtfCqCy1y4B6u13KF9erH
VBld9H8iBoCIe7LftoZ9qJYnyNyzBJa/D3fO37ZsgzA47BJMk87LhcStwgVFMo3d
qSX+dxKohGvJw+MwvphQ159Wb0Qd6sIVm3yfU2/lih13Fbdp8f4QyfRyAswHzYEY
JFtghEehThoXkkonMvyarVdmPAInT0DpQehENwFpYLwo7590AMyxIY4syQBVFj6O
hkvMtSuOtU85GQj2Z2fn+f+Dx+Ajir3hPKsqFnGvRakSsV9Zvo6N1tCPcXSR/tah
IlUvrwaXMmLctg1XI/63q4Oc0HNpuORg9N+w818BamzaDTFXChAXoxoOEX9Assr3
MNlJsH6BD05K48+Fsu/6di5QaK2I8gEa1Zlnv3io8+bd44u8VSx7iSXc7Uwt1zA3
1UpSV1BXf1pq3d4pKAsrYts+vDiZqcu+6Oak9SwWRhvy1gNURQCtnD4v1+YDxYup
SiEN5l6q8XPXAO+uBJZtQtW46HB6t8va+bOZOSHVwtmu5LVszckAhZHVNVfvjN5g
6Ouu3MLG0JJrWE/I4O9ABpSmoffTWhoCH0Sh7fH0V+5zBuLmczbUewRR1S2Txhne
h79ncopRZep3PgJl+eROnrm7JKc5ThNxLauSsrOPmbug9Q0t2fewhBz6PS6tkTFk
zSaswJVNpBuvhzjA1RsbmOG5tVm5Zx35H7xEkAlX01xel/KDFqlmQWXc7IgAU5vu
FIbiR6hD5hN/g3LAHH3awxIshKOqHJOK9T+6OvhnnhJEtSlutk/pOPwgq1AThuMK
t9/vGgvypIIlaMD8GkFfUHZnbKYMaRublJWXOSrXU1vSQgDW3Cbia4nwcEnaFK4q
fOOGHIkIu9UQEJxDQWyz2V6sSmT4BHWmq5hnN6Z9HsWbjwYX9oGVcwlSd2dO9GLh
xNXclq2YtqnRAg8PhJyR5MX7dBG1QX/vbA5WcHCZhgMM47dHCmn2/J+icCHO9YS8
ZhJQuMQtHYTwh/Y65MM0uJJZuzJzFYWHwOmLS+5qRpH9mDuJuTkS9BNp73KglN7+
G6i655qQy44EQBCQ5zMGNa8ZnWxuBxI3CZ+ArmH7zXyrWKE/YVprka2fsst8gqis
8urKAug891xc8UoZx8+Dy10sCmvJPsOanPGCDHpq9iKLOK1tzxh3i/bssBhIiTRX
aoq6Vsfxsi/KV+5GAiykJLCWG7rvyw34CcKt4cJyFlp7SmB2CzXZHwsZHBowYUS+
tyWSLdrFl5xWRwnduvgiwXEWHWhpbJyIYWznV0gBoJj3A219ER54vGCfEZxyZB10
p836GDJNJcitGwo3VC3RSiVgpDz8WOszf8OW72oBOPCPsfsNFgIKK0kM9Zs82a1y
84TB/6vZkxLJBXJIBFh0pm40b7sHerao0oXqiewonEfcRHBwNaMvevBYmvgfSQrj
dzVDbNu8TT0kyur5vEP1ybLvznP+d2SulA8R26YGbT2NtG4+b5b7v5NEJnF7tkKZ
LUZp2ELBwNbNJYz+0n5+0/RvjtjhEuJL1/MDTGt1gcyydg+hB3PIbs8YFVAabizB
QSTs3+gZBVr6GHBR6nm58TtgF2gGK1VmtPF/xqy2ToczNClDzqcEUtYOwe5udW7h
URZkB5E3em6W/kLGyKxj4Yt8Oy2L+MRSQMu5hX+I+nZdE2ZvGB+cP5+dfS1wEDav
nwv7MPyXlx6xvYv1iTIO2ppOpvY14X2J7NnT/FLUu+7sKUL1pQU8F81J60h8Gd6U
kiAA06zL3btFwqJ8OWYZCZevmQDzKDGEFHph6qF00/6jnedYMoSZL7Qy8xRB5tjj
vNgJbe/KqlRyBh3BT0plxUm9b2E3VAWk0DryiU0YtXKVbR6xr97jSenJ5pIhHj+s
NZqL1tkfzvhFHTviuQ4Tx0D0Jt4GqWG4wSH8j/q39EYSc9ZeJNBfAwP7Torf/3me
kLUO76it15wa3c0FhaLQ36+w44tWZ444Hr/r2KV0zdtdP72hDQg89Zoc9bgAJCLJ
+ILFQ2MZ7s67aM6ILyZB2XNYay9V9OfC5niQRVCl01+BZnV967LOD4fwt0/zTHCb
fsuOftZaoq2LuB/bRDM8YEh86LhjxRx/Qg9rOXG/jZ2LvjLyTEdF/F1HiUTlPH3g
zijpgsXbJJPHIDwxpTsvvHwnb/d6n1PpFESwq00o0tiT9iGyfnZd30RvVHPGr2fg
aRKakDiW3Zu3xhcjRhjVxBOXfbO3lapQ/jfE8XQFD87lO2pzUA70gipufdwnTPuu
/xZCRI814hKO7vsE3AqdRRuccW9uJ5WoMKNcT2Gw+vU00iPoNnm/IplydwjocEes
7HHje97DzRhvnSoZ+vUdq83ylSG8255QTCDTvVsz6ugPnXYR7aZwwGFKbZp+OSYm
pv+8oUcbyJf4iRA8kl65ca6LrfIr+VdeSplDNdnq0BAtVVIFBsB7hC5trKiMfrG9
FIWptxefvmMglU0h4DTH1asnkSKQk7sd55GFtx8PiREhlYgAnqESX8pIhBiK3kvw
e7v/bD0TnAsieMvp42SzDrhMes+sHFHf1tU8GbnI2alkRNluprftNJG9icly39wY
dltfsVSnauipdRQ4Z+YIWWoVfi1MC1d1H+rAIGJt5b+FaHkuKCR304A87tQfYY8+
No6OU/GuQnzeDwLmnQT4yH4fxXrhsN+EZknOZQVEVFthxLKbZByDcoMAH0GPXTX2
B9pGrl1wuZBvRgrdzztV6scHH9db/NNPfzLXL9DwLtThv9fVFrCYsF7GMNaaUlOk
e61AnqImiVPvFIZ6nn+DLA18R6wI4yv82FA4bfdCBTvfwWqH/XRBivL0kRoLHe17
HvpcOn9G00kIZs/SogV8VdGXjjFzxeBrwd2hzsVLDzksL86IH2E+SKegi7LKIT9g
V8oNAP5kof4lKcFQ+Nr17ccdw2DbAueZwT+PW5VkhLID57rmavfYIrPTpv+FpR6Y
geq98Uqd8ELp16Eq8rM2jHbf+N1t45EmUsVzhVisky3MjbOstIanRly175qzM2Ii
RjkTc+MYj/n99/0wEZuoA/8M2XowzHuHMFM4Vj6Kj2l7HMKLE6HdDZaxsUWuB1tt
wkJ5DDtbRU46O7sfsbADrXrw4YRmwyagQagbUEgyUouNSAasqT11y1j6r7+wWgAC
Mnq7TPPqb9Rh8cwJUTmwbNTFvMUOCS2Mj4wd4yLpnaqdKxUzJgF+FsWkY1aKBTnZ
RUi5wBIg8DqIk1FjOjai2N406eym/Tk3F2SL34F+W7zPeDCB2OfVzvkgcySEZtgK
TixjMCsQKwFnUM8uDokek2W7C/9Jd4elbtQLkGdDJKBsL4Qg4u33VZ9HLFoRuMFD
Z6/GuWDygcwLOpnxRvqHlu95p2wnoJCzD5PJLPkl7FT/W73McKUbe0bsMEnwo58j
YXiuTCIFvbfm15Q8bHu2SUMsIYg8gjfM7rD0FGGPUBsnp/L/34z1C6pBg0LNZhcC
agc8jhJ7VnRMv5ajwNRF+REKUe04louifqbwtz2GPLnzK/GB/g2Kic8R2V2xwRbh
2Y1lYOx+TW9fa9OHKTnnrhJ5NgbO68MRwFCo0M9+zm5X+7WnV7mXKRTChyWGD1cu
NfN7JHK4NFt1hN1iSHhGs7/jVpn5Kr+sdH8YKNvvYSU09Ma0aaDTnRawZ+SSjQLy
6LQ5CXbuufkBYEZFvnjVIyrrAOEoHC8HhCKeSk4tOGHKe/2EOEEw0wTQXgKxIL/I
eKWKdjoH8zjzkEXNVPjgj2FewaV8/JCHAAo7I/NuUFnren911GE41qQmC257kuCy
IODsCL7ufPDWORCexSFRkRK8OOxUTIl4XfGJMi0oFJUnju/zhCphCTcYeOw/UJaa
A/oCR3pEqA2ZE2/SaS9St2lcR/P7sTwC24GxDw/RUpSQNj0h2KMeu4ssRJxYm3ip
31YQTo2sX/pCRnacG9yDXby6jusRcxp0lAZPyyqtSPSvesDLBxEe/FAZBxN3Hs6O
dpGYG3VLNfsreKl+CFOVvm1VFrG5ZBUr2nSppti0l3SXvAgKwpCD3YUmAFA4mWPW
8xmm8fPxHk/Bca5KMbkpT+wVCEluJG9h1kQuytZXxKPFY3mzTBtXsj8FCySI75k1
FFI1DWwDjMAUFDubUJrUmPOKsjUsPfk8ONUOCkgu5OKjC+0WJPmvr25PqEihSNOc
cyb9I4v3lahiM8dI+aGfsWD6MIM9qLDnMILanG7GmziYppmbhDR2mOsLhzHFPkBB
C4kr9y/jC5oTfTt6XTP55gxddWcLamxl2JNUfiIhLizd04Dy839YbWKynG5onn1C
NKyt9i/AMOMkxO5Gx/q8Nx00zzE7vFKMtEBcNtb5hh+V7zCFkJILia3+2tHyP+CX
8Rxeu62LIQMcORPy54fGsAKRCj4v3m+jYNRWvReLMXC6iOu/jre6KgTZ5zjUjxao
K5M88hI7JscaJB6FrvLFBn6Qe0LcoMCMNzYCURLBd8ruyJIPLuWayu2J2m8j8xfE
mDWO4pM/fgnwID8pYYaKKZ9MVEmN0099wbGFhf30+hoPpYA/18824O40lVBzyeN7
rBEc2h/Q6DP5fTIj2LZDFJcOIUyrPOqgOtzA/7dP5XHUx6A59EYEizPbicnUZ9aO
wCQ2NbUErmzj8U69twob7uDhX1IZFQmXfyWvHyjX2PgFzJJ8ld0sOn0t53WEKAYH
7drtmczEDllxx4BcjsgJHUxZkqP5x2+B+Sfm7ePZ19tY32rBfXqdvM8xy/Rqr8yD
Tyv79OrEyd5Ymw6sZeYAGIUXEOBqWX3jKVwthNFOJ6x3gt69s0Cpoy/nKm9w8snP
6KruFs0zO2l0fh1WvelDF4+BfwsL3tK/xpnC+DACDfOa2iOSuvGiQb2gy2tq2T8h
XsVlctLQKCTiJhIdKVZ4xJLepw9DmwAORrU7sNpJCzcIatjPTYAMCv3z4+uLKEWg
E4dnUkB2JUO6rvHv710plT8GoWAy1VAEiHo0b9waCqWjpemGFNNcDX+MikR8KuUx
DbKfnWHurDIfUt8cSCyAJSobWLAw3KCN6agvCeNuutXmPK1WREzNmNOe9DbbThSC
mf2S9aFK/qM/Wqf1iJ8eBdL0wdYHqQjowMQafXF2y99MVElOo7hrQGJPM0bC09yZ
HQLvXnleXCLeiL5b4tydcCZzi9BYFrtiLDiMrnn8B9tXknVlBcRrzVfbhbAUaHE2
89xR8yQPA1q346RvIMmDNI8stHZ3SSub3+WW76In2tGQL/8KNtKt/WryCNCT3+0h
j2h+41YJWN8YaNm1aD7Pm6s0uQOwzNAwyqplAdAIWatjJxd9v1w7f+rKl7f83dUJ
c9OoHlldQkW4Sm8yYubrYaPwPjaccps6WtvmClV1ZhjO7sNXFXUlPA6FlAaQEWkK
ubhffPY5wmkAcPP2IG74NQhrEg+7+IDAgYBn9Vhn+qbZLdbyCY2HvZtOv0Fp37Za
HQCtgfa572GRrR77l3b6dg4wzyj1q3HH9SFQ7pHKLBOB2jgl7EG228W7Br1nI0ER
qhMeXGYA7YA0vFSGICGEpnXUeNtE7Fsp0/rgPewrENGemp3798ZnJdSEFx6oFfQy
gtP0/0pz/RdvA5vpJ2eSTs50vq03//bC9Al4nT4a0LOQHho+EFCawCyiddzI610R
3w+9vfp2JgLusWobMfhDov/QQy83sgP0b6Fyox2C3QM+pSSpMA781WmVZru2QkId
jYOUMjeT0ZG3X6ROXbLboGH/vmwWfAcC/87HhaYoWG5kuXiJoGWP4bWrk9D03fKr
LCaKlpMvE1+Qve9ffT20nSGrIzJFnfOEUW5e9lsMlau09kE/bBxHwKB8Nr4bhWKz
7IQZWarxbJjwXQxPOLrQuNTy1tDg25p0aIeA96XTqBS9YtGg7wGFvQ3l75oZ3Lya
ytDGQUM0jsyiiGhQ2cgFt3yJ6VcrzsA98oKml9Y40UTXaWx725nNoBOQ04tqd09W
qml/4kjWcJRE3aeF5HQ+scb6ehCwUF3eaA1MlQzwT6JcNc2kW1qoyX53vzUSNufh
MkDZ70DrdppYVq+W6FXt4kNKi2SLO7KdUnO6i/mdZUQkYDOp2K7EYTgInH+AZPsc
OQ2cgn66Go6z8ALx5XS+F206IRn2Ox3oIWd+AEwMfWQnWO0hbiCgjhLdRTAL2OxI
oPkgohzHsglw4B7UCreEchkWBXYIO4MfRw/a/ql8M1gKIB9X2Q1J5a09qP+3FF0e
A/FIypAmT7bkRkUslaJID1MSf8/zZoWt/Q35ttFtGLfKfRakPU8c+V/5DoZUPRzo
FujZvI2RJljRvXO9FH+Ux98fCqZcLKDunZ8y/2cSyGwaVXjlhWIWQkzrPvFqP4xz
/YPHdsfc+MDkH0CZRPDzzBx5vetq9POpKlUnKMIXDJF5L5S97GMIB5fkkc1q+ech
pOS1owvrWnFNkzEP1VXJf4LQ+HqMSnYtjBD7RhldTcnI/cs8XBMTahLyDmoNh0Ov
hlimdcQ8odIs/CqyKkdxqIdv+W7n4EvG5FAxcvBYC1hd4KVYFYelENEQN0W2C2EE
LBllF3D3gqgb+2/S62HA65tTWkYLPTISGmH4P5ggzHUZ84vGPFNz7lX3hoxzjo7H
wT1xHRyrIMHl2FNs7eyxYlguub8UsrS+i7kpHK1cuV2v6O0A7jPkSecWPKotvtzd
Ai+Mv2J7q/HYi2kBfQVs6PeWGbxct01X8SSjmYtp7D69sAhS/0g9lfsZIL7NEgZf
y0pTY1YwFF1mwV8ZyTUQoHLpj5nrnoabB6EcoNyXWvLSaogiR94154RSHKEoe52V
XvGAUu4eWW0/jiBMhj8YcVaWX9H5BD1Ey0hfWcZk1PyBKz1gqyehsWOSjDu/D+/j
dk90D8Go7WplP1cL/bDnvrSZZyCdqICe4fVpt1pFqR4Oa4IFgZhskEzmKYij/6VX
vrnxzVO6yPuU4a+5QBs9AWHQnQ5MhldoJeG8sRAHit2kkz+W/qGiC3VZEF/+Ye0n
Gd5uT+F7+Wm3m5UPI0stKrd4ilQ4+f9WkLWJLPJ8swvz1phatTbfTxuwWi4SHYWb
XRCu+IoB4z54BegudoSAphv4AbL9+eImOYr+cVCy7+X+dAhVko4olxbCv04g52yC
Z31PgPH2WDXFBfBNwhugnzp3o6Tn6fuCN8TeMt5WejWV+bk/0rpd0BSdwqjHCOCb
Lu3HpKW8EbJNnBGX+yWR08YIKHK1vJ2FfSPpFD2Wfgf8nGmTjqt3cJ1kGSDDHIio
Oc70EdTZW06qTHyIIKPhTDgC79TxrfB3EkewFW0qr3PH1514Ft9ABUoj1NLZeo+u
3yH/hyszw2CzBZDhVtqVCz4qH8JtgtysVN2OH75q/YYwL5Vo9OdyczrMxLamY2WV
PI0bnZSPrLn2DXPQ6Jjh5NNb99WlU2TEVGVFi3aF4V+RmlHs26qdLsIm43qpncQS
LnymnjSaEPi1MBrrEkdrkS4thBXCjVw593ur85hxABynal0GFb9eUfBKx0FDsaMd
MEY5lGnrEcJAzhVrfD8giOihlOmXLO8rBgGl+bCmqLPGB63LcNPPjDh2U0gNjMEv
23DdmyXDnOmtzEfz753hhK2/6Ac4Q2HLV0R5ISD9ceOBd7GACdz2PCMksaQM8JBt
ZulShS9tcvWi1lqt8uQnxDziIE6Aiw60vUKWVswGXAFbd+t2bG76J1N7ocW0e6GP
JlewuXi42OprV6X422uWus3zUe9Csk1xnKIkru6WzXE7TVSaSBtxLyE0gSHLr0tn
6TppsUw6herc7UEbrfkSrAvvAxvBnGWT20j5sS2x0zBK7F4xzoC3r0DHIwT7ofMR
ZGQYuiCBZihrXs9dMuchxBQ5FSyZyRdXIDcM0p0uuSFAlfvLL7hk8hGiQ6q5vZQY
t71yRlv7b5SrjTtrC/M9h2fwFpkHMgzxBCzjSXlkcWLn39a84cl89jv8x7yv8JpZ
vZtcxAxiPugU+XgtspAD+XE6TzfPLf7JV82mSl2CkIxDWxzuotNt1eQb93cXAfcf
CWkCDcHJNv1ag+myMCTi1l60qeQ1jY8iIA74ieTNhTZ3U3XIgQpc/3atmOn74jY4
0OLhMe49qKFdzhQRCRXKdzBU6CaD/8EotA/JzT7j9Us26wRt8S2trOHdX/cb29vk
3+bCFAAa+1aLPBNQAr4jSlgWbhf+7Df1hHek7czj7VPWpmW08CcSEW7yh+lKDXOh
YheRWBbL9inWIyV4Q48U+eKq8EEn7w2neVWXsXkmsIQU37FsuwXLExKIPHE0WGCJ
p0KgLfPgXrDJcwXhruYNnVhFRMs5QVVwwptuKzOf6gTGiPXOncBz3x19aCnVz5b4
h6d4sQgXcLIR7KUY+b9xLZ6kfiFQKCB12g2VB9zvrkDI1FnkCoeAR/JGD0XQdPdl
wQ+irIuy22v/m10EzWqN8suZWWpBzq3gOU3Drdx5K6WpqQ/uIBZ+nbyLSAktw7vl
AfFMMqnEXuHr5X/R+AZ4MX8T35zdBtcqKudQ09QpmtgLDoVPDNMiyNWNzZ5wvB6X
KZOIbIDX/mZ8Yk+bvOHtWbcaOyiV3ymVC4L0qgBdMUKBTynQZ7XZqi8jwcxzfwQI
Xc3gw10ujd+NJDBixtr5d1uUwxZA8mMR1JgKXN1TbI+S/s1wwv+zDziv9SI8xjs2
Widd4fB196n/FGU+fCSrjjXJkRUZTbYhTTpe4h0zaQzw1FVjSvaQC6JHFmmqQaO0
9FCuXtOAkSeGED21ZCRTPe1wDjoy6TC5/G4sHA4QEst2cd2boYgX5A0O+sCz8l3o
8jfGDumHWM/OrfQlEOnIzfzbZ0iHIeXZRNJSi4YB21keO/4DRIgNDOrXEHc5BZpM
EdCPBP6KqVToTV/wGKWsZ0EcngcGd3O2iO1EwVp38Jk6+Lrbz9qc+c+uKrzOEFPP
Qcb/uMSGzWmB5I932QbeB4qEuTjw96lh53FNS6WFwOhYZmgjRJzByemxUaeBTv8a
7RXTRoe9FHmcEeHef6+HL8N/W8GKlqtLSxrbedpxW9D1OPcVmIgoaBBDhUHkR3eg
W4gMGlBg64BPmbx0KKtqst7z1pvqRjHPetmWtjKVky65CZKFBuUkOoNZORBp//Ag
dKDYw0j/9n+EZc3y6Ct9uZu+5uUmvkyrnIT66nq86z6gEn72ZYErFOu8oHa0Ko9h
2/Wlj9e84ovTR9h1qPTsw4shHKJp5rTyAmpZfnf8K8TonULDHLSOkdCzkFYjLsfx
VFS5zQfl7ELW8pxy9GMZ1BksjgEwnthOI0LbNHzmJ6AU8ES6/Qt6eEzu+WQFXSiA
fdftKSv3Lxx27qj0A+rag+LAx9BCKysVQ06kk9dzDUzGutvTvyTkM7422VxS3lAI
1rTZWRQrZ3f0YbxnbIuigOWhbygl34WrtH/0T7v7cY/hWa8pt5fA+vR4oMWRjEQR
iJSink81f1pXfwt4fg6zvB9mQt+IfhhMeqavKh5eGt6mqz1DjVRrMTKKjxcbBgah
vINqQmV2/DDBFEKgtu/kWsxSutYK6i+6ENQHcUCa+9GebTN8GYt4ls+OpGqsGJVm
8fazEGh59Nlckb+316bFrye0eyVLXGzvtKWkZD5aEWeKNLibg0NUNi3EHWG0p/Wh
pP3T/Bw8pEl5XKGdBETBnVwcUyMSPvzxtNGd7S7yma9Mz6EzpBsiKh3ADcP/8CC7
36oF2AfB5X0aOYTfxYgLFplNSeevcrUSCvsEV29LlRzcMdrtsRXYOcH/awaymazt
XqNjqHh/Vqxx+qigVDat1wbJR4T8b5ZQ0gGny+pjhCJyeLo3fCGeU7RrQERz3Bad
Da/G24T1ILAB35Kav24tALcZ+x7E0gEyk7E+mLr7ZQidNC4VZFbKf63yo1S1TWUz
Pwa3xMzBB5RSyJtXMsWm97NrIhMGWNvuaxynoKMRdsiFiE+a9c68YbhliX7oaR2I
TAS1wLMRScuOJd3QLacD03NvdORE9s7mj+YtDQ7zGg8gHFy+l4RXcF/ZKgUr479Q
fO2gy5ubcO5nrzNeJqLhVgPRP7dmKVlLU4YWExzPGCNT5CKeJGR/7YI+/2mXmUQa
d0t2pU6Dd2s+E2jS1ZOnht7HC1Gm+m/pS366Tofv+HRuwAyhVcx5dQqeYRRCbh3r
CSrWLRDcFn74qiNfCP2qFl0SOvMpyFqR4NH4u7i9zZL3nPEo4EkTb4ylTPhwXafw
U/8918ztr837lF2sn98KNY47PZzqc5QVJZEYXNdE7j3oXTPRs+7yz3H3+s5CViCf
AuL+D/XNHQUaiuPaEqsQ4PRkNqSKJWtztB09PU7i5AWRzPtlW8KSsqslTaDuhnPR
GKpbg44j/KMk5IRxjxvcOserwTXqTiIsQPuo5MK91cyL8cVyfo1rJ+xT1dHFYqLk
IX6sFy5yDbQnt936IhmcyvYrFmeJ2rSbQpIAdJURUg6JzhQ0ceXuY1n/TY5FygH3
ZNHcBih8M8ZGxYGfBve/2EewlYh0N5dCOEBwHOdXJ6Ou+kTRHan2mgoA8Petcpa4
ysEdxfiM9LQDtG7s3flJcEKpCGaes4U7dIet7uhaw/wgeVy+7GZm1xxI1WrVCVw7
BEEYHkGgouzZy9AYXwSKxahpVejGERofiznkh/N1fVqXKy/LSXF4pzSTdgWQUsA3
relZ0JlCSTVbo+8zbP/XEES2y3zo5WTsDAEQjK8Mlf/h/UNg1se/FLStkogtEuBL
pbf+BsMz/8sl2APJ1O/G2Vn4mY+/abLk1wG5yRyj4xTjLzTSRJ1iAoiliERb3c9T
Z5ibxk/50ciY0cZYYnoD+QoArw8k96ZzIcajVS0K4mCqDG68XyH4XQHvHimy2v9s
mVUoUOwIs41ZONVH2r+UqfgW0l9v4bqNedAJXRXTmu8wnBzgeQylZC6UamDted97
9cKsiPuJul2tVlfEY0fscrYufrME5DZhxKd7rQ5pNLod9PagjciqRD2muihbt6QE
nKQVyPPrcEBGklLqUKpUbam36E2jvTzjeGyaOhT7uCFqrKUURC1nP4LTGq94Dh60
UY1FFF/XjihKfn85NZwXQENnms1bJu4it/dHquQgZqvUMF4iCLYkupuXPX3IuzA1
PJuD2eL3vlK3tAoZ0FY6BlRUt4W2dqDa56YgATFyyHUDuU9ihYKvmDE70WDciR2x
5sycc98V6FcPjWTF602AQBqKmmbfq/pn+4y76R+NCWXHWXejhx5SYeZ74g2r1KX/
928gwEVpmijqHAG822rozUuuiC32TG4b39vQYuOz8xmRIw+XAAJisenbjhg941ub
Pl5ZkxdPYUVZJWJiqYoKk6CJWurTPrpkSDAzTKIwrtvF0iHQr7F0njPzdpSLJC58
fGqOFiXjcdMuuCNNZKOwVKhzkrcuRHujWZ85CYFGyDCLlPx+5y9TMJNy35fK1k2d
pVPvgrZJ8C1AsYH943XSuMqnZXITpFi73LRU58tdJ02K+3z+bffYnsTT4k6U0I07
kBZWcBtlWoyCCMDdNQfVwe0JxHs001D9YgnZoZk0JHUlOPfbXALR81xRGg+yhdSh
hJZtU4BCJMWVSCiyk3W06CmX54DKG/eRXKP9rZ5j749TYvdEtjJVipF2U5HjBiyk
uSnnjE60ZBezY9Y9ahQCLAonYSDR4Oz5xqXs9oRTHz6hOXE1Af3073P6lVTGEG1Z
RexKvai+6Y07WxggKhAIkdtOIdwUXDg288l/+CmUvdE853x7gPJNRCeA22dMaozb
7XnXFYsUd8vC2m48aU4vNO6Th6LSX8Mm/dA4fGrdvZu8HQnVcjhy5u6lc0SKyP2v
VabPt5nUwN8DY7mlIHozhzKNPDwbKkcB38Wg557dgd6WC1Zkr7Mxxj8FcX3rVV/q
Z2fzd5av723cGVGTVQ556MdMjNpf25/e8Q/n1TjGRhubk8Ak/rmT8Xk+R90yWnTv
iAQnMPS1aN2IuSqqKa0xdTxsP9GCFpGybX5zJVHqWtNKTMDBUU538c414dfo27Gc
Lz4tHhPBfT/3cVaBP2n3t1sYAiSngv8sFR5ZZjrJTAyzMiACG5UI5pk4GiW+OlY7
LcZ6ivMeagRAcfyLyiWTfaDsj1Rc3v6oqepO8McdUMoPn4C5H/3jwaENoced+e87
BLiUtCQF647qK7nzUk9yOdY60WYBrVl0zzl6NDyQzCJ1coAZThfsbui2k6Aig/Ha
9JzoSLLBNgWVFv77Xi6g1KuTI9LuD0IC9u7UysJZ7q6N21t79KP4Y35OofGj7Ito
yX2euWTiwvNogV06w+MBiphZL1My96BM2GbPttoNXkuoyh8XF16Y0USeJqX5eOhz
+yvBSngt4zQn4Ms0zPBFLhFk3dLk/z566GTU2fOeSZLHOgJVwlnYslmYv2Tgd/Hj
k1p4AnyNVYo06+TcQxbSDPh+fEX3E5i7MGyTtMs1KsPGcaXcdPsMtg33aTbU/3p1
SxhcXMEzy+I0Yv0ccHFsAb9Z1jiTRnuC4aukp+Wk1rRWKNxHyzYVEjU0uhSRkvnr
KUW6J5TC8/qy4JwmoCwvIrs5c6q0zrKsmsKhpd4RTMOqU23fjx3govuTpWpmwpAT
5Oegv3Bt0AM/g8kNfcqOjmVmZr3Tivm7rsrCeQOZHe/53/qxNvq1L7KVO9ETVPeM
KX+0mvpf29hObRrcXfCCgKbrPM99N+py3GrKt0WusPvt8eW/VSnqpGNfjsMr8ZMW
Scwidk8T6se1YQq58kudI+ecXXgalteHuY+pc5ieTAeTHs+CHOUUYAwNdAdm4phB
493oqrtjQN8l0WiwcvuxF5KfyfBZ1WaOHYXmpyu2gBQmmM2j0B7G4vsd75/3cZqF
+kScG6dJzQ6N2Amy4jQ1nplcRc5u5WpfITqw5AE3uEKZx39KEJ5cP/XNlKVJcfof
0iOXtRJpB53rXA2qdnFG0pimMVb7S2EaEsz0LmV6XCvoZEYgfn0oQzrLtBAj7ueT
4wbmOQ1e/FNDiQsCBfbn2f/CNzfnUTYlWwGbNvyOrLHmIaf2DbQTU87ISxetNlQk
cNrLtOdNrWQx09ui6DxzT+7bakZJ05taBmsKVPcvGAsSWM4YE8waIkCiu4scrNaY
B5faXyODT8Gexhx/Apcrhs+RWj2df6DhF9iXmBzoa0aiIv1AfLf1VNnNCWBvPtTI
9e1+ekepX7A2tc/MnaaIPvLDPjkHmshbhZlaK0Lug3YoMC6gPV67cvGlDGHznfWm
hmQYLnllNYGBkdMNVpccNu1raRMyom8XJXs5toyhI5RxaTgvspBDKDGAIf4FLbEb
XZIf1tZIUOMR6OdC02q7QvWJ3mrXEE87ZT0ROF4NK3xvSsHqSBOffNvjFNvu4gz8
M8sVp14HLN50DSlBfewZBms63kcKJk8VN5EKka7tAESZwRvgbPmp54i6V5posYfK
fl+EKiCqalOb1TAVKbMRM3EVF1lO5WkS6kZBeCgw4Yn3F46/Ky5b5J3zCBX29bH7
MCXCsZdGPmYDdAyRxFioAHPC6GC6HlkE+/o1ZAlZpKBKIOg9PVpo15m2gZee2mcS
FKCr0OAWC3r9AmQNM/lb+XaP9tSflBtQjcyo1ds1p87MbvDyY7MZmwPvUbfVZ05l
UTYVaxORYb032t6hEnqrdjX7zkGZBxdATJMaXXdjDqzwaGIKAP9CCssHEKz4z++y
w2z7Lqidq2aD6nGiS9zpn4A02y3rippUuUDstOCDYJ4hfTng2xzUL0CAmBM5Lh8I
OxA3lNn5CG586aBXmPpiuhhQ/F3KhTHXEGLaaw2zZwXw4Wol0S/wEeYth2QuCDzW
QPdqg/iFVt115i652qFYId7WL/x2hwMaPGCmAAzR0q6MvCs1L1aAupfLSGrlUAXR
lieuWQYP9BTC9VAqwPfXpKkfW9JaggnZjxMLL/8lS/mfRfFHvM8oBSkwhMcYo5D0
EyqNry6tnmTS03xZshghCBaxOrXHUJPDMFAdJDBhYdOz5hFW2hJBdi9lThjuejne
6EAYsd6EuFTTHOkcw+LIcpu6SyCvPYgEbUr0r8hATjF2YTj3Tj+xvIeUxthpwFaA
lORurr/U+3tQE9HQ0nOpX4hxLtBtNwijzIhdN2QbYzSlIA7OdOv/2Xjz3Z5zfl2T
7vV8xsXiXUf+d7LZPmja11NgviPvaVi4KxQs6HVZZJuNO1KkVPGNbosbVL4XTbAg
yaZDn2g+8HYr+V58THnNZDL1qjPzLhI5z+qwgWHbvhjjW4xceoDz3l/WJuNI84XU
glkY6aPy7XdfXStTgFHH0uY8sTNIkCfXZfZEfEPzVPx2tEiY9CM1md4qhsj2FJyi
1kiPVILk5zFP9EoOGBlQ3pSwvdVtzWCjlUjkGp2RmNHl0Yc0Ld/NGQTmG3RhwseU
b40x9I4V/NZBg+WkiBV7Oth5t+eICwdPMrtjo68iPb2VAlkU2pVSnhH5fP8aIqGT
18gVc4IK7qWxeuYDuoL8ASop6vzPgAaHUsY0pZkwx0/XogIk/sbb8ibozHBlVDHV
xPbEeLpXhVZ4Cf1En4WT63RSoDwjmsyhXQYchniRFWmBIpFboZVuiiWgKEHi3GIr
/ztru2kxO3HLwieN6uElsNMUXcNEEflpK1/p4DmfdFbU/MPq9D3MR1Z2HgUqHTFy
kB0V6up3bfIprvnjCIYsCeOACs7XU2hL3ZPlQ+mI9NS+LYf3yHLaKZlbgsoO0pqp
OIxsok+v7lHvc63Z7bBv5sr3ps2vkdNFLUCbm5qHdHt8sVI1inJ/n4bvfz755LFP
UGRpgGTqu0d+fawPhyvCBhRs9EwzOCcnNByv/att4GicxFkxeEjbS2y98E3MDxPL
C4HIQ1bpZo7G+EXi8gfgFPDBN/9qzNUBD/uyytwBwVVE8YNwjmIGbJgnc745Vsjz
vGlaqtkrG+8VjKWm1mhI90P/Y62Jk/2jc8uCjx6aDlB8quecsub/i3Ozl8R7YPgP
4cOMBRBLygt27VR78tVHNo2kzZohnVRl0NNiLn5ToxN7s3/dyFaPtq90b+uAHUbh
K5gQ06+wb8+QNw+D8qMXezwmLjDcFtT9LdAfcVnn7q6189wkTNX8+4Ejw3DIIui9
f33F/+j6ruKB7rilAkUOPoEz+XyCXcbORHwO3R9wPPSktlYA92dujuTguDjiSRBt
v5Nz+hycZ9FahIvU0pItXBc/pAfR7UrUNYedmLLgsKh3GistscoxzfQdpQKH8L0E
5GqEnziLx8F/sfinsYmlx1ylNKfRT/av4cplwyxv8miJmn+F3HRsLLaqxUpnWi+x
fBnG6aNh4h7RDfLAk1iK9brwk8fZreRepXnShzsYUlvvkGOFnPdkQXPrNASGUwZh
KgbsVhkaVkxMDgxaBumyTgKXYCn7ZeIt9+il4QiEBMYisL++U22jt1g/yw63FSkG
RN+IALSwTW8WgeCBG9ea4Xxx4kCo3QE3HKQ/FpO9rnwpjhWteuNIBD8mnNFWQiAp
2U4Oz9VAOcPsTKUDoNhMXirkrMMpFSgK+/82BxSxpOM=
`pragma protect end_protected
