// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 03:56:40 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
G/vaF+g9NbxFXnSQu2jtOd+0Vuchx/5FUfjx3NhLP3lwRMM4Q+y6TfAInAvrh9j9
dAP0QvYnerAqWZzrVMyreq0sLIhUVyrPgcHDFDM+uJxZS+g5kKYgHa1fIikE7adO
M4OzXCrkzI939an5pJkd2tSLFUBiwZhydPu8mcQSDvk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 125456)
UQ39ZIcruplcijf0zk6Isdvyne66gmACJF/+usmiKVpWeaGpHyjrdY7+W2y7ugSP
2LytA/Gxm1ZHaoYi4Kw1uCTDlA0QMnXh7zuZj800QDgPtEw0xHW6F/KHoLgHOrQN
GjyifCOxjIJ3d1MzAMRsQFBrJhZFZh+mnw6UNZ6aaUCyaAfnuYTE8mwLQcT13BBc
HoaYVC4f5K8J645+DmNjc6qiHm06IvlYMQak6tGIJLd14qx6Qaok4yjrHUAv4zhF
5nSIyLqk3D+G6IvlNaAjm5ANpgLcICwwqQsm6h8KfIENPkSoVbyq4DgHlkYvZpd0
MCMc+dmjJKAyeYg6RUhVY3T2wIf3mA4XuSLbhKE2TgoKwDXCzSwdXugZMRM0uCLW
rBfYvgh3hM5lHbe2laH51OqeAdu5YEQS3GwwgT9UGxNpRUMuovLww0KbNn1kIGHS
Exvtwll7tjn0UpzNbwfGHIAgrfCyvoGreO2/OE0t0SrBAF1XX1RMiIW+qdEj1Jsz
p4oxXq/Vp4reCcZY3b5SxqVYxTAmPLkMTMwfntwMgevjcuwvpUfnMVlAcGJsnjWy
fd7zGE4ayFQShHHZ+0xJHugxuLjxLnhD+FtQzNuvek4tS7CSLaSkntUM2i7s5yA7
oGF1RYboAc8gJoMCh2e5N665Jkx6XYhrhmeyM671zlsUTYpb5xusruMdfVAQhepG
p+yG4cd1bTYWmUHlY/zL3+pCEUmqn5ZeLR4T9qG9icQSIkOr7ReEL7od/NQorKr8
+S6GCnCXJgJBsIUqEZ+KIF6IAnVZ5T2AvqPVuMM6ozlQjqF/8yOBk0l5/3jZuvBR
PCvxzwINwKP4Oj0jGepbZLAh+htlQdF4ZK04GA14frvbbUEUbetNIqgBQVdDyimP
fyxeBydeV2FFvibNK0jH6Zn02foEibDj2iUKEJEvfbOh+gtI4ZGIXkNTn96+Fhvf
dzYLMAmeyLttpyxIE8PuvWVXLK0EQq4pMtOymOpWPdlynjGukQUUfvlA0c/64Lfd
zwdf0kwfJXw9c0If1cgTqt6lD0t1SViGy24CnFJf7/hTwLk2iERbpb4sPbd24ccD
Wcb8MRmqFYWlDYIDvJXyWPmeH0+l0KQIVOESM1dsHW8RNgmjuFslJPmSo/ExFk9R
OhDoRW49B3Ul4jUaptBtTPE+c65yyioKRI98ROO/upT9l4lk68SC6lR9bUXZTpAV
sVm/FRo10WTbineMwDbkZc4wKh+HPmvtjDbVSDIoDwM+50qbalF0HDMgNMySSPJk
FKSQVuHS/BQXP++HdMJZbJxuLfNObspSBSklIBJleaDgja25DzDaQBBoARQAD7g7
iIROgxXy9LekTP1+xOT0h7PvFg1mja7u+dyD37RgoYkPSz1Wi82ITZbM/lWJcYo1
R1UX+cA/tzdlYqsWlgWS3qwouqg267Gt7aP5tPBtGeIZYCa6gDaDGftDol40L0YJ
3xR6PYU54bHdAj0iCIW0QLGzo5HIpgAH+uGlHAGUq+HnbSpJAvv4LMVPsuwVQTPL
6omjdTmFs/BiXVmrE3vteevhiHlrTU92cQXuyX6ud04DfXyJB+og7pDn/EF1+eWk
ZPLvgYFlO+SZ6liKY5PzGISAEyZ/sqofqxuOjPoex8f3g96ncCb+QV6LowCwe9Bj
MnCk08+VMQ7j+y6BJ1HrwOSTOyp+lSzmUkfub30t9/MfODznI4vKbURNv4lGbuwb
u4rwhfOP6p+TzUC2ACmj/pty8+dN5nHlE7ajp3BurK4kiALQFmbPDlpxkx4TUkiy
6MCD09qkQkiQydqYiFbr3HZJZmm6XaykTZ2mETFA2SiOJrEIrR9nIqqUhoMgrDDy
c1WOLARoGBXd4KzQxAbc7sob8iuTUkieaOgWpnZtarPAj+8lc1Berryo/yIlywCS
oOe9LU77L5Bs7Exq9O+8g6lEWLARrfBfcmb1tdeICxQlt3DirFI21IzQvQGmVbS8
N1JmFwZS83yuMqTWV1HQAqTduAdU4RMFf8s5AMeI4zof59oe8ekjI+k6QW1KBOaL
InX3oJg6aGXE2wi9seYreN1eHyYYCUGYI/Tk9XgHkxwRDPlItt1yeBPhMu1Z+X0g
I60SJuGKX3OzS0iUVziXZs2PK+mS8qL25+gYgmhIOt01JjYG36yOHVLoUUc8oWBb
H5iFie9rFkAIgLJTGrTb7P7TRPY/ZgpbcMciX25ImaBM7HbuFAKEbCzLXZxtzAr8
SmhJhBx12lfKR4LGKVcWbYaYhQMsiJlrnD6zMCGbSZKG8EantJBnriP/FXzKk/Ry
oBWold45OCIBz6lX2n04Xajue04GvS7GIuB7Z+Z5owNOR1zx/DwjcynAN0U5ywJb
w51Ta9dLPrIuJTvYGWoGfySr0LplGbO98cSykgeHLKfpgLuk+t1uRY0OQT6m+efR
M5cmWqcHiaaGcWrkt9ssAsuSW9T5dyOsd7jfGOipKoDF7R+HevtWwjkDeQihePii
ViTMZA08V/vGeJX0kDJBUjhdeVFghFpPt4WbodLsR7VNEMlHIuK+dG85mAeLYuAQ
A83vFx5kyfw9fzOKJtgcgsUSRshawM/p/EXlhA3gkhnbk9pR4mmSVZ3/DpNvXGF0
3aqMFl5y7IPrS76H92Sz5L9TtJtyWGI4GLnM2DdKZQf/l9c4PHsLpUxe5h3rIoFB
LI1rSUwg47DZLoAqDhvuvQoFSAwbuSqCKhaziKGz8DG78QpM+iVXBUyr5nAOQv3C
7hrSE7+fVYjNKxqDdOnd9gWwHTN+jDuLnNcZagYnBjXZaHnUavUGcZSekRcc2yMi
976wDdlBDNkqC7Zmyf0olNBOipe9OiyZ5uJ5mlmc2/pk6258SkNh6h2G8bSAyJBU
wk1GVIwALX3VqT+R8RWwtafS0PDa+n6xH53yLD8PcyJNCt5gBcZvqI0jbajbOKlk
dUOB0BMnJ2rVn5AxOhi443pFpihnQzE54nnb4UQyE39elggoFNUcarScqRWhO1sD
vaBB7de2FgYcif2pxTJMjbUu5pRIqGYXDNAhEJ++VKtjOmt9BbynQZxx1DttFsrK
q992xkE58UOxKxRn3GvRJGXiickvEIn4omnhsgDpjyK4+nXc/PQYBRO3HJfsHlw5
uhpKd1ZO7D8iAdvtKcNrTepuIsv3pSRPEG/AQpkXCVvxeNdujKK5VdM795AjHGgw
6GM4JM6m8x1YwqSfHjpeYy1k/xaruuCle5bxCnQItH+uKCV3x0J7cTz7QqjtE/CK
g/JEjKFc0kkD2NhaumteWEzI/anLEsCYg0P1xgUziEoDYlUz2Vfg9nWPDryGf5HY
/xGVYiTt522pCCbfdMiIRy8kxsAwq5dixp4Vk8ijwrGgMd+7Or/UauvieyC/hvEZ
AxW6hyW21QsRmuuK64IV+sppjsxosc8AGZ5KNk2O3HuZqA8rTVx+LVWuC40NjxAk
VMVfwdU08q2+YkdAMlK+sMU9q/t+r/Wos/t8e7udYTi7Euce7ZdNLgHCPIkQQDvl
rb4ZokaPIOrlz01Hg+HJm7BcHQyxL5Nz6XiOXZuOgAVG+PmtIF3gzQ56iCi9Mes/
m4ms2yTvpzHr4/Y12whjuv7isiHMXnAN/UvKBLKaMsXLPOCMM6Xr2ixT7bSn0/Nl
JJQM7HLAv/bsdMz96jhknDJa15pWU1nKoDcR12AVL5cWM+ZJbUlnPPOWCIA7PeEZ
hMQ1UY8cuj/HmczJEiRajHpQ7lfFElnbkBqxa7S0d0FbWWWWB/GAR29dF9dzfeF6
o5MOOhTCeidMi9VaynDB2uOELaOQw512688yaRaBSf3VDuH+X0Fb2HPxBc4YVdvV
FkZkFE8uWKG562CCqS4Q4jCw3yqHtw4v8t/jcRdcOnNw9c1DLDfOGRcZdaCRLGFC
wVevgOczIG7mgljI9wyvUuhEm72k0cc8upftIKJYDgfYZXxYeP3iBOdMvYDX/6U4
r5DxItDgmQ86lVEmKatJigLZldDKZnv+AM/2awwrCvqvmyW1xZnqXKGdVIEG4tEu
/V+hxXDggfBtcPXy68+MV2sCdVuj7vacA7QI5AIEp6I+CIj42Zu2W8dsXX6imuUk
C/HBV4v+XN5777lCjLR+kakM4ZroenBeBLzd/Q7a/1xE56V5xFRggHz0Cdl9tJPR
52jSEOTkAsHMrLTwkCAAlUu8NjtSUO4CPeBc7fFi3Srt7qC727dTboX6ErDRojfV
E/NBLBHQJL5p5RJCI6QCnVObUT6AUzvpFIDZal1PnCc2acsFmRBBPj09qlDjl9MM
yt/MQiBaf/Ew9w9lUFQhtkSzzvEJZylMF01Q4lpdrcn5JM/xPUJYbKL7lXmci3ee
eF1SjuxKlapvDJGL5hAzCHRofMMGhhQngnEO0a5/1PTABlcHHYV98TXOlwFl9+oa
N9WU2AdQAttrrR1bqkuphfZd1svvSwgpmS1qZifcKWVfkO/yF80eVWLd1qSrZBgZ
BSIPnwe5irTtvC/d3mVwlTMrcoPlpHo1Rsbp+XUe1AL1ujf8WEDxuqFVehfrY49+
VE36LWOvKVvKtDn+s0JLo8FG+vbDB01JdYQFV2tWxiZb1pU7M3jD7hMOE2k5d2Kc
yS7NfwUtIPsEhqxTvOHGvSKJhpSvQ7KWX1PktV8y2mQqPKqWc3E/iuDoA3Z9rT8q
+RnepZaXDqFn3mLfvPABsk0JzHZViriPuA5x8gO9vGqbRf384zLSDy8ygj4O9Bg/
qR9E72KgCEmL+CdGkL1dSjThSWuXG2pLV2wYUIlVVgTBPWqmKtxZUbBNW3nbUzSb
oV15C3hSgHweR/owcINSEvVe4AzlgdNvsD3odrUnmLJcT7g83K/er6bA+zwfJ8VH
xk+sTXSxCK69DCS/4zbwjRmLuBxMN/YpaWxSo+XoWo4Wl6Cuh0Qe/EOvC6Z4SU7Z
nH0CBLQiKkaV9YazBL1LhddLngU6ZgD0vuFF+tZHc+NnL/PWhOqVM0PdRtZIuZZV
QRDc+DyNvuF+CZbrfPwHPTK/8VgIJSN60BkU9Wvm8akXCSnI2VyMwIPc/b0OmgDU
85C8FXpoqprhdHvILCPvfH/TPhgk+SGWFoFO8+WXXxsNj6de+0O/P5AzqDqHT6CN
9nq34B+btT3MiCR5W8ZEl99M4/acCx+pCfZM3R4vNcmMkaZscMnL/Uz+B6Tf3Ohm
1wez8FUsFdY6WCpaByrZpdljAWi4sJmTRv2KiGNjuciRZvNgMyMUIGE2H0UN9DO9
FGPpG7V9F/+aMXWFJdjDaXvm0f9tflaYT7ghwHHsGvMk95EjDYuDPKsStFQqCI6I
3admL+bcdXI2AV0ilCNDYBwjUZQbwFav2F6KBn48BLo9juVxW3e2LQf33rYUlh20
nSCpdn19P1TDrQWTfq239J0TySPOnMcWvPlSbRjktbZyTXJ4oVtZQiwNb0chiPAg
odA1TB5KLS0g+YKgFrlVw1GJZV193+SjT7uVIRenp6kBa+7H5UH+VMBV9r9poC2s
U2Hrek4d9w13+T/5KSXujN2KBiuseyuNZM1BRmBhJhOHThlcEVXk9bVDxFlY6WOu
geWAJceSfTXhQAp47wVpZHAAbrLK+DRp6pFythb23JCY8ZX3YKAG7qgz3XJjX0fN
uhkQQbEfkwQguEcFGyeoMYfOHTuggpe6ZxfSl6RGUOj3Tb/Eg3LLw1Lbh7BKLr8d
TF/UqpT0+Q7PHbMdMj93dAUY8bUZKBtG0BGynVPfLyUjWMcza5fLw2K9NEbIwiHh
PxunIJy8fMdVdQuV42v9EnRej6qNUV3uXhI6XkVShpPkMdt0G9gxHLzaRmtU3BR+
s2OPrcz8RXU2e6nHBPqWpmcXlPRKoQPVQQLV73fpO3GGFzXrMxHkKnfM/GDxxGg7
uDh1E57XIhAvNdigdo+KTGafUHENXSwgCbvjSh+fWTk8rQNPyzZda9FZf2B1xzzP
nl6LrEm8evsVjFk7kB5DWlKB1a2TI3pKx+u2HZHxjVNmi0KhhnfmxGg0NrJuti/W
RgPKKj/rYRrdGOPH7XGMPXg7PTcX3IsXXBiRQxTMBYCGpoEUtKXN3S2IF1rNpPN6
+Yn/Ds/uPP1z6a3MPM5fGnF/BJ3idZX8ABgIHJk2SMyQu/4amotkopM6iqzTmyX5
IAt03Ts9afW6d9m095ZxUdhZadxU8l62QA+2BAPhL9PKMIRzLLQ8M7a0YA9gFYYP
fvx+zCd8G9sgEdWmEz6FIFU6rcw6S2gn51NZoAq8w0QYiqbw1GGqcZLZLgMKd/yj
rqYfribYFh4ZH/cluDmoiE/CsVvuDX5wbX44jpPOZarYeKM3pYTMWjcw7zwkPqj5
iZH1xlvYaC43skJVG38oLyBZHnghpjOAXG+Cm9YGCaforXdzS2txaiArAxMiQc5S
Mqi76jViZuTDPlKMu+c+xd3+BWOX76LPJ49OL94xGf6Fhf04rxl5iAKcXWNCt+uq
39yJxa95kR/GRtOpzTYRXQR56YwBQGJT3B98Ugqy8JqwI26cCut4JdBD7I28+qQK
8XDrXmFoegequjkUw+bNgZ4eeCbHz/TsBdLx3+iBbQwJNe3o5o2ysuQOu0ECVfbW
S/L6nyK4gquWJltGpddp4IbfmaPWBHRdxyVkUD93CNNO+m7yw+f+ObcBUy6i/dzt
G39f0gwbtgxsdx7HZUQbis4Eg+HvHIyKpzsc8OjLtkD2FScOuyWIeOdFWhQGgagr
LDlsbOVBMDo84MKqtojq2xZ/rTHUgOhGaT1h841yVXk0Tk93SFjskHYkzeTVFtdT
oTPbVVg20DCO4rntLeOqws29HW2GBSmoYNAteizuqZxYTJJ2wlDtFm4Yzalz9qvE
blEkjllsqfQyGLZSvVM6pqMoJR1bYRE7NWACaQHJEcp5RfztPy8qWpIqjEexeBv9
5ZUIYFRfTU9GFt+niRxmVj8x2E9b5Qun+6g1OZCFi8gQ0MeVyej/rt4kx5p/Stzl
eiKJeae3atDzFlo5s5EXctZ/DikGDVZehDX23BzEPZbm/T/T0JBFQA+dK8KNYYDm
YC3tytsHGjGTLthB4/wTAohAknbk3v9o8x8rmnIsPTTjdrqD2zCFpX81MPkHuIae
K0idjTK98o+M29DzaiG2Y4lZnNYouzYZrYuqh0SNlyhJJBjhYaii22MBPZKc1Ngt
W2cpTpgyHOR5C926NbrZzkpzh1IV4CAjyycKAY/MGc+CTiyMnWRv0SXD3ZJ7WDhu
/+hf80ZVozzA9c9VdXPxz/7thqLDi7ZhVwpmyKGi4Grw654bRxAy+8bklTRbJhdG
SDkwNDHEyI/ou4wApjM/iaL07veIDmNfYYeuAiBgdext3ZwfpaYkLkmp1oeKjYZf
qF+cTB6H5RdsnAZBWx4An9dLyQ0rMOVdxuyaYlXzQ95nobJk6qkgd4oi6DdwC04b
lXyb5QIJjynA0R+d9BmKh8/EIVEdtdxBlhq1/aPDwRfFbLZsHdPhJilOpAvZ+p7S
Wae/KXoUk1aOqWq4BlG40lWswK0p0zME1mZ3uDLY2832GfpAApBa7vEkEaa1ANME
zdwz0R4zCGxLW0us8qZqUUDc3jBZQoG4LQcqiNKzyQEAcvvsgx7hSkBciOmk5NDm
l5fCbfh/nDmRHv2qy0oJp/jkogKpYpOOa7lkZDzV7E6VrxCI6u7a+X5OXB32MdaI
2cxHKI/zGc57UW1lv5xeNvT7zVecEEJ9M7otarxb3oTAe1kfk5v+XHv/saXUTFde
AoikWL78NJAwQEV1ROJJjCxrekzkTVRpjm3CQh5tbigaiJkCd077wcYhqwNu5Bpj
rqbxCbfbrSIxh9dHzp00hkPeIaD34I6omcyjMuwYv+kvB9Rf5A4qAn9cUh32Iafv
I4ch7D26V0ZGgttOmQwWuw5xE7AqXjZj9it/NA2vQsoxW49UbRaFPZbuPZqcMHIE
1acw+kLb4tNipkh/zNeNT97FQHijInhy21+NeNEKCw/stNXUqgW1kj8VLEVaRvAY
Bd0h8BC15IdUoDkIbhkgC2pxDy7j3e+B6suJKJ7KKN2i8iwGvLTY8VZihYtMkG0P
bUmZTHnk6QVaRm5qhyd/+Djellj5yeP5Wt94y0D0WmmC0IYF3iP8wqrvl8MTOCOv
EDy9A1pBLkdOwuBn1mQxTUIExNF9Kn4UhQ94LsYP5g/Wy8cWzcSbJzCLoBvwOTh2
l8aVRI5lbQg6RCXgdWPYqE/b9p6l+NvxaUsdWOzm8825mei1HMnOLymBYGxxS2G0
AUDT74eZAMUaRtMcCVUNLsGBlU5YXJY+DvH9vFzVuRaIObPndJJ9jqpRMalIg+PY
l00rpp8FfywubbKRNaNaNyaJA8YUnki2bpPihk5ZKW20E6KxqaReu94lY/DRpDdL
ZwlJYnO1H/RX09w3smtE0UMFMCa0osLIpdJHcjaFmjRrskJl1XxzrpZxBsUOYCIv
IxC3VPyzv0PauzrEP8lzqfPsw9TC6gPPaQfOg9YKH6XnmK0zbSWmy1cZ9J7YQD/w
QRincgNuzDnLVaPQrZADZGIZv5KOarfFInL2b9UTzhXYznmmjCC2dtkEzfHW03Ly
b6bxDLzCsWW2YvKzHMgQUqXbQv1V1BNhiLMK/snktfbr85hZnRsZ4K+dFBOTpQG5
oOI2WNUuKYGnEifbkDzQxIx0DQB6RkDBQUYIOd6yqP6vukHHR0DrcEAMrMBz+Zep
8JW0Y21KULKaIkOZln/dkb3aYuNnnDi0wdY5BwN0U1CgtfhjVMQIVYkTIESYS9om
uM/gFgSNFYuRp4JlFIt8JwZRewhzt0h7+ux1uyGVocc4/mL2j6CQOroKS2cvt2+o
gF2ELE+9VR+YdhKGAznpCfaqYad3LBAwcWFtDl6j25BxaZtUz56bQoRsIscdUW7p
rFB28PCt682PvFvW+nqTS3oNkLYoGm/xSrtRU2l92IBEyzT1n+ezFm807VBY9juu
i6oowNcEVecLz6paQVKf2f+BgPxJHAaVPR0D+yE2FyDQRrUHtz7Q3dhqpBwjvm/m
68nQXnZqaoXwcHfWuJPusKan7qU+gVBLdpQ8Q/wc2dv+rzu3Uqs33/ixTLsD+Kky
al4vs1J/LtLrLGPcfl4XJtDgVqNJrX+yJ7OIvBMbax1B15JlqxaNbaq1A9Q4fn75
yeu9EwaLjWV1x9dI7BM54J763XMbvSMYLr92qT/DSrPOP0XT5etc5bBoA+H92wDA
bCgdxmFeO8eI2mP2bUCaFReyl6k/mjYF1kXuSo7Xsn5VcWK8hEy6K/wSueKFjwan
wX9iADuLVP6gUIjR7ZCdFaV5uEP3orECYyiKhiiiKVw0VdPbGK+eSmf2axEWf1uV
IViWTuWwbiT3539jOokvYZRvfEqNO98KmXnvfeW0CCM0n9j1gmJHcCSUhmuw7DJh
74xz9/kAY/gtkwRRY39pP+aCoKRs/mmO7yecrzE+/6JQnm4jSAYGolSi4D5yGlVq
YqYBlCXOeS1q0u3/doKDRv58q1N2rsHdVrOGBeDX9tjfDxacmzIzfKoCajtRrB7h
B+0tYehp0jO6nYEiBS7aa3V16jDji7Cst2Dz7Cgx9mQTn3L09C4nUZmA2bweoPUl
VK+FwGwAbvcGU9r1twsb4uf6ArnQc664wYlayJdbgVbSHi9Ro6jI5F4TySnQkif0
Oh50Ytt+jOzwMe+UgtBYCeu0RGzkimLed42PcU4TDQ/gNAqVes5zDa/P4Hg+23Yk
xmUnpNFudEQPX+zhF04q+hUyhUTcoiCIB1rvorwxBb+wsJcvB+ScTqlgngaUEgFg
grfSdi2XJtMqVBiGrW9LxknnShVpUAE3xJTnhnL3TPo1ILCAIhBMXVNXnlnOxLq0
rGmuNON2pzA0GG6iMvylqxPz6DVh9GS7XrkhKoIgaRAXvAp1r9l8oGCdqcNp3tyr
UBoC2AIggcnJlElghfsvSrNlE1XAe1kBkSR4rQZBmc821QWRDSND40M+2fjd4Xo1
D6D6bpbD6TqmwrgM0Q1fOePus5pr0FZbv/VaDBaejSo8P/+HUlHC7nkJCF13r1uy
BzKbFLfgZMA5pJRsmreGj9vbrfKICFI0EU3gek8PjCknQagjiUngAYsAa2S7S3je
SUQvIXLVNzL/twdpvnwQ5YZr97gbq6YFmjsJKUTtSWzrAejFDVhhsyfrCgg/4OXH
eBI7xX6djHj07ExhtDsUYj6LCX6V3FNitubKEKrBqzMCPCbsAFYYJnfAPTlAtjmd
+oSMw49+kwKqnF38uKWPlRXigfs+cmcmlHoK8a/nddNPt/lV7V5YnamZIhS4bQU2
Mw1S/zLKxgYuNgokERINogS+Vp3+F8QkygIQXR5UWCQigoxbSyU1XHsoshDQfKQU
0O2e/C7f9Sq6TpBfgM2cF1NcyjQ2ZFxY0CaXscSTdRpS6eIQednf3W42s3LCYeBm
+fAhQYubOz6ICdkYZzQDNAHVVNht2xv7E0TIqU4EDI4Nym0WQ7+3CXsbbyDiFPTj
JMerirnyGyzmlj+tp6uXptVM71WbbzDE9ePvPRwqN/dt7j7hD4JBtxmphtExY5dn
3GzSYAXpIJnXxsuf6CrPz/ifpbcV+k2AiDzYAc0CnUFtY6mLATmoYWdII3zxBf8e
MD+JQBJtkcU/u7GTHeQ0sXt4jbuprViJGmaQFzChb4ThSD7fe3CCo58h+UnDbupO
z6Xpnwwdgx1oRVPLKQlOoMcpfpRelPE4TpWlAVxdEDFKrhszfGGxKtAKVISWZDxk
S/GoJT23+pJhEOyWY/SMUww6m3Gh7BazbKpLCh6yS6SngS1HOzfBPJkUB0IQfUda
suMHZselF3pHk50vGbdGN9OJ1yxvieRHYuDT55fWIHN5xDo0OiGOv3hfV0/P0RnU
3MMIeDCJbf/2xWNV9ZMqlsT2XvIgJxeVf4nNTkzvMaexidny2lsVGXFiV9CLmx9z
VLzVIDhy8qh0AJ1REDZXDX3HF2Z8fh2vqsToTNd/J2IsvXixn87pXsuxWKwmMj0Y
rYKBzvdExUZGYcL/rGlA+gIe9GiH1fz2JIkNRsIjrwnW8fSXX559dSeNMpBJrmsn
HIs4G895LTBremBxQpzcocVXA4d5dnS8FsDAQr0pya0yRAbr9ll33WpSgMtBh6q3
uO9jSPGVQiNRuDQk4LPrmbnt/4Ecw9Qgvsv5FBIk4SEGZSy28aHOCi2bouhwwhEs
KcPyLsIfwpUPD0oSt/usEDDHyX6Ym1nDvDqzFujLUGUWN6ANUlfdP82cd46a4pX5
9CQcTWYGH5Oc6UDOF9VmcAh9shYZUyIhpiAuAt2HUGG9G1h/BZj+Vqr8tRtpGdPa
FckhVVfNAwf2YlPKrFK3eXwivkW0bwD9XbORxwWhfLlZSvLA3Ie9ymrouq4xAB8s
OXxhAzHIYwYlWorXYke0BmmL43cAtTNPifJS6P2YmeQS+m1yseF8REg6BMdMx0OF
HDUJm0DMuFoQ1bNhKPEU42lNvJQADrT+cux+MRm1bu+OZdSvFS5AoEF1LUDx2BYl
Y4pIxBkp6nYGcBxlyN9l4OWRh5nXtJs8rGJS33QaR9xSrsrc1Afj6lFAlFTkEbwV
YdBkmEAcx2OImgHFa5RJEibKMUxNctvObDiUZzeovOP7yjPpMRSmiEynHWnIcJPd
kZZ2qfg9p5aesoR2v/E28mrVRwedILi1pAlaNo4eeHKq0gz05s5tuMBbUYLZSzMq
Hyj1mAJHzimy16EoRmUQ/vouw91PGNf6EdxNczEI1OH2MkhDT4mx0oJjStDO2w6a
wkoBoWM3hNOd6cn5xtgUUVAxSNzZZvgSq4JR4kg7+01Ya1GqHamd13xGrgzp+RtZ
WghDZWnntcrCjP8EFBNbeBunQv9zLcCyd0ZI0afTwIoW/GBIDh33evL9BX+qM+gL
EO6tDY/zOKqVEUF/dP8PwG9RlbkCkTR+yx5uTAUVa6PFBaRaJw7scdNixt1taibd
cqZ4PQoO4O0Zf0gi+gHdQ6WddDEc/LJUTdbTAnkyWVoOJEWeMILRjnV5sozif3Ie
cEVaSI9m//KiEFr8k9c1DmYlxEHNIyovlQffydlrFZ1Ak+CbLOwdHnOtRxOJPjq8
UUuId3u8xY9+iwR19waQij75Ff41TA5M/f4FljEWhcLiOYWiI3hT9YsxtzGQvftP
TU/ad4qbIzylZ0j0xiLL4TlNhxjjckVK6+dounyJ8BDGXOKETVQw2KD71nntc+hi
FzkVGKI8gqvolfhKg2dV5CSl9AN6i2h95jW2+suFKx1zWVZAitOiqIkzIyLRc/M1
VVn85l+vjnPLhArMCqNaOuNTl4J9rxadCpMzv2V5G3OEB6AAet1vMpLzv9w+Jj5X
QflPGWwSZPmRjjlWrpLpaFE4fYkKeqZxtDKpK8YnWwk7DpM+s0wAbvJ9fxvbeuaa
lY2FGkJYPZUS0OIpOSfRA0qt1iuuymxae4SVdl8V/SuDGWxj6tX0L9+U36dhr8qN
h/kmQS6G5GR9za+Rq2KNyBkro03eBWNAiKocRab2aZJrWtzU+Mv8ukY34i0WRCvk
pQdd5n4mV1x0V45rPpXAOJ2sMmYtXKlXe/3LN1sJ9ZD8hLERpxs//zXQPNiD4uVq
9D+g9MTIpqMB/Ctl0wZa57K1QRvtY2HMqtxxfVkHQib187vip4fuZoX/cPUjNq46
gEgNsmjDaPMRVJ2A8xHyRD2LdIV1qyUFm9Fd71Yd3+4xav74bChrW8uwMYKN31nb
khDpUCjipGoksxur6oDAtQct7voB+5bDen4qztQ3MYvYFbEMQviZwaoPDM6FUO4D
GneS+/37T8DXTJXRO+1PDzZwHGjoqDAlpyrml4zLMwLJ412wZmVl1MIJmKydzJ3U
9SqURdqKGmKYMoOJBQi2BgdPf0+gI7LJWjTZOzZHmRKzJem+BsqOoh7rPq0UwrZO
onqFtWzsaenR69bghcaxLJOluMmemDxzbAwitaRGPO9wXx3pU8fIhXwmFPiotVm1
jdps8gVFQezKlJKVSx5pDVCY0osHNl+/4+S4AR5TG8Cg9LYh4vNeTlPfCva4VMuP
C7CfJIu7lHKp+KMV1zSjIcFwfIcJ4QXCJUL8lOf3bH/OXI+6ITcPALij5JXMPG9N
AtyfYWC/men9CxIy8TLDAz7HWMaB6PcpgyT9lKv56ilPQF8IDU3aTQXYIdVX3cvM
4putsAXi66+z8ITGPC8p2hnU3l00a+Ur2Tz2460hLsPhzu+vZ9/8kDqp57R266EH
+IzGZKzgH1qh3cEv5g9RV4Lve+zvJ9LP2Kg/mFAlH2yL12VjfeYnQ+enP13G0Z0P
0jMz50ELrOcPTA/HbO78Kl0i5uq7WZTfuslNRuEAEdQmx4KIOAociiJO3J7EX/Rj
z6zf/a0IfR+ATZVKdUCf1G2H66SnlP5r49pPnHlNEHEXRXpXFx3c1Kq2/6+7Awpm
EeSrX/HGrEweKzobLJbyttGdL5fscQKRJk8wz8wKr2OtYoMXzaBxeTBXI76DjPa1
8zxb7uOWrBGKySoIMF1QoLDuEjFGGuFHBFKEKc7mGz5/QlnfS918f2gz7BCPOcSc
XanYclRUkgsugq7qyecVJS/F40ZMEWSjXdyZ9uEwSC98QKFUjQ8AywScxuwB18jz
FoOrErTqOBLaCRtWo0AbIArpx6WaVtHMYdS0tFsQRzCJMGlMzdEPIT6/VnroydDo
cScmWMvAKD6tF3I2Mz+OJyT71qe3wk8ssGP5UzvFc8yCY0aXvwunuWmdXeu0WJEr
F8gTah24Fy+WaOhNUtpFw5HKSypSl6JTuOinEwFmkMfbF0415K/xEVAwSTPDL34R
otTneFJqaJHvAlSzYzqDRkgrD9K2MX6NXqIdKNB7SFRt8lJ9t1FaOTlA7tWWX8vz
pSlC+Go+Z32V8dcBikhoqhX65t/n96ZAO6iLfg8JzMxRCFRT3q8KHDVB8gSmFbDk
Vw4kONbonuxqbSoxjgZ/hc9kDuyRcSoWybjPaao2GyEK53IZkPXNFg6ibL0OB7nC
GGU8lyEke1sDLz0AG5LbgHGB2GMpZ0HIsu0XtPfUcNlA46g3WNek8oUXaIpsS00W
Y6+nqdNtoWzbfOXyhNUaBY5Zdi9222vS6a88yqZNQ7MoMjJRp3fYhbH2pw+9nnXF
L6VgXACclDhAs8MsT3rwUb1pPny1scchXbruoF296blyd0kokpVKiKSGXCSmjChG
WOwr4bMMyUhoDqY4gyLSj0O4Y78xNPL0I/9rro/f7/KLejkS69h0UTrX1u7gTeus
3gZstW5KKSYw/ZXZMNg8461YmhlwHn1jZDgo/jaFayHADbcyhydF/zyrToyRpRCq
NP4KXGCr6s7qG5IUxO5j0Now/uoeUNCeVaQSAp55p1pexHpwlGJO0N6zjwDrJ0B/
CJfhnlmhN+8zapqSC5ogJTZ0FF/I1TsluSXhZTdJ0sSPod2w+r0X85WrGcHWXgC4
jRE6un7HKRmfaKIblef/Q9a6xoS1vhlsTcTBL780ZJkEugqMN3q6fnw+xyaly5iL
BoODkJ/e3EbCRAfkM4JUXwATsxtwKpIrJJwfBC9IvRPWh1ojuvEv6r0xc7+IcCo+
rWnxqUUDbkCMTzNCxkKFZz1sL75iiCnRvF9MfyD6coOMnaRkt20n1gpNj8Il8BuR
pgLt0+1N2TJjsoo13dKDRaoyEufVor/zjBZykcSjkwWuVvaLh9OhrT2luFdIsadh
XVWNmRcGm949+2RBj/aubR9hyLidjLpWoC1B/fBT88LHbMiFFWWN6Mwk0UqGXeNb
iOP72WJiFXU3o+aR/ViLUYrR//02Y5wZG0Lp4wvQPsPS/AOh/wjUU5oPeqMPJ/kk
3ZegHlbahTfAb+R54QYDl+25ZCei4Hj35qXkCgbm4aeyoN0b73g1HahJ8d9YG4bb
ySkQ9OnDbrOlvG0wo9nZM8WDwk+0SRZ7t9gpusJ6XTGz1sB82F8blsv7W3Vx/eeA
VISIF+AIoD1CruF4X7EHiQ82e/z62rpporOriOxaP++H9YtKJPxgLK0ahShAhR+n
/IIq7iZBqvMIbUmO6V8F660HFUfyVvVjgQVhvO32jhIRFgzA/218tnUWEgmUkjWv
I7RMLykyQ1w3WQ2ay6D3EGf1p0Qj9sxMMpAtWe6Tq0OWja++AwOmHmDBtJDQwB/C
GgXAJjzT0Zwzav5oqI6bsfYZXVqN1XNVW9EC6xHfTfUvieEotkQVkKyWGF0Us3F9
h+QgPj1llC4zoGqes1rb0evzftcYuhTvr82T+uXZFhTuEahuAMYeArTJOQc5wCmX
+nyROpWT5y9WkpPR7UttZiSALeVCM5ZBy9dnBi1qL+I6SD+2qzzq7JfyuYzo8/t2
v9h2U1NPVIDOsoSheSvaJ0j57GaRKCZy0n+pBLP8mxn9eMiPKGuiOwQyCbezsE/s
AGtcNifRnM+sZphmvIFR01kW3eFPLYouRLytfFw4ySEC4FozgKErjMTtLU87hruc
mgVl+imy6hEjgfc1xFkmzO4whT8MFqAOLHDu4xODlZf8/q2AOYyul5AWHVU3HnG8
XBw9Lz8v22RQAJfMLki2CpHuwnjIXF+EJheiQpXplJoJ8DtV8CMVhUVtDTZDbPx5
oUJYdrQ1TTXf6t76J1Wg9pK5lpvhkOAs8tgA9QV/aNc69Rpq94teEI4R/B50zw56
SjIY3OGJk2p/HkBKpEnpGVPL3tisvIpUFsrbpr2Oe2lHfnEia22ZU8/tOaP87hpW
Hkc3u8E00M97neRFblNLQkXTJMGK6Bha2O7dlc8h6MtWvf05xo8ysVeagDJbfoL1
HoPVN2wApIybchsRH+v01ubdgJhmm9BAtC//8mtwATU44rRrv+RjNnIECOGuE/CC
hJMYcFiHNRpfxAkLXHHmRtATtNLpnHwKoKiejFC7y1hNkkCXwA3fELMWXTToNqTS
Ws4J6NabX0tye5F1Tb7BvlPD2BIzjyI0uhbNLQQgbhVXaJLLh906WSYc7JMlQgU4
F92C5ndCqc2XQVluaW9xutb5Qx6iuS/ljkCD5iYxNao0ZZpWmH2yUR2F4h+rwgHs
Bhn9qhTmz7BSIikB/zoePXOQ30KhmFobSlIqOBqoF4WiU2jNZfIlMOs43LUOFjaK
MpGJ2VFGDdnvBv11Rrt3IqUB7OBz1/i7mEkpT8Zw3LRtAVJ9YcK6U3jA+lX1b6qD
SfnHZkKz3xmX0JliB8GyMnCEKFnTGOF2BRF/RjQ/QjL6wpXMzzubu+LMoTTbWw5Y
e1ktXNkUQ12vgRU47PY3OB/GrmEYGuHai6Z43xmFL2mvVko6HoFwYgceRjRvHbkJ
VvpqhKS2RnRGUfM2iuLk2KlRW8Zf2Fd+RBaThTNuUuksri3jOK59UbBCbxU/VDDG
VTHXZij2WPmF9P/LFOIo8arpKtpYa6SJ+p3l6j2bx0uHY64wT5h6W2zifTmGJeui
N39zlpWrnnq+oqgr5/Fv64PIW2DF5wROE2UR1fV/5o7aSYRubCd5ZdC5KbauOgrJ
WT8XJOuGz/WwEuAbAFTv043IpG6UUIy3GytkUE6TR1j7Bxhtm9Bx/jQHHFoyXEGW
eqgFmDW2kCZhMKB0Xt92jWVPt16OeXyABUnOUk0glRk5sLsCIHejy+4yaKvqVnkl
BYIcCAmSqr+ssWUmVxlIa6wRrowloXXBRfqDts8jC+SmHGSl5991fFdqtyWozWS+
jJlbW9+2vvu77tmHRqf2JcTMmBP15Bfh0CzpalLB2M10j3IZoJkePyZ51qbtnlCB
r1lv+BJsmFawP8dTlPAKo8JLdGIgJwpGuPWU/ulQBqL9vVkUZSfhCG6WpxITNEGa
9D5L80tsV/25nE2LQIfCO4OFJzh5CPKoDuR+eA87HB06rpiUcUWlm4/L2qx8Wb+6
qOnFGFQ5X4vLvLAapbmjsQKOFyD1pyU+4Gm+HmRMUANL5mymIVm0do39dc+Q6+gx
zMO+q1b2CQqX6HxT889qO5MP9Mho3Iy3PA6MKMw4Lh/Rb8tAmk2PdYZ3znNx/faj
tI2ADc0q9saFEkwvpU7pJrGlfRJYcOu67xREWSpdWxO2he1fFzJK/raXd3MNAVBw
OJUaZYeMr+mraMsrT0S9G9oMDQE70fhJZPlSZ0GtbjGTTa8+xnfU4jreFkMb1eVh
w0/rV+y4fhiOiOyiwC5/Htmgc6vFqHVGHPwUcDvGvvJxC58PUT/SeEDUEZxXovQI
/LuXKBodVXHqG3iROREaULTcIwYVY0xbZrgPdkYplsl0qnvAosaAoLrwULdZVuRq
QZ4XAvjR60vEy+mplZ4YlizqbJG+aWB+XZjRLEkQuBlpW/ZPPfaBmFRTaek/sPNk
TvRzFQSPnreaB8jzzdS3n4TL1zC/MC279zbl/fFkOe0Tjbi3kPZXpKpYePWsyo3q
kxDjTu0YE1c/FkwdZuxXTpB05+jZGj1uili4oHNVc/tiEyMgJdFoFzKCSmp5ZpH7
x04K1fO1l2OoFkVUC4Us7IcYAXIn5jF35jq59kkW5UeH5Nv0XoY6k6yrfjCrG2mk
FwlIwib9JAgumP6nFBntclJ5OWb6FrMh5C4DKkXRv7cK98wPXN5l9nCksEyQ3BRM
fU9ew4TzNlCMB4rxNXeehBLMdJd0j3G59K78TDOx69rjBroF/U+ePydZ0tVnPDbt
JdzxTBN7sbqMUylwEpm2ufFOruFaoCH/bpJNG8Bu0zL13TbFxjzmRKe0XpvrKhE/
dZgTE+Hx8uyCtBuTg92D6WIF0MHWrQaAl65P0s+FygT9NJlveChKFDkE4uRTYvia
ZI4xjO04WRMZQ6dCz2kYkP7+MUvl62PyWmVlhoRrJihVEwAZmolhbe0OAGj6U6Qk
ZhlU29pMFO0gWFqZkZfP0W+BbZMznf8xnUrJYLCQs7XTECzcB0u6mIYbrV05ug7V
JjhUoBMnaMb7H3wtOB30Sgv+/4GME6lounaAU7p3zkWOfVC/pSXwiUh98gjI7N1w
FyeDgg4Myx20XlorB4UQmQwezT3PFli9+FmdbPw2GmZPq6fQd2lZnkA7DMe8vo+Q
OIcC60/TpFtS5pkgz3wicP69Xw8PDa7weRiAjQA84hmb7UTh+U9pHl8T38Wm0WOs
BtHtu41kqIcWl9Co4ePH4MPnpWkqpR37ecvMCbIy00/jc6biHiS3qU0sxvohMwJm
VrKvMp7Ln8Rw46xalwPv5nM2d/SITG+HsAtwzNeKzKut/e5aBwAceR03M72dtc0R
8MuEwUgYMZPAw5mH9aX/e6g/80Us+tniAiGnOQKLBn9hcHt9aE3RrdcNQXKhfe3x
sPqVVWADfifYRlUPwUNyxPu2RC7dNeeea4prc10RICK4GW0R71y552FQF8U8e95I
zf/70AIRXwKgxlCpLCb3lQ/lKh74KufZmSDfEr7jdE4sIZDNM57BsGfIqleTKf3g
m4anXrD8501UifOili8OyACSRRmyCQ2o3xXcEFiktNioUcII57EcVQBlW3Enlonw
eyUh/WO1qdeH2XNxieuhipPv3SPGZnbE8aL9reTNqBbWLQjdu2NGsu32+px2AuRQ
PbkAyj9XucoUu1JYviI5MIAGAmnvlDBL2Hgilkdr+xt6geOuj+K7pD0GQawuqwF0
x36iiSFUIOcnl35FaJ6Cc9aZAHqU8WEh/Y5gzucnBa9e2VuIcHvUdKZrWFhutb4Z
itge+ANq2tKZRTQpIui7yDKOdJUIfPb+kMYkdz/SF1mWKHNIPp0hwOBn8RRoepDH
mAF4C3nA2JMW94BIC5nndegwAlWfN/oA6PBzalwvdi8rmH2l3/8Z9RGx8zsCNVvN
XrvLrhw8xlic/tK3WDolI2WdRB2IteP69tlDg8zKjKR/PumTVPYmcbu2KHpcDm74
zWNRNmMj71w6i1aPpcO187enz/KP95G3QUYYECOzjrMHFXgFMooKD+i6cDY9mb8x
UQcByLcua1jy/ZHVScrx5x/Wy5IuauXgqAA4COBf5DvCKlYQCpV60IqxBQ5VBVfE
hc/cafbpzX404wulb5BLL0ENVXkrI3uc52Y9ekr2sO9NJcZGG4/md4sX/da6Nxmd
m6H9eUsnM87tTjx6hz7ESwIiR86XjRsFYmm9+EnMLsVgL/yhXMnlj1H6LHjwgSph
mx5RRSqf0xRE++6GGOx1dirrzR1+XGYUUxWA/NE9UgjAf8uEqcJ7JiyyZ8Yi6Y/B
z99j8KN612pANAOmlYP5WvVdU8znBl9wLvwos0YTiN0zKW//tGateBmqa4GcYfZL
Sh6jLDjZdSYREJQa5B9DI5/DqjNkILhvWmHs+1c7xoyG1pTzO4xbWcDRLC6gcmd9
I5usU0yGcJDkfIw4iKwQJaR2yJCjxbu37gLTvvwRJbRWG15+bYfdI7fGzXXr3X36
a4KjyBnePX4MS5F3DsowCYMD75VzkK0V0llLKvXBQEApidtwYErjn7KDHluuG2cO
YPmyif25g5gBnizsVamNuk6EWbYtIpvlwl6nV3+h+tlYdBA5rVLKtuyNh9ccm0o1
3WzvqLbKO04nS42o77gVX1SkwRj3GEko9o3Je0AFOpqNcpLwEdB5AVbb5YZT87ag
5QRtQr1gg6/rMYGehtiUDVRT4QHdjCogL8Tc4lt4PQQnCEcTl2oQCQjOpQBgLAOU
Eg6eCf9qSpoldME4g0ItMo0fuA8h2t4rPzg083nUPsg2xmRwoeS2sCBAM43xCd/G
BAkjuSh8BOnV903yAmCDz2avNG6Djg5P82JY7QuKcLTv7ZHY7q6tnyZkaNxAjFzb
NGmJH1kgnF1jWiWwx3N41OH7YBDxgJJ7qVnHWIUrYEmyfBNGGaY2b0S2cDCOwChG
EULVbOlOjm1CPc62V2sQSRXqcjc85G0sflQa9TmGO1G13ot0nAuOGqyLUQbaftm9
OBwB45fI7B1u4kOSz9XX6Piceho+cwuvisWhkXwS35zHbN7aQ139UWd8ZvVNBJMR
00MowyTpPZaez+X1OqNR7zkArElE9wmlgPloJYEWxq4OwQueXCyTKVH36DMX3Mq+
NJgSvcjgCe1MbqUai31+lzwX4QYt3zedNrmWqoey7vknv/x/7j3oHv3AfF0P3mjE
/Smvh3lql068wj7oxgWmGc7BlbIfDH68IqdvpziuoRWGJos3xT8KS7gZ74skLzF+
gAycURhuukqgOIolzr79yeyFHoaFNBBl1A8PrULDaqXCcFLd2rHL+BPIrndCy1ZW
owRo0b/j5NyBISMFlD2+JecrkG1nb+FpHAAvWIUPVJgO2B7AAe5eO5MgMabaxDuf
B1R4T0SUQOmOxqm2Z3tZmhb5z2q4hbqBNqRfJ5jzIh125/mFp/lXgZdmflY/JBUH
hezSXDdtgwsbzuy1cMn9I/rEu98Kqj6zNC/FqR+ebTIc7xz2D4OmM2XlKa/5Thn8
eML4xSdBR06QrXfbOKWCc2f0RGxMJeQM9FJV19IdxPZBivCQdHipUjQsFfcsjONH
0QnySUB+PMFeJ3b9WsUIGCof82rDaelp6f4zj9zqAMtC5moAmUCE9HRwjxSYzURi
KtDg96hESI8GyaxNK4huX/sNyvI98zzrHYJQzev5DXHfq5XABw0VOq0L8oQAmBuG
j6cjpN0uMyge0XeY8wE5poz+vaICVM+GyVgay8/7WVhbHf9+j/D0RA7TUJK9zskS
25UEHw55Ak/L6rSdQ+4b/V2ARsmSWSX457xDQXbJv/tc4X1rOrJgR7LWdcWNL7fD
annCvugEO88lAIZhbTy8iINo+EIYSh7uNKQrHcFnNKiIrK6pWlwYa6klxP08dWtO
8+LvPoysBFQClQo/NYRzFEb4f+XXNS5655n3Q92T51YjAw+TcVyXdswxS+v3VUqs
Th3Vc0exAZAf5APs0CjitMu3Z/3rzlvEATSFdc6Ol2VV6XmfZ5yLRYQ4RYfGX4V9
MZfZV5+H117ooAo0tt238cYaTWp1QP0XM/wWHv5bXXdGJDRRgbKtd/tW32tfaRKD
1Q9V3C2IHMGKXHb1Ur5waErKsZaVJECkXrkv6bhlpVMECYSg7hiCV8UYLwF0JNm7
Eq1BPiMu+nj21CnY2O3Nd8zs4VL9DM+nWZ1Q3nDYBWfSRNarVM+h5OxIUJUXTlIt
M8WxOHclSkul0fnk/Y4vS2yFM5EymU5FXeVY3Y/jXduYuycgW0GTiTJjWATpCBay
SrmFQH37QUMSgeSbybgFgWTEKWW+6laW+tmAAbTu7GL0pWmJmxoAjEvNnVNTOLTk
Xhr5oRTO2DXHR/dPP34Am7aPTAoRVHcK/lx9ue5xjwM2GUNitCXzDTLaIiLqHlkC
zb3x/Xi0RqpuCqP1OpHXFAZ4Wo4wX7C+M97EiC+UUj0zx+11lziiNFAZchcGgY2P
E6KTddEkW4MIQNIHOlQ99kyTZfVvNzKnFyc0efdVhOp8d7DZ8TxEDif2ACtnfUxl
VirftOIWz7zuwKxHMhMGUKhMhwflP2oH37IlpT3vwNT042n3Jn0bHepUi34tCAyg
d8Q/2lSanoxF8x3HfDK8/UpEPzwPfw4u2DdxkrdbZCLtHtcaTsEoJk6L/LPxN8p/
9s7dMWwaJNp7OisVGzsO7fF2JbCK5E68e5ZsNjjDVgLF7rSqmw0I1xsMeiPHZ9+S
PP/8UvRfrt0iLnhKbQS1e0Shja94udEKA5cqG9Ov13H4twaVH8DVe6+T/vx04v0s
HN6qKWRGTWmlOlJR5F6fIZBvbUzVEpMwEFnMx/JWmH4nu3JC4qA7+Y/hrpGqnQo5
zkkZ38W4OpHqv2DuxLmXZrnu5CqOK2J/iCNRNTbKiamP8C6YPRzSrD7Nj9PIv4an
axnspSBVqR6v5OUM/2wKtaZp00JHT1kDgmsI42RGmHWoRNE+TBqe6GxJkkEJzUiL
UNI4P93MAw3lLOvrSPuLgzOHoGi/pv+kXZ3LEue+rZ8p0/XXM8pvZ8PlmbsZvorE
fGVdd+3+YExsrewH+oogreXZ6ICltuj3z3/EmoAXQBS71Wtor44V34aW7QQpQrMO
bbLmtBW8JhYsNkIVix1RiEguyT4mWGfdATLgmWUvs96sUogA02mk25LSRbzKHzyp
hk7q/BgglDkqy1jykdCfxhagwhP3QwrdpdPfqLuIbiH1fjKVwwOr05pg94LznGGr
ZDFbsMV8h/3DqiaSa5S+uzjL95DI5wtA9niX1u4cs8fcOhvc2QXrdR3iBHAk80kF
KNGjB+CpWemK3lKKrU+kRF5EmfRNyBDhHaRR98YfdcVWaqDaGDfBbM3gbwf+TGdr
CFfKLhVUlNERJ+IcIjg/OH1R+Z/A9VlZaYDfaWlesTiJhHTiVRIM3MT5wBfJtVWH
44mz7jmEAAE2e5VKDj8YfRyYnRut0gEwoU/8SZUP+KB0BfF1gvn/15rxnNM5u/In
OS62Pkv6QAZYkNPaKUSh2LEKy5hA9R+7Indp1sdJocorr+EQ44csu2R+F0R91Q2m
B7PwCH/jx86EgUbErpL+16lIIh+Ia07D9BdJGj7LTSX2tpx/XaDaY/siOO2ymj1n
oI64ObvbNVGCP/dpHC0wMk3GEzWRhvE09uOf0GTnOEy7ba+umZkikaiw+3o5hBSB
5XD9CtesQmznS7pe3S0Y1whJxUTiQLJtZukuuZ8o02jhGSzS+F4nuXaKi1ve5nvi
ibORwbKKvv97oGN7wFMl++E8WBXYOjI4Dp/Cf0BqQvjRGh9Ea07uC/yVfi/Z9kqD
7ltyZ2EwnOwHO/YZWCxwIrTrKW7ZBsAZNdCPP9yf66wq/vAipnj9vzmdVE/g+IjX
zkKAg+P6girYxwCxNMOwg2qtW3oqE2fko/hPVnNe618eok/uGnV+Y/9A5dqIXiUa
hT6TJVWfxqjc9xqPbVN+HWvvqQAw5tVW48sFb4PhGsB360BEDRKuHGT9Dxkgwc26
/ABlEDG4emcfOyDlXN8Ymch9MDaePBil6zFHWVmXvRsn0NJqjXYbFf9ELer3vaiL
eSb7I7Djwl5vSWGdaEk7suZ9O+fls5JCncHvux5xhyVsp/zdo47uoM7BN5Kwb173
cQleGnSAblNQxcHqBjBJSDlUgeoe2CO2ezElDPOh+DkNc9H614xNZ2HjUslv+jsn
JdJkm2YqdsEaYa9Q7wBQMqopNi28z9+C43h6RqgCKHqDpfF+ug4JaNWEJhMCRW43
biRbw2wBDTIomvFXcF4J0w1fhg1pVReSVsMY6NdLMuqeA6qn2f61GJO48fOITHS6
2G1haxQnkK25ZTgwxSyH/Pr+a7CI8wAvOTR0L5/FaLLlDo/uXcVghqJTbsmmJEol
RBMP7l6GH3ZqQ/xB4yBK0uEZHpzs15m7Av4ZvtcQfRjtRaKChk/sGmK5t7dQe3xo
M+x1Bh7GNLTTzltWzV+0rRbkRHtbPKd3c1KLpQb0XpqQX7pTPzbcrm9TyKF/SRmv
u7eQ77IIWblWElO7dJgPbZU1vxLKHzWKA2Ugg3+fLPxZpwIfbmUSrDS3LoJpb+Mg
xFc/gktfz/7E7vZNzVMktcnQ8EScYTjCHwHOThsYgLR/nVhWnwaBG5s9pnpfDUCp
vcVz1LtUlRWepSdp6WXjzWRDvcCu6475HUo/6pRO5GinQULdjDyJo6/Rxdwfd/6q
ltRchmW5VdxOud88EFk0AErNCZ5cYqHHvf1m3x8LnIcetwcHYk1/guw+paPzzul/
zJqeGo7gh+TF1+r3hnvV008C/apVfbFvoidpX9UyD3bUpU1BKOcu6yR3uO5eYVlU
fM6rq5ua3jJR7ZrI6V5B9rWQUnlZudkHjnNiVuEuVhUM1id9HgqauUD6DRcvAvWY
ckzIO8lVq5AoYzODEYS/FDaetEQDzsaW9AgD8CQtWjaFyvG+v2jmzZ6QDF3iRCKh
OhSvRoi2jUWyr5YSg3wSByfpBUY5dANnkxRu0d+gmOghsTG7wf3gYBPOWebKxAiF
WZCvTQL0bisSkRQ6gCr6efXi6pI6m0Gm9YSRI3CwF57oathxVw7ekQ6cCLpoFnCp
vMdIoPzUYtNgy2zvQZkfJW7nLrf3aRfYU2HMs8SrQ5lUFwlZM7XhVZiyhNMM29F9
I0XMZ43s1YbW1VT2uZdEaUD4uP9Wcre+IhmO9FRG61fej/WDAE6K/DdAIyLFODrN
eoy69BqN84QhtIn8vhWNIuqpkmcUcyhcicv/1rFjJ2BrzTTxWqdJuzzwuGdpMuCb
YD1b/m7heD6ImZO8HO/WoglumcK0HtnAVCWcxeOS7L3E5Uyiv3mO4OWu16WArAKc
F8FJwg+1P0LeCm59N3mc5ijATYlsfZAVTI4s4UMaHlVTkdftHhrIlwAhDdA6c1NU
n21Pf2sEZwUgs/W6a+kGVhpvLOCRPSlVH5cgtJyLBZkg8PdFMX7yqMgEOaJfixkP
bz012GBEpXA8VY7vW9u9H/DyuwlQ3YVoBmy5OLcka3IDVLnJXCsmmMW2Usq3scjV
nk2AgZNxrNd5EXBJD5rKBZJagDI4Zn2Ja7lWCaNv23Px00u13GTVH06u5XeX1MD+
a5OS/5J/dEnaDS1eR+vwHDVSgxbJMPScunLBvw2WLSPPKkIswwYv6q011/L1wdxF
/letJjP22woT+Dt+OHX5VclyGc7Vht4En1RW6588zK1EvRVO1BrSEMu281ZePq6t
NHyh7ef6Y5T2+HeJZ/Vmdc1VQSipIsBcKOq2CsZcMLIWbpn0lu7DwwXW95epv533
mjsAuwrj/gY/QSjrQIsTJ+gatWh4AGYMt25VlQRFOVZTTWRHSE+vjCSegXMMtIxA
yit71RdL+Q1IfH1fLe5rigyyGVrE1iKcOfCMOS4K0xLs+3NBUvfzIYtKPgzZV21g
E6j7hUuA10NXLueKdj4DdHTdmfNo1Yh28GMuTRprT72aR+6ivc2dhOKO9GaFmsYa
mp/N5QTl0IPC0UYgXmmd19+jakSH9wfy+O5GkgR1tiOO3H0WLojQSEOfbUb9ocLI
MOPRJVC7LEc6CBbCyFc8f5kV9fOIPVJU1oZBAM+t2kKSf/e+SIJK63U1Z0l5gvLM
cMIYPDXyp98IgsDvGNUfyrGiF0+aDQU4IxJxgYpxGxqWg+YlCls9Es9fZGD6JmMC
O1Ceg5zm33yVb2NB4KUEvJRgZ2/OeWg79+xxOwS4tIjxbW4lUsKKp1vaqN4Cqvpx
/UQkj5WmE2pp30gitO2DB/Q3zSnfBO51zUCBkIcALbD5SU+AmpzGjIHjBwDnUqqy
5VIXqghEYebqAL3xVkufRvtvl0gsTJQYmrvvaFRwyWPt/L7cPg2hm6yf//0GH4AV
/Tnc3UMlu1cV6USyXeXWIhTUt8i5q3YpAKBPyxLpRic/yYf+A+RMTBIvEDFapPNP
QvP+8MfOvSe+i2Ir5nZGebGqp2Hvv9VAG25FVP7zJ8IJ9RrNhrpzStUpCE6FhpH2
1zNjHOUOpLqkOS2yKZkrQcfdbRbVhwEjT86aES1CaMaF87hA9JQ85E30wdza9I/m
MYteyyg5oYG2KmblM2sN7Q0SIEcimbNkvSSc0WraGMpHRFx3W7Fr33M9+ZwbRN7G
SX2TDOvzpnhMMcre+XxeChNkQWp961fIpRgIrbeVRShf08Zrff37pTMmilPSn+df
JDHxsZvx5t8amXBg+WoyzsCBP9N71Juh6lk+amRWMWDpDTDzi6rx5McdMQ94Igpa
iNnynGgwPzoD3O4sLDNK7GBab679JUaYbg5XqSzTQy3n5/vZ7BLEi9aFT0hmcZme
QAdJr9fcrmKfE7VVg9a6zQpLwwO/5iqcbgNaCqnUuc3MHhSVy9YEdNKk4CWVIg+v
h/btq1EGYjS0qHzmHt050FRmdhbVHuGbaOOMuQAwNbEQ/kA2LNXAOHarC1+t7Fdf
wIoJ2aV7b+BLATxFxkhJdIjGmqBgmqe+K9FnrayAYzd8FtQ2hf3ywExG4KR+wwT8
d1oR2o3oVHHucQd4rEVk+0gfFvSpOSpgFDf0oV+BiItV1vdRJITtEBnnx75eeR6f
LwTqGpAjEPpOy2phtkf2pLWPb6nVRqNyLqo1hNQT4HhzKaL/H4dOr9xgY/fAIUb+
v9Dg8n8CgeMXUs/1lgM9x0RdtVeZS+m8eV9zNAkbeMHeLYh4eJDr5R7wnwmRL4jz
oyDD4PTd/IoVENaaZ11bdgLBHh4lwyj2N6C0jiFyGv5EFrNljMitV2c/79NRr9Bw
ZKag3LhbkCszr/dpeI0DP0oIU699YLd97Wczg5r79tG9WkZRYu+LHKfCpesxdfLM
DF8ZlVLU22qaaFSssBIZ2J8vwE1YXkVjvnt/Na7dKblo+B8PhmXQMq8xOc+0IYVN
LAPnoUksa7gADBKJUYJp+u0WbT2VncG1MNhh4bF2rC1AqOH9sgwkCDaAuG8TxhQ3
m832FwoBOD08QS/8uhqWYMnHJuaVWXF5xA7cXhpgR4gKfphVX0eLpFwZfCud1OBU
L1GGitRPMVGamPkdcLSzN69wJtIKGvoMgiOi1xpgtzGFTzrJfzf0ox6UMOg65Fay
ojCysx8kvaVFx3mGFtGBbILYYJ9TdlSaCdyI0saPSkFL9C8k+BBm/H9Ca+O1POSo
SO+RgXawUMsWxZOPPDFj2lknzPYWQ/j+YvC0X7JAEXba2dr8BnyD3He4nNEnPtD5
iPcSOGw0I4uU5ZMuklN7obTW/QEj48lKdIkBD9+oN1ATi2EM2ioXGASzapD3vH9m
YwL8yhEEoHKw8tt9TWXjIr5d/enPs8/rdhrZWmmMKSk1LL2NimI8fL2A3dP9UNoH
l/f/umEnRwG9KRvmKR5R5zdO+QEJRJDX3srOGY0r+cD4/9XNU1lPm6bCCeol5YiT
0xixzw5oZJDry5cWVKaEvUeuL4tPL/DhJ1mKNaaqrmbC3X9nx6yFA0LiIJQyGjQL
lfO3kitFMtuKn7nWIXcV8CE7gpiv+4uPsNWmuq1BJKALvu6cNThDlCzklK/WXLOt
LT3BJXCK/VhDqvr8Y7FQ0iPp5Dg2OrBu1d9FUBIHEcoI4+V7g/6lSRlqJxkpGywv
ymX0x8TO6Bw90Fi5zxSSTXQXEG8/SqzkN9lKnukJI+Hf5iMr71QiquUB6kwegJSU
v6Kg+DmCC/p25Ato4UMua7y7BSR81edQQXF7TTRKaXyoO1EH9JAnh/QdaBnGJsfB
3SfY19YPdVzeq3XFdeXaDNEyD9v3a2mTuyoYLtNw5o6DexeuGWQMazr0RbL5Oc0M
EDM0bFVDnpmC2Ui1SXHeU9aEQyOSV9fH7JOwzXrPkHkJmbpV3DqqxA18xKLgvU7P
ZScCJTS/d2Uxf9GG4evQJ8qf31uqxsNct4bUyadejCgEAI4VjQo0+Isw4OIpB4MS
bvhb4MoOxS/Bk/ZV85PvyLHVehE+16FkpGPSXgkP7ElroxfVBNGDT6NCL11KzIiW
FvnBeOhR3IjUVqfPw5GQycRZmjOZh4DcOZA+KmSqihLTcop3Kp08veg8GkxZrdA6
q7FMfUX6HI+p6zTEQ8ANGdGzEJ4FtRWUfcdgoVM/Ya8B9oPqS3mrgCJu4bD5RFOp
kdhgt0NKxZ3+qKVt16AGVxgd0m2xBubME7j1sMYTCPkcoBcx70lR+8gVv5cvZccf
3IFG+DcdwaWqAZFlSeGIdybbkdEpzqYpUsWSIejIp3BQ3pvISRVI8sCkq771SikN
aRC+iPE4nY2WZATxUfbTJSOjmd2KSRPt/q/8HhjsnB2LJbPoSw9OpAWiJ/qXVkO0
wyr4eldw6v3/OiVtBiO6Gxp8k6/G+eEZIP2BfXJqtJLcfc09cNIFZzuVPXhuxUQg
CginhvPQUTeNVIyO6I3tfQfisx/CudcvCS8Q6ZqVlfBJ7yAzZOdzzJeroeK0CUW1
DNa6xQuNvucb62mxyddQfuMghUryr9KDUpLuCFJ9/4eiwvPBfj9hxgmGvy+I/N8O
uvz21Q+uoCcVh/vxf/zl5N/A/EThmZWzAGj+aGJHnb3p0ao1UFFmoW9rvwZ/svrk
qGp4ugrHvF/yBsSgzoI+elTk2S9o+je06OK+ZlVJuK/znc8MJodzbq5z9MFXECTb
l/R3nsmW1/4AWetETg5UVxhEtFIgx+lX62LEm82XZaFlcdTDmWBtI/zE5Wh362AM
aP4BIsJWFsGJAGPWD9KqZRfWWk5rnkuQ8l2O74lwpmmlbuRWAXFJWO7fu5rOIuty
ATnPdv6bMYzBP+RXEsfiS/wZ+UgORbKkNhWrLqaJWld5CY3r5tbabY+9GYxm+y67
3QT3Xj981sVeklRxEPKidBsDgPeAIfvuQQ23j37SiCuN+hBZdTp/3mSKMZWfZ6m2
Vr2/c0WqWfaH0QU4xqInHqNy98SjP3jv/nL6Oyk9HLGOhX4eBmfcyGWf8YIdzy8N
+xhbc6OE7JrMLa65UitmyCsg4XgIF4jDWT79EBRtppFPLNU54uLjYFPE9A6rL1kh
7cGi0Ig8yfdPH4/83G7nLkl1PuAgjUYjYFsg7p6E8vPRP+hrXBkOJYJAsx3hOyg2
HK3iGOcxNjNjZTGub63EdbkXk/b2DZHkpQtH9aSiCAXP+YFYaTuRpE3jMqbbPovv
aauUNPF2hb1m35fVPaUuO6NeKytwjeij38jI1wdPaf2yJf3bS80F6X6f7b3jxtl3
bpOcWumomf2/CfUqDG1FYgMjNfzkRIrimDMazwKFTDdE5lMWcgD8nYN9ovhyiawh
EItpIB+u6RRLx1svojsa/wM7tygCe8ljwgzSUUtw0h7cFIuHNbrqdRycK5uAh/aO
8BUOyxCNRd4UdqKbt3NixbjRxj9w8FrHwZBIExd4JoAKe/W/STYJ9fRDWXJL5/xW
ddqyDgbusN+g5O6M+ZjAUexmXkdN5B6xTMTh+k6efJ/Npa7sN1HhBjY73h1AmExw
mPQz7aHTS7hyBvuO4ETScNn+jvIC9HH8bM8rEoFRwep/VnF8Hbp3F5nO81ZX5iIQ
vNbgz/Kqdz19B89fDAlnO8PjMXxfpyulontVUIy42gNRymx7EKImD0kBkmkJCOKT
dj9Mo1+iUyBIEw9/Ppo1QqJdNdMhREsvnT0uQ9LCNov+nyMyIdohHvG79ZwOxCWg
7V2FZOYLZugBMV9S/OeuqO8+OuAts2Jb5Vjubwxs4RRQRmSjwvYbEXzmLaUzWTPZ
Aincm0nsiqQvHxB5lTefkZqoYxEa7n/AAuVsO1tgzLAA+GXbZd6vwnwj5kz7zeGW
A68wsCZdfWDMp8B/XLUp9cpxZIt8eCnCSWvjKLWLXKRWwV5pG4Qfl2rDaVHAcwa/
jBZyjqL+GPsTjg/5F/i6p6WjkSXrkhs0eT3Q9wa4Tk3MG6SJamO254TrN8h0VCC5
q5GgKPFV7sxSlo1LzxI+aaoJ+z+KJvOweJjeLHE/kzWgzn27s7tUnKeeAbYarlXs
dK8z3hbT6MGjYVGWgV/ZvS3Bnnu1cd+Lk1vgBHya7RxjmI55FZbvyUTZkqlRvtTw
ypgBlz20stPoffXjPjTlVlQeiIB8OgeGM67QwqxmG33OPfEj9xJqoPUeTNLwF92R
lRCJJML/a0xCosy/uDNvnUC7/EpUGH5mH8b3PZGIOARp6AqrrqJdN19A9hlA39z7
DcDi6DCoYVZ2MagLl3Vpnl6jcdI0nK4M+Ao5zAXGep5kgZbBodgxo8hltwfG1XLR
8bIldCi0o2jmOQS837E59VBSaOleA9p+Hs2cVgysXZhZoM9t76V+ZZUNVgM3RHaZ
aBN97WJBhcA/yFBToEPCG+BPzyld6cKqU5M01kBDPBwT29gDbu31FNW5hiwzy0vb
+ui5Udk3q8VdRzL8uKguyKfNGJFTqarpw+4d+/9jBZJDFnjD5ooiFo9HSHiF2cA5
L1bqE3RtOkqWx1ajkMUzVg3OMylVJzsPfkpyvZ5vGbweGb9v66gj/um5+GqclN3T
n4P44sFQO86Xpto+svz71FRUqj5ni9Mc+kEM+qfCnsi6tdz9p1hQieA/DCcRhzmv
U6xAWMDEDT94yBgFhUJyJhQUdnB0Pp1POZUQnFftccZP7Jvm0T+9GVxl3RkNu93V
Lv9iHe78jCAE5mjlX/iTA02bAuQNuO+YHBM5tQYFdFNwVGpAtxQTji+2QUFjnRYc
MsehjQLOnXGfq7cr5YDYD3Q9w0u+bTJ//OIHwMdwnYgr/mdcyw9qMXuRS7ZngK1q
vcJMC0EoqT2QaH/n1NKpZxSz2nZ+SPANgssdHW3H7c1SHlYlWOjknQeXUQ+c7eGM
mECnGCfEzbZ4ViX1QCM+IjNxgrlCsikdXVgSKeLK/cfifTwY8RnDLCuUFxGZfAox
Rm24H8k6+WKDcrgz7xVUWdkRVGwRrkiBdlU39R3BKKQaSMc8pUZ5KJxx8lSDYpud
i6DVJw+QZGYeWkSAKw7kC8Z3xco0IXzA23Cos/Qp2rrT7KwdKCsztRHQc/HiJHbL
Joe9xvyP4ltdgavtXKtRFAUxCh6gaNbYsN0gfQINkENQk/TKge5yz8F/l/dMcYho
Gen8WbTXohfgVKb+QY5V7UMpfNKtxFddWm0l4pywvuLIH/W+LptriTD5ZxL4fFKz
UZVGkIBc1bfeL3UORTVSacP/J8rsNKw26uBieF04uZpxSMZJUrunjnpyIum9qxKV
0iphsV9V9WwvO5mOzeHT37E5gfBufl8LVdMXCd68NiQK3RauAaJrYAk5dyxOPsJf
8zSy7Sz5SjFI613kkxw4sjl6lwZLO0E8vn3LzElL1OxlYNhdqA7Ygohech034Hfa
k3/hiFh2pm0kP744pQ+XcJN0JTGcB520hkCWdwnQrOXpw+bq+8G8D7FvaRNfFdXd
ZLrt4GUjqTNbLmjJF767AePIVqM7hadIhgvJLf2ukaT2iIu1esSFvWoXtvPqeN2o
pLx3qI94QGEWDfEqGI3xFMRI6tA4IhUxLMjOlaae8uaoohQfFaNKcdhg1yaFJ5aP
w4JQY0BSunxU5wI/QbdqL2YcnaG9J1kmwcMDJD4wEQh8fwY8EEhj+CcCSgtJjcds
MJchnJWTFkjK6yTrZo6r+rvM81xIybI3eNsBJZkUMY4vXbysr9Zt4DkKoNUmrEX0
Yyjh87UNj6BlUqACxRY+hZWH8WKbIXJ8r6hVLkscCNMwd/yNG9RlsDs7D2CztTLo
RBwMg0xRi2ggDT7gVvkqIkz5riUcNWbxQ+OcIk4MRcRiTaHhJNnImOkMOZjB1cCh
bPmOX6nHbtF9MWJ+euQSqDMZbncE1C9T1d37NImEipM60gjBehlj8JSqSN0YBGWQ
Ev6f9pmWPHEBN0tgalB+BPmiLv9vcqSOG0ENmy3Tc2Eb4CjtG9fqZP27TVI+YvLZ
NoMyPwU0to3ixp0CMljAUj+BjPq9T7cmy73Q3eO9y8GDroiNCM4/ELbBX9uCHwaL
PljHwop1nJRZfswXhi4kpvSyUKTwge0oYVMoffYzvn3h7NUyOJBNgYJ+ebzIH4D4
+CefFt++/RGT/tQDdZTfwhh9N5M7nd41dD0ie5g4fhdW6wy6yJVGmNA9Zgbc7Nmf
9NNTn7GaGZDND/AN1xI7Eo7il2Ld9052SEN1vZCQUIMWQke90Qu9nPXWsWcF6bMB
iTf/VLO7rJuOf5sg9nwKJt0DfIfVJB/bbNEgYca8L3t4dbDODywtoHKMEn84AES2
Ozz0/EeloYo6NA4QbLngHoqP99NHDRPea204NkeoQ+tQ6ZWoZrIA387nziR6DwHd
sqGyQeAaKP3lWRTmV5PkvBJ/7K9i0+FfDiIrV/G4sWVSQZR41FJc12lAtp9tea86
jSEr6XDS/B1hbu7MIHgja4djk9muQNt/tSjS+/m91PcAXmHsZtocJbkmvA9a7IQS
Ghp9vj99Qqo0EZuaDwzPjorDBbMqcUSULMx1CxQtCF1opC+QbWhsfbayVkwqQJsY
WrANUKCgnJWleomxZC872nRGr+Nti+7ZA1zSgYcL6ILLPWDQgZS/9LzCFDeR7p7U
rckzdG3bKafBXcg0HnIxbeevIHi7QJU2DnycejKQN24tCDeUu5Cucnp2Yu8bLUl0
pjvNduxvCuAoD4ylHOs+63QhFyh8mx3K+Xl6gVgzWv8GnQU5bKU8jaErcEPFcYnJ
v4Y3489E2rkzqyHfH/PU3SjETg1rGzr6r9wrIpgmUMG2lAXFtPKt+TCCKuzZVDrU
0Q584pscxr6r8AmmAMVTO4nb35PjDei94q3RzRx7uefD5/U1JMoeCjfSw7CNJbuO
NoizTND6XAfUr9Q+dUtmFXuehacdJ9KEqJEPX+zPcwtcVrqfFxfejkgP7Jk7d8Pw
BrrbGLcbvbSQWBw5bzI7aca9wCCWGvZgTZP4qcslONslsSHzif7jB7VxEYMyAkre
PwXIqikUCCGvmpW57MQJ5ZVpiSztVkIRzqb0bqN30RakLveUW2hfhiFVk/Sak3ue
nF1lKvoGXNb202e0JhDoUKEO09w6gdlE1uaBgQvS+Abfd6RFxE4l+myydpBuKxkZ
4kVoqUV6Nof8Cek3HbHyQ6N5AbHu9Pnuc45ILKvMCwBpVugr3S/G4Lq9FC5Kgyhr
ODtbPd/jtgzS0g/AU8CLaEAc5PMKxbAd7Q7E/mBGHQmZwf9bieQ1Ip/1yh+Nn1cF
rHhwWW+KaZ7Lzx5/+59qeKzT4yNUs0DO/6VpG4qTn4x9LpNKI/deCg/Rw6ZM459u
kRlFWiCVcwK+8bbm9GAeXjjFqpiRhFMVpBLKKYDsP8pmUUF1T2VX7cRS/zLiMa/K
B8g7FZ2uWTX36TK9oqIQnZMZaj311Xpwxvr8mq9qpzU2/fsRSABZK3gXCpUA3TPT
2WBtZca8K3V2u0jNfJTBXYA1YlniF/a6xC+QBqOXhrIFHsZfFPquGHjSznP2yQvH
1tPaO1CPd4CYVjz68sihW/hKOHLxppAUCQWefmFygc68XQaoxcYu5/C5PGkumNVB
SbRi1TWjAFoq4ZKB2rZ8Z/vdxKPhzfW9KWrydqrS1u33Iz7wjFrRYBZSVPQb6fIp
Lp5IyySRWe1XlYmlwZ39+G5YLX3qO8pyUHYPYNYtOR3Op1OgjS0oKw8An/DLHNwQ
sHBOzxSDWd4rr9Hoh6fqN+ld2Aqy8BupgUvUdya9FUfbnSZU9WvoU4JCXND1HDg8
G48YPStYLPUZemu87KkEaAwfmie1nCEKKhRmOYsKnvhFwmQOuY+L3O7FcOVTECpU
AS8AyPlVxzw6YllRY8RmxSt6igTTe1cTHUezNXpqaTGkie8z+YWSq6BgcpWqZX07
1js7Ixg7w28x7DvYXbb3u0IRnkVEenUP/HlrlU2sBv9ll2kWGIEi6OZgp5bl3DIm
ljEUYfCXi26cEokpBzdACP1R9LKDTZ6LKTX9C9uXGud51VSjJh2b1AK5kmk0lAJH
p7fEMWtHNaLwHo6YQ0AFqjIgEX91lUJDzxGPkUANJkhs/hYAwbubTfQSPxNlNDg7
7dX51MlWZi6gbicpEMqIDqdyjeT1Knd7315xUirdQYsIKpcFpDVgLZRxX+dlp3AL
ErXJovnRoyzQiYWr5YFCObkrU9XSzYCZhJMcNpF71/mQuCz+Wadq0ogz00hJriA4
wOt2UTdZuF/jZ9ov7h5p53QwuaZxkhqKXb6HRha+CxTLyXDC0bCrKnulaiY2PARV
5vtPVIKgYwC1NfTPPwRhEPiQ59UYqLfeZdz3aCPJ/0ezLZ2AZ/p3eEDj/fjFMXus
bQIU7oawu/PytlhhiTrtXWyCtGM94b6Sfn5GGmLCZS2hcDZfAgtwrpQqIS4OcrdI
KrrxaksFgCSHkQXni6wlnK+xwYNqeMEP+zUUHQpxDL62/ZpFyYzGg8ah0X2o3ARx
BjyNVE8nKTGen2OqWhzZGlc7ZVEmB6Pj214EeELsZ+lSmxj82FRq+YgNiKrC63HN
ykE11+eoBWEMgf+dMKelJX/oKj7j08hHFafTf7BgiWUU43xpIe8JRHoJ+Cwb5hI4
vfdAzilZN7DcxInmvwmERNwRJFXxeGwSbWtrkNFUlzvWgO2YBDLqJ0TC0C4F0ILf
YUokdVvhNervxRbODiL8YCpRVjsIKJ2EMCWwNciFADO24EIzsd+fBDy1LEjxx2ov
ozZkwYK3TvB3NpuKuL/G6tET4EI9G9hF1mY95irlSdzAJLs6AbpIeNcoRSeTybg1
PaDu+HtOsmktWVbApC6dS2+N0XTz/svqWL8uzaHCctqYeT4z2jZb10B44NvSK0vz
uvxkjm7gVwCH2xe2oBsR371YkjEGNsWTWC31IplgTnmhLZtDWpTG98tqU2KfA8ma
B6jUHQmckreQVqOlp/v2JUg/MsEYgm9J/fADYZjxmNDSC2TP54gVlPI5iEWUx76j
QULo9WYy2ghhwPNy+/y+xXgmvYxDKNx5oJOq+VPZXGdPDdTThkq8p6PhL32wetzB
00jYgb4fkLD1EN3DvhIFHDh3Q/fwAakxPdjyP+JU8wcmsA9Yln+b7yfTjLzQwtQ7
xZPn0SRgaY1oTlepQnccbXOJG0GPCPNvitQXV59ZWi3gEEHMdpS6u87nTzTG4uKM
bUq/SDdftSc0n+wAyXCftmUtnYNlaXQwLKucez1DbMhQg9qEqUldJ95RTKqLXMyA
0QbMu5m9e4EKDvaetCIy+/smz00VTxlCwjc84w9fn5man30A5dpvEW53MweXArlY
z7N8FPotg1u0niBzKLDjWPm/atL8SRNeZvhR0u0/e9ovP+e3DOKPT+Ag1wBAm9L7
p5Dlrd/Z5WCbezbOncQEqX/650V0PpKC4KtiSflqw3UB+bxzVrOHZwvZ7SAdJoRF
vms38D3C19m8Fr5alhqZHZ5XOaZd8oqLeZucVzzcbU6ENIo+GPs9rIrKHLn5QI1T
ih6zz1tIACgFSmBoL3w99S3bv9vHFRF74GjUtFeFc/kSyVLJpp++PWrN3KtkhjMJ
oOTTQi4wBibjgDs/fs+HjpjMSHym2vkTxvJd5jun28Iso298crMVPpa3H6apoIe9
/f83ZPZyEXgwj24BC1UhVjCjD2T53nA85J1u7hx/NNpp21CkVPsBapBPHxOpUh4m
FmnK9OKY3mOXjFTEuvtZp2MJwPxWxCobtkjbsiFipKS15IXZynUMEuvUPk7ZaW4q
6UbCNdphm8vxjxyVQ+eYI8IBq9UmqoORLbqOgec/aZRn/ykQDoRio6IEFLsikcgX
F3+B0gxSEoK/Bb9VSKejNHJhbvGmMOZi8kcOMKWzUYTcQhRGsU6bEbEUkF/XnDz5
ZdahBTrpP0DVUWNPUnfuX9AS44xNCMsTF7IEPretDhqm04TiI0I+YIg41ClHtXOf
CxaNhk3dQIHJmV3LAgLQLoI0hW7MvMqQils8UlZQJUX2npICbW3xF2Mp3AEmBC06
FqqC/e0r1bo3Jw11Em5qrqyKxNK5bmC7M8lBC9Sy3kvvokk2rY0hIIlwWgYDhcyf
GfvWKMS44yB5a4WrqAhc7OmRNHqvjHtvsJorO7FUzysVIqg3/BObxd92Td47EfRY
q0yNVd55LAG/EWQNRmauSFLC0Fb5cO3rH4ut2ZpiApLyLCdtIIgKrQ5wwuXsdsey
jPvSdAp8OfzD+PB+uWRWMNglZPgSn6LdWkRi9MNPSPuxqi2tLl0Uc3KdiG+zao7y
Mht4/E7fvqBVexJEMU3mUMvX1SUeZUiAQWTg1ZBKtJIZFJM4UI4bRp6D4dtEi4p5
s1Fj4n3G5M2OCBv9bp6p+YYSvq3qAChMjLk9ApmPKPc9x5woZFr/kegMnBc7v2Hp
PuLZxwFffMrkWELyQYc+ONQ4NxZv4QWilMBwLiI7zLI4uznvC09g2hPGayFAe/aW
4KyhPy3lYuW3gPwt54OKG/uxWP+yjhOCR1iidZQVflJG73lGyo16MeGTB2uTgPlH
24utQ9buq0nrTtpwP6zVZ7ElUPIjQhDlD4yrGjREJKwAyrWzHgDyRy+mWKV5vEkn
56YlluR8qVHeFQNaWY5CzHiMJ2EqTtRMK9kIo3aFO7WGMBiJzA53M3NgSS7dbWAL
jOFWMsi7qQvYmiD3QHIN1qZq69lVj1vubDbYyCPewRdLEC/LLt/Khl9WDn+LEAzB
q3YFjje8srruo8NCWdgR6nTQhiUSFQ23rLtbycWJI0dDK4FaJ4c58HGO0iB+O9Kg
buwPZBkNu8BtGt1w6IC7tLrvN1Z7l9qLQtasIQGrVQvApsIgNo067DE/3LF7MwJr
PDNYZevPYDG5QFdJ+lpQ+rLMg8IqGQpd+2RF+PHAbxJZfdjJ2tQI0OjTUruLuCIo
BnRf+OPqxX51n+m5gv/432C2Vbi8RINU2KYiDGe4Wa6Br13nrhX+gqqLXOXw1yzG
WeLEjbx/5sItS8EqtPUeDmkHgdjtz/bp+bS3DIoYbkzDiU0JFP8OMnZfwKXKQbjq
XhZx8kGVkcINy3+94vVlKwhhCssK84O/W1EFr4ltfERLjZBIOgEhERs8YDNH2nQq
jDmeQx3Gt5nQ7+IUd4xlATWPU0nmmtqWxVVDzWfQgCtWD9/a0NwzQE51FrNn8pC8
xahf+HvkkzcszFKoGReM30PjeZkH5SOCfxkC3XRpWhMvoRjjF01O0rKxv3naCPPh
ltliv0TvQ/4ApWUmtnINmLjxR5xh04ljD3dsTczsFaOVmI38AR/atu0uybZSEjLA
DucEHaHJaWv3+yfV/o8tiK+MjfJLpVGySaI0RCtHeURAZ4YL+8AO0pRtUpcOB07u
kO3OvOMIZSv+jcxpkaf35UXPXLAsBCX1Re97l4o+wDEey7Iq3IEYEQoBYRqLGCIO
oy8g73AfWX6DMFC5bFSpCQTvWRtffZK4NS+RvOqj6fP80bRjTA9pubtWhgP2CG23
UGXUxopdlytQPTiJpb6jj/aMnY5yuVXh/EKEdtSII28R8xLOJTxrXjZxoer8z3z+
koJ8xDcw2CJkZ6dImVfj/0n1Uos/fNh7ZNorIrzw41VCUvxR/aAytDiemayjX79g
FQlgbGnd1jN7Z+DR3WJUAf+zqchmgFG/oNvjCn11uxpizCWl+N4v4b4/ECxe7vHr
gI/83Z1pQo+7DBCEPAB7h/dbMcF28/829Kurg5uoMT8qfVPTabIMcaJKhAW/fCua
GuYl59ju+Zea+rKZW1nPxucgXZLyuLAQPf0azXVAmrnWEKsfMEwq2Iyj60lUV0zs
+7pQWx8S1EmGpD3iPoir736njiJ+YU0QY5qrrPwybmz4mDAhZ+serPXicRQGH4yF
1Sq06OOpjYUrUz4usCxMFWVi7ZKfY/Xvo5+S6CYvSGWNXsnsbvtiQnBGz01KSjkg
DVhPSdW7ooIC8WgrOOEKiCxaRsbS3jV66kJvDfcWvHE0oZCpzGLdjA7tka2awbq8
HD9qm2GMxlhDQIb9PwZLt4zIKp+i1p1UoLZ8S/sNPce5DeWMx2gfQOWwCiI6KgDv
9aANDx2exfMGiNIRVaqVsHDLDEhjEXwnGOJYxhUQ54MEed0rQGdV8CNqmXU8oRG5
s8hv/AdeuOJ9neH3pUZdB9GAd2cSi9401srkkNqahr/Jk3r9LIwueZmNH63S2Lz5
ReQ4Ymu26f1BDKyTQscX/zwS/Dp+us7MT+DP0jZIaxqYAdtEzuFGnODazGEa9Kai
SZAejaRm1SaUNFWAipCtA4GyVtOTIuE+dvwF4TWcy/yXp7/epMzJ9+9KvkJmrzFJ
qMJLBOUvNRpzXKD7NBxx80d7WpS8UuafRKr4hNWksaC1b0L+xmfwX1AHM4xe7j0X
7YNwK98PY7BtzDj1tDFWHL9qB/iXDzKRqChCW9jCkjy+tS4GA4jJLZQegQvwU+5X
BmFvKLbSTs6pFhoNru6vMUCQxn+UmFDeJuBGsrJ75dImfEZ7JqDq16q95zXuPzw9
NTafLMlgbivbhXnW9kuM5VQNf3zFhvZ/rHK6UENGxecP2PISQaQZn30rZOdKJ3xQ
VlFp+eOkH6jHYmoUje7D/t5HalkoaOM1LuQbxZUbi3V78EiSOswh0nnW7y7H7u9h
HmTi3YV7NBKEclFdNdJOrm02MU9lOISCRSMRIzJoItXEsta1F3vMzBqntso4jWYC
nV8JXvVIbt32nfPibYgEYSmYLFwEN3BRmp3fF709NmfXMcjc5HSrvyLHvOMw5+gO
JjacTkjvXJp0+fgA/v5CWM51ik3tYCw3SJgI64KjQ7ZCRKvuD0vH6ZSfSaIh2hFl
oCraAC99Xtr+wKkiMR6/4ZhjNMVw7ZbxvdHDaXzjC2uMeSsBwmBpeNoZJJYHHtkV
2w1Ju8Nsi4ADtEXDNPAagHn+/GZg2JuPLd3BZrLw90S8Z3/8YTU9LV3q5EbqVuvf
uMQ/YUIZX3hkMPzKncXNXxgIAGLClkXT89o8wHElmvGIXVuTA9dskdlCADQEmG/R
n3T1USICWsGEMlHrIMN+QrkPRQZ83SXig/XytPKyNvK1D3qfCiv3hJmljzamVvyu
GuCJudK3ZkUkXEe/o/iEJGJrAdsOt6HlC7mikDtC8FGqW2V0yVbGP+aVhSlD9s6g
eFItE+jzMxyRsbT+FG+FFnNnt8W1R8mvLwzgh1C83qi1ARV1SsQPgHJt+glUOwm4
ghefqfifED14coBXqpHUXIY8LxUwe8YIrcpjaTYEmsS4Rn2f1RlykOPNVtM54jl0
QWvqIRezk8ZT0UNZBulYw7ho0BkHgCaznbzX8P2vYUKUU9+Ew+bOCn80Z8dRPk6H
bY0/yXEA3gSKLINg1gLzyZ4NRryX0cXzCnxtTtoJHlojtx84yoxz7Yy4vH8wUbWs
djOGqfNxOHX/fqlte/YnUT25BpIFgBeUiDokJOtf1NE2TEvVmRVXtt9cxCJqwfo5
uUR+DHn6tDhFdLR1WzbQlzf78XiwI0Wt44PlAZfgvUVkqN/HBORotcKYeEdq9X6L
1XANUeNy0js/Ojwg+hE8EAQOVgSccMSUUhNhsZxNCkaupYp3bhtpZHSM2ybpa3YS
bP1PlOOvCfjz01GLadeQIA6iJGHVTJKqtaJm3MUHG5Qjt5kmgMb8GiOFjyY/YkH8
TTvPmgatYygYtxyw0dPDGVfkjYJhO5vrI5hnZqJFWiak1MKCUkFs5GNZqyiVIoTJ
oakH636ZzDOLkuJH8TLoyXfihyJjxAM/NTw4nFcFDDgFM3JNNlXknH7ycel5Ul0V
9zxzNWERu7yD1EZvPVNtFs1fjiE0h1mr5EGhLQcUO1lpRWYTdQRidZIb89cIw5rg
keSzGlmq3eX9OrLdZ7kF19Qc8bIBsoASZE7hqWR1IDG+trKy4ZsyUE2QhudjZMfm
psgGGEm9dRh8vvk8nyoBGZz3wH17hw5MPZyBSRbvoaCW2emuZVMMh+AShUDVKBRL
6dAdf3SXGRfJhDoBGYQDo3n8QdQvd+fdlQtUXPg6tYI5vkLxFgxbMd3CHBNTUZLL
7yaT7MiNgTzu4FW1uLRoxRX7gDZknU4S6Hu5X4/pijn5e7WyfYXHqrGSywfJurCY
FGkiVIgmhn0c0YCICrP8NPehxaW2Rf/w/EVO5NqD3r+4YfLLBSyDykBYfFRd+KMj
CWqPF9zoktnVvAMI86MZqmCWJhol1fNuufu1m+2n2iJxhojaoNvZTfl5e3+WS366
qHQfndqJlyzbQVSJsB00MTFprb9LP1nNdrGI9tg6La1RwZlKbB8/cEMzaanvThAE
7dXKBtAh3oZe1XKLq2n8eLpKpK3ybXKFZW/2CK3zs2EhL7s61QYDSfistZmz2GaJ
A5097Uoz2jV2akzinmsIOjYHMig56R8UA7Frly9RZ1BLFf8QZHUhQUfGMsOfD0y7
NEy8gKzEiN+G4uo9m7JJlq2KSRlL9QB/XJlxMq15v07FC04y4hcp8ntCe3BSGmGG
nEe9MSo1b4lIjqW3VPpFek/Y7Xj1nduYxO5hG6jD21S8Syeke6TmXJ/gbOXiUsPw
IvXI8mbzDA6B8rvUTHa3aGygbTF7s7+Ig5OYAR4mqrucIbv5RlX7da80Kjk+cY8X
MJ0w6VbOLfu3rxUxqpyIzQCsUT2HuqMj0dc/KtWmKntvb4HtD1rRXlUSt7CTn5Vr
qFoJk0Ivz9RH/3Z9YJSsbjAinzVhMtWiTgtsvTibI14TYkpUxK3zgIYmqRvAVUyk
8vyCLAsTnUsaoDsUUxxAtiEyP9YyDk9RxuDtehRfyPhg3aUJ9ayciE0AoI3Hg+8b
tLYQYiATR3KxMkUSrBcKgOfaOr2pMLDLLqlU2n9WWAXnlMaQ9WSlwYELxhSUlr4S
LDUCW49Vay6jSO9+JvlUW3IGXXUQaHSFb97K65ISwbU9sB2D80W89BRHXxgRzaVx
WLbCqJ+HU9036+/F2f+j4D4xEL8w9qxqJy+aKUnzjk+KhypPBcpj/4sICfVQ32Nd
BhSdzMzL37GygztLWLHNfw5kQpvi4CkP1zxahfYjII+PO8jdwpftV/Kfp0HlxJFw
GHmef+YV1EhD+AnZASDrBAoXd19WDon+LL34dcrOL4+SY38rJaEiU27hQHoFDlvW
Guj/ADJpzZpHCGeYX8cMC437wUzzT52MmZnExBOrZtH9ZQThAv4MMPgpex1h2jbN
IkUUlQB0zz6Pc/HDKUKT4tX1je7kLqiX6oMyCnzGbsLWWZuy8+vxABSOh5e8iST/
ralzOXlxwyEU+l9eocH14vouKaCLdv36xFrnCBbwOiFF/HPFiU0Sg0yA9sPW5vZ0
cnKwjZtI7C5l2jTgS84r+8cltAVtxlo6Xa45+NPv5moHsesWk+RpqQQBF2WC2evC
5+0EIZBDMoG6Xd7nmdSP0ribknIUQXN/fJTKakQiF6GNllJTQRDl+151IixjbyOd
ouNhZ6KYosqXgkDpytGQYPFG0E85D6VEQ5ETArN7gxAtbkyH5UBbyKIJ5EJzfZ5n
om+dfkj2Wl87Mny11GQQ4Q+1sUGZDgM/pZWZlA66bknSZLgaemhqIir8VoxA1rZz
hzKuDj4xb+DRFrBA1On1b3cU74Ly8+3fpoVAIy5qBv2jodEV+CT8ra0yTPljxnCS
pUl35a2wX+9KFINwbX6d3JVmkIra8iIp+9zysEzrZ67kLLgOrt5SMI987rmHA3PG
5NtcnaevYY/nzIKb4oB+LC9PsBTo6x6nkgJ5uhByHJpGINrfJTsef0FjbkRDLZ7W
Lu/jPJDOTGWzLGqxVBiS+X6jpFLjn2Y0oyvJeD4KhkRXsFjPph0aV3id61pXYy4N
jXyUlUj+dLzQA7/xB80XnT+h3Nw4j3MD8RtOlJwRAHYPFERCs7sM8xj3S7DgzrS4
3OXSgwZgL/0eP4nKJMln0Az5SDHiewHI9hSFiHASm08Mlmc7HXDJT3dDM8OYeBQg
mEuU6ptPoh3HktGFZppMwVhLIOiifzt2TfZvLrZTeBucben5rcEzQmO9a8RFVXXF
n/cG2v9wExxqJ/0C2zxq/rpUIH7z+UZ49rzbMympR1LboKLgke9rPNfv+J+Ri8Li
scX9zskfr4n2koi3/+Gm9IaHZDFXkiK0Ze7RYNxU/ksJdOO4z6j71ANJzC46/tKM
n6eYUXOpN+xbKlYCtJWm/iAuNZnSa87J9+QLBtTOPr8oGazV/dmv5ugayCbGhnra
ATBwdvo48PMqn7TP42P2ruUYN1HQCcgqS8XkMzu8OSI5o3VExjiFWclotAJWkYYI
u1Hjrq44R5OfUEi33AEHIBDFtC6AtgXlb2nwThuRfhu07tgPcFDDtFOyaPDipIee
D97bWhRs2fQDZTgoD70m1kC2ZEv16zICOseKuvaV3peHq36sHvfeK7SZr9cDQln7
8NxyQ80itM99byuHgc9Yofxcz9NexhowLT9eS09SnG/ePzLCO1bOL2RmEo/DkfAy
IRlCbQEzlMDKsSvi7KycPrbSORNEqnM5rWvI7FQBiD9GWfjFpvw4g28DDEa76QK/
YkfpWtgPyoB8PqvtWh50Tx5iAqAkdaAcg9dLp1BASDri9yJZNFPLAMrUifuCHxzj
Rl3VJQ4E95wA2lcTstgDGavMl95q6tTEFsDH3WNKLhvD46A8GiXWuvSuWICsivF/
9UEwT9GpAXq2Cnh4UGRGldF7dpsr3Fnk/jUAPlCi2O2/mGELDV1TpRHPk/Y531cP
gjsByky4J2OhmC0+Ludbp6asKj9yarCLfCEK3ROabgs8cwAwgjsB21RQlynhmdHe
q5xyQh8UMqephnpQiGYrIxmfOO7pbDongDcW1QbdRCVCu7E3ppXYPU4088R8HZjW
Jb18XtvRsIGPZfaXpntc2m3d0Yt8IxXzSjkSYfKzDD3MpLL0QFt1q8z/gFJmGFro
VHcak5hoMCk7MdDsPc09sdQs+fIBgZdYVZxExctjBbPKUeR4a9ORBQCMkgZ05vSX
Fir1RbqXySLTKRc56RdDsRsa9puwpaIdAVsCcoNc4ioHm3AeVidswgJbWEs7/mjA
bUOHJmWD1ICRh0iNPxGyc9uARfnc84Lgku1mnGvNkW2Q0qyAsC3S0LCNM9rCJKxt
1eHWbAXwVpJIZ9d1tf2TOkiNygS4i1igPAP2pAo3b+NPQyTKhCos+1mHSq1JpdFf
xuSoXReEB2IzJeeSy0GQ1jR06adWZ0uKWqslVWrat4r+T4J/+YsbCCNuYnhwTBMy
SEEULo1GrV1DhnSFoo/qLuD2bwomO5N6rNgAPCrIp0BtTo9KKv/zvReTK3bNc5/j
Sz+ZwB6/BI2/Vb/q8iPkq44WIrJ62K1VnwQAKcY1zaXVPEHcjseMOttXhkdtW+RD
wlt138ZKO0l6upbHBSI9zxhwFMy06TSYebNUEaDRsKdxfWxOE4PWcDrQry6QbDNN
Me7R+aKXD5Mbal/NTCIrk8T+SvAaHU03S+0VnEU2XAJcNaWlk9yD8nku89OK09mS
uD9X7KKdSdeULC7iAQP6hvxvYR+sQhjOmScRMpmTD/enC9u5PYnlgJzAZx5twuZp
tmy3jm2IvIue+Pq1hPnKap3z/Rpkhhez9h3NxqvSICJrzp8DJvsn193Tt5jH79pV
LIEKtQRP9740LjcaHhTof9y25OVvypsm73LP05i9egLSSQqKpw5e58tEPewr5DTS
FLHVdalt1aOpANLEkjrUKgILYXsZqRutWN7dfEnSu0Tl8loUVQPEsXF2VktRY7ZK
IamKO0XX+6ZenZ2nb4DB5KPFOhJ25c7ttCKvzOKqN4so4sYPPQrN62B6akil9QGG
U+azQcC4pQAWyPNxl3sWdEVh5QtPp2P7iEKZxJBcJwRFl9Hbd4pOS55X5COoWemI
Rb7PpC4cEbSfUIYBT/3E/nBi027YxWVqpe9jW7a+8a8i1uvnAxGBSmjTfvy7EM8A
iOWNl05bDrhw2Md5+fccIJjd5HClrNTFrz2jAQNbeRAVtfqCn3VhuiIV5G308dZJ
pjS+Crm4fnqq6mBb3h6ulu8aoQNJSMhdPF2yARq4ntgAS0/E6ZoXMf61mBffRF83
QRsmzifUQ/lzaeUxsSM+M/C2WjpKJIQSt2phtou+Vo5WcQs/J/B5JxFxVkdHGO8V
5GH2SnFi8VWQtflEy6n2wzsLNUNoW/4BGinNrBncsgXi3WkrM8l/yZucjxxgK6Sx
JixHcRg6GdHpgOhNXOry/P67ZqHh5SVE8t9s6hJ6EJ3bpkSwkE0+Q+9FLI1EdBvp
mOAyefuZP87zf/5LZFLWFoNbogU6pCA+1NBlTBu4oSh0H7Mkxonu9gsm1nRZPQxO
L/12ORKwETawJ8i+lsWhH0wFsER5dJmw3bgW84gQAIowyeZ/gf54IS1SX2LoAknQ
/6dll0/R4+V0xfGg4GMsk1F2fz2RHDFFdKnz5WbIYAy0WUXcZolE0Y2dRRocp3m6
LDNosRSMcvlUMUpe93mtZpMLS6efgbHsH+ZD5AByQmYqZzJ9pPY+jIiFcBSmAJEJ
F/pXGViJCn8rh2/sWd1lyomVfb0M4fQbZ0Cfv9d3mXNndHNIkcLTNU20FtHajZUj
PfZpCuqDowWeaRzmvJnPShzDBJxskCPmopP3FTTmtEVaM6VaThXI50Xi3tXdSrHI
PAa77kOTraR3gDCAAkP9VLsiOYAhg7TE3iV2PjqsFD6soGzOeT9hAg2fiDBC/zBm
eyfr6D/2ofS/JfgUgKLEzK2JwcvkowztgpOE6MQWWKqSWJpNXZiIloCV2+0r2ikO
Nc09AV5Y7zFBCCNhP1g9xIfiXIL5sIUlhP9P10ztZ3oxBhTd0Lkdlz3vrQRv83S2
WMGPT+YojmmmLo2xLT3KPJqIJz/lqFWFBa12ThW+h7J7+0GnymNvXycFl1sIm0CC
YgAWrQgxVFEEaMzZ53mLL6akr2ahoGSv86+PyZxIiW/1NR44PvZrOLpc6nhclucZ
/ZV1IwPLvA0czKrSapCy+mlDSorJGZQRkJ8b/juPgNRemD3/JcrcWXI/qhwhgE3J
tEVmYOUwsYYhKDmofX1MqyQMC1ESuvRYsoRMrbgbVd1qqF5/vgSLzlb7i1YL6Oe9
UB66dgTU/mhPut4wF0odBcndFwfZe0xv/sbiD1n5CbBP0lwLSKK8UpvebxeIXlqn
CZ/LdqVW8OihcjcH2BouEbHN/TKdm1oLN/j43MuBKOObH/qTU3Kh6cVQ+3gTXGb7
TYyrVlU1lXVcqdhlCWdvJ+fPgIezYHyZ0BENwEkg7bu+vksejp8pA8AwDy4BPDrG
ixBHmCqOILLPwfdNrIpVbqpkPw5RJ4s+VjYgPiM0HnTTgc2nyAcTuVUCHBqNQhNw
2YOri8CEsx5Z1nGSARPBdBCSwhd6Dp14s1MB7dB3ghvFHmouE1Ot7osJgSf8Xo7F
z1pAkfSw5E/mU98u4t4tq4dHKmQfuJ1gaWaTG4eyaiOvOGxa21qQct4DkuKUCeYl
7MsrfSOrTKEKGv+WQpRLPXskP0AeutCMr+SEl6/7K/8vlyBTGiWc9lLV+q8vW0+T
qD/xEMQtI9LjIvBKNj2ECqwbc/5ldGNC6LW9MS2Ma+NVU77EJh8U/ionryaLLKSQ
2fmR1CzXfJSeD4QlCKfNZ4YxA1s+OnT39tO4FNkTcfku427H2u98GZjQ8kvUT/fy
8AQoM84/17udRyo7V2vWyhseLxnILrNP4Zk8VxjMgMwQ8AadYRv9Ppd8MV9ADtHJ
WLio8FPiZYImubk5WXWiV/BoGhBDVIde/R9nSHdmVTu+xSC1hIYth9i+4T0WbW1e
Uq0X3nmhh5PLfKZxYP8m2/oUobpdwmcsb7IPFiyHa0JbccOEQDx7XTEQXoQLfPDB
BmgCT9R2hWBQ+4FFToQnON5UsAzUAqvuacUjYj5CtwgRj/s2Ap6CHOD1GeKPLb7j
vco9lra26BcyjQ6gFZOZG9IR6s9Nbj+6yrZH6EAxyrpItFBjQeoYlIhbYl5wDNrC
jJVR3N165ajbkU1SqKDAfnpN/dqVyiCS+eLh6fpo/w/ZSaemd+CgrpXkcymqnJ82
9bDJMeXPLDl6RZ+wnJzLYoLsMViKyhHJo5OxXT+tLhj1cOWRNo4u6ErqsNXqMeuo
SLtwUCYQ7KuGYNCYpKslh5XKexVOzwGaET/UfDA5kyGLz6dMZaUNDf4YuXrBVj2V
QzqHTLgdJFrVri96FEC8vEAPkla2+idgT2ybQn/Eybk2d+DdhiA/IeGzIFUI0uKN
tYXHv7p0aMQHBpBTn3IFeJbZNYR8ISF1mZdT3Dwz0Ow7OUlzAv1OAjpDOLo2v308
lhklMuEAttYR+60MMjzsET0KVxlXjBsv3i+Clbg04V0S+Ri6jh5kwW/h1pV6VgLD
cWU6GUYgX8VVemkTtqmBl7D/W/W3l6R7IOYduBqEqGovDVjk/YsHfpL4AC1mq3aa
A2yCkCe+ZhFCZqB1ltRZXrXDfxIrFk0a9cAdoH9Gm1EmNrdPqPRb10jz9PvScUM5
54s+gXH/AQjZcWcdwoArwjTmuqkvq+Xfl1mCcKGQ7amkoLJbNl0Blcf1LfSBnMat
GLE9YiWnPDuFzwvLApFm8EsoSTLjox0BorwXlPRp2wZGyObt8DBAU5ausTn+w9SY
EfDcL6NGm820we706HzduH3IzI37sJioKqUPd/XHUcH3Fp8YdhTO1+soY4/oH6nH
Hk+/vxEkIwF8cYpyql0TGqDxBbYzid1z0RKI38ttV9sWS9JvN2LvKxccYtRcZSFf
D+O0RGvbVODDiZq05pzVUXbykXwQcSA3ZcFKdxC80iSzcV1E9evSKludDKmBrc9g
eQ+OpFuo+trQ4/T1V9de0rVOXW3ItUbpFsG4b7uIqW4+U3t+y8hBf9F9sV6ds3Fm
g3OHqANX5H/N3IDgfLCytnvoKKkqgX+hweEV6K5qxXTojzSVzV1X1U79gLYUy3DT
UokainyvyIbt0axmDGGr/PUfTkaaSMyWtpJE7/F64QBG2/hnlUdQhHQXLAmjzhiJ
UGoHA0Pb5A0oaPFI+D/zAaA8wXwH6Bi77r0pLdMxZMzc/FEq62x3KabW4f2o6wB0
TeqqdOoACVwqqnWpfvGDJr3xKRSg14F7eNiPaZgk72mWJFmdS/w3wfAJklXSEg6B
yr/Tdl/n0pkX7/Kkc29QszqjFBau+ULKTpKI7Xd2PwzfSvbyF3Fr5mgDJseTMItw
HO6p14dEAZ/L3n6/ha0hSJiaDEqzpdxFBN7+302PMeKwC29YjBYGaQyNhZNqnxCo
ac9ZxQhXkuzFxWOrJwDPNZUvS6ljn/xck/iyS5R6cgDWFIrsL0Wo7lxe2lsHY0q6
uWRRhYhbrxFBLuxXsCXoxgVUw+K6BxcEI/Lgq/VEtE2wa4ALn3VvhardwlaHoiYe
7fB2ftZPebT9kuDp6uN+aA2gFCBKOcdanXavZIV6OIaLURueTnYPUrQQmq93MLGv
sB9M0f64n+VYAhTVQV/HC9vZ799WEtrckXRQoLy4epL3eDSV6tRIko4mcaAEggjv
5HHJnZZfWTfjB2f+JcKp2O5bu3jx7CViLrktNembML2gJINsL/mUZrfJiqKuxz6x
k5elL1U7OEFAlh/VrdxeMGxAAkewq8hEtWJaYVbATdZmgbtYsO4OqcEFlXDVE7j3
xgJkVhp0kmTvmasdjzLucVusL1+QuaC6k0V9JoR97PX4jBNmTgcHDQ4Z2yKjGxqm
0Mgd/iDPeze5M24LPHxtNIKqMkrDcHeG2KpztlmHE0EjaelBBLBggadiPf+kczD7
6azsOwaB/4RObYlk/du/I28n8GTyqJ/pjatPBoBM/ffe9BsQWusQnfLthDhVuIOL
CST45cBfmof2g8dW3VqSo8ZqAYHJsjoQnm2H/a3+TxQIxY8DMaDYIcb/eun+7viR
akOyG7VtUh7x8jdxtlPs8hixLeYwHHNh93TXWfYE9Qf4LRFFTtGAkbaheqzhYKU8
wIMrrJTRnFkzxoPxyJ+huqOkKUevv8/BLQ6Ntv9ipzjofbLPoil4mLRXML7LkymW
O0nVJH+ycXKb4CaXtTShe4I+lvgqIOxRBBYt//xjlmZxT30nMChJQZ9tfAeCfOlZ
H/OYukXFt9Rv4TvtWr+5tb6hwGzqiDJPAyTfzSqMBUoShvoQJfNhkzEWFFbnAo55
gNs1K49K9UhTjWJwQyECHMhzuIWVRNR+Ec67Zd3ef+migTvuO9sZIGHiB81swzk2
qznFKYvX0uV8RqZjCnyWoKBZFNPOK40H6XtlbGKQqdV+40YbxulmPDEd7KCyDPbJ
BQfrISPhRgX7Q6FvhHrG5UVEamVCwzcsVBxOrU4t/74CtR2hsi07BHHnRg/GgrS1
oyJym4siJ69wvLuL0MQ+LaXeAssSGjrmn/PGlhPpCKcq+oX191oP7sV96qQ0B47T
Cdbnw0RRbKOabBKmJUNdbJhH3RcoWStKKyE1b+UwpG0Op2MmtE4/y8xskycX7VqF
9Dtl2nXLFdqsgdMT8MXrxJHVqZMeYSkLisApzSXH9hEAeeAq0nnbgcfr0vAvS8JX
POIl6NHpFzyCjIXSmEMI17vdE1WiAhFVLTBO4U+81KbAJTALpfPf8vI4Q01es3V5
ZRO9dZ8/vXm8+TAw7RNkR2Hl/o3CH254wPJTNrUKPIFqWGd49zUquk9dh2/TgTVf
W0GHTPru7/SCK32kT6z8jLNyz4i22lKi0vW7f9gSeJ4RFTIATWvd+ml/pnAr6zPd
WIRCvpkfAw+uYU6/m/bJ+kJucoEhznN3CS5Keg3WuIDCSwckY+l2mvUfbgXj/D6N
IBmcj+Ie81v/eN/Pa/gNsp7VFoohLjYCI44iAfQlnd4qefRhrBX1om/ct0AcSrM+
yfVAC4AuR94wt2p6V372JOoQzFMdEH/8UaO4dKF9bxn3NYgUiy5gzAP3fNk7hWiM
EOCCLEls0ZSN5fIN5mqME0jyC6475eS8EimMA+x28kiim1894v62O3hQqxWYjWQW
UDwE7OhQEIsHUIsjHdmuOAnIf2T0oJk6CSzo9KE4rSVhqGINQNlIz1UQSJ2PJ1bd
4ntNVlqActK86P4urCFbX8dXsv20P+mRvONkjqEvbj4DYA6PpeOfuQMWUTt//8Jn
QRVP8jwP5x4j+QPmvxGh1bYkMizi/nNGe0G79IOFCTgc7h4Q2l7reWqnceJ77v04
E0aK6nHGaaFEHxdfdorKb3hpeQRczsK7vSEiQxrkQ8hLWwY5QOzN6GTsVnZLqay6
2jkpPKocwQY+Up/xBXdoChZ0b5lBUe6h9ZpCQoN85/97v8aOFCNIBoIOL7cHgYIB
cSRvowRQpALLuFLyOL8ltwx/rQMMPahjonggdV7l7wJoZmGGD8tyvD5aLv5s9erc
WjUIb8BlRGp/hRdhkkc5YNOMxBEURJxfCf7SVJFQCHYNZA8SlE/Z4bRAZxGNyz5N
DnvhUA4zTDjhYQa4bOrqul2P/l4B9zUZSyac4DXG4iU1nDP8bIgl3+RBu/6qG8Q2
vNdAw9h5D46LWEzpMP1rxA92zjZAhBtb6KGqmbYWuRVxJeHmVMbAVV4IkJKVQYhz
8ymI+hyW+JoHl3AWwUP161+qQ5xoSaXW4Yt6N7qmZpszQwqCkfWujwezmUX9Jeoa
crzs97BM6y1iaHfMQ8kqDs8HCDmwxUUq15h9bJgUnTKm63rtrblGeUahhQJRFGag
+GyOXtKEkIgQALDKlcT9IE2ceZy+DKX/5hDgqIqaz9+5SLRfcH6S87s+Vwn22NkR
2EOdUanA+1NhTjTe2YVe506g4epqdXOeDQLJA2VU982dQR6p0H8cIzTdArW0Cfpv
t+0pZjNvMud0Vv2OkJRwrugJUYblc5KaetdYQFcAsDXAuPjAUehxZWwwi30o5B6g
ghmTc2I7G4yv6PJgzunod5616ffZJPZZMhWX5Zw48R++MHIfWdKRwp0iN3psEr1G
W6GnFItMgZphXUqHb+jN49TBWghs30FiM9glOTDm8vnWXwT94B++IbX0pQKy4SY9
uXytXA3Kf8ieRZRrXhVZOtmxmkmqz8EmnFB6+sR/Gp5BQ7lAVu676bxuq4ZXqf6k
p5/H/K8lUYxWcnYbQB+H9fi/Hi/ag7aM1beUeGZcF4WDcIMvS7Dc45kIK/e/SjA+
YY0VuiRlJ1EBb7VbeJ2ImLyDedLy02EOlPvasQdPArEjC3aP1+I0qp4lBY2K3Wvf
XjqctLeGESTxD26HVwzvjfOKPLS+rhdDicalEaGftlPOKamR3Dl7qRt78ihjQq0e
A5bJmhTAOULV59jvlio0h4f3vocfywHoTcAImmDN5YelFyGS7+u7eNzZsZe9EWkw
rWF10eGNNgoCos84JeDJ+GNixoLUT7nxe0qFT/lrAdwEMuOXyz9iMx+6kdjL9LLF
iylD3FBMh9yyzJJPTETOouml4YQsXE5JuTbeCREs58dt3aSFPcAA7rCmHtkeLQFX
hQuJXYMz1G5wZVE4kGd89H7wjxUf1gaFTggoYDnN4PTh+SamC1E3ez1Md/LPzCBH
MTG3/YGDaYS/Lq0d74rR1boIJB8PI+pdnnP7XlfMxxfk9x2WGqbtNDWIFHhN+qXL
mKz+58xoYUJnSLeMYgkq/d8doygtnh9wi7ARjBAkyF1Ud8t4S1zl1zz6YQQ9kxYU
w+KhIHJAXgAIB8/68EaqVBB4UM7EcVoFlrG6CRheCy+oZPzfAy0mC7kNAOzHVHO1
KmpjLbAFrY7xfBj11VhSFv+APY3x5eJjiyDezOli31NioHIwQpzdNazkP/QBjcON
Pa7vSG2rpZJTQsp6E4EW7/PhvTihB0f9FefrOmB81YZtnesUkVVV6cs30G+kLEdF
2QekUbfJP8mXca1a9ecQkV+cnOhEjSyWX+wBS6088WBOSiud03sQuz588RPST9O0
qpcKEbxsfjmUnaDyriXmPnUi4tuGZhJ/OwPwnDPBN72xZ/h+oiJoBAYH4T0LchzG
GYY7eatOm4qdG/Tun2MSZzxPUIf+YpPrsAk3pARLblsIx67iLRbTj28cJM2zwYmx
lQKMG05Lca1vtB3F4gCavZ6peJ5s/725nC9O1HoYNten0BKe/5EBWeHOOxN4+RTh
0cFyCsIdEJSENqI/rNS6M02GrJUJ3gajCxOJGKc4UYLaFsick2glOHLoUUifXaYj
f0WiqQgTDCg7xuevDK49mvUT7p6cBEVIlq0sgIMamC4Ovq2b43tG9gzV/6NcgkIG
88GFuslZFDzKInjXgOzBDlOftCQhgxIoKsQnVoGHtr3sck+odgpcxBviAxmFJ/8B
eo35Da22SFxkTx3Lg8d32z5t5rT8h+uDV1dp9kHij5kpsfXOEfhKIki75RSkRTdB
a1j0ILegzmdEtjnG30e7Ib0/ZdJMjkaixrx9TgkR/cbXP/1S6kthTBllvmiNJY2i
nQm1rXxyxbWncSnA8YZPDf8NjJT0WPeFKYtHASfcAswVQsjd4yXKijfhQesiuGad
zdnWG8aww57CosKk4eVFmSS5wTZlKPgPDwWGA7YDUtgZUfFmIyPYW+sRaq6jrB6f
rl5foiII/HKMLJAS94wHgAxIfFyL8tV79MMj2mgJ420oa4oZ5MX+7Jwxtty7qxry
m+aC+0STTtEBDW5Lsak5LPSzJDXvoJhVZzYZPRDeh08Qe2dRjVjRuVr31NLgOv6V
GKy6pPEjGF2mPsHlfcIiD67bn9iWW60DNpWzuy8VJiJcPsmtXs01FvbFLirvoxIU
eGVMhoPfAt1Ff4DJcPC05qWm+GZKuzuMN914HJOYSQPgPzNC10v9uckL2+0+u1h3
FSEx4ybH7O+09zefPvKWxulHahD4mCVrIWdtJsjHIuSktBvyIMkpLu5vpRan1KA8
1CDE71YE/Jf4mszXIJmwcJoCDUHXQhxql/x2gmhegZ5qBB68nJoZiGHdt7o1EvEq
ZNQiL0GUjlLnOZv99YH39ZIfm9SvKO4QFuC+IMCcQiXRcuTblfMrBrKKAXHaxv/H
VVmnOwCfmhSntw9GxTGL9APVcn6UbzaJzyYa1ks++QPCuEPMD+LVQsAtYYQioaQh
GW9DWotqTbR3dG9/YwwcJmcUf4UJcxEdxhxX2z2o7xNErIDa5y3j734yEh/87ZFW
LxjJ7ilhpu8QGVwXCb+ePnDQPUUuvYBtD+peOvCILxetn+wAZWbyA3m11R9UapfL
YTzz445DGsJ5TJNK7gvK07IAqd/TmqaSzmSxi39h2VNpIx12lnOKzhlJgkg6K1wn
fFiaTvPKCzjwEG5V4a0zvOVWPhkE7Hr2N+01d9u34S+e9+18zSeEomlp+emFdMY+
Lx/o8mZzK9Y/v+5//QI0GAVxsNmWddKW+zRmOOX+OSu+SbuTQRZq2AiutEym0qRp
SJw6UP/7GGFoKZRH1dg2L1O4wL/ekL8hafGJLwP+5f+8vRJqRbO800g2jcy/34/C
UC0z3F6HHxAUT1jj8r2/OCeNQ3slUomoJ4Ma6BiMNbRZReJMVh3XcHKXpeWZf/8Y
DkhLQ0qcsHp2BriqpNiXT9lweyf5MzX/jZBKhZXaT6+3gQU2pB8yDKk/dlSApxhT
ck6baJEeIbCXCTHA+7rQm1iUqIABxQ8IMLN7oznHWRz+fyihjy5ur+252g+js0Pk
6d5f5Cij+om9aiwIX8L9CioiPM8M8JxcWiwoM2c0hgAmL+IptV1bQEN0BOarEK2q
mOemlxHluXzd76psqfXSNSnxgHt8LqFnCepIp5cWl3Y9ey7ruwKbZfYkeqRvNwQE
E8D33mmTV5BHdRT548wzc4Uy85cF3d3eDkQ81eCmCnXel330xJa9Udl+ptdfdhOz
8a+RKKCYP+gPYVyJ3i//Uv4QCD2BbGutAxtYBjMZFli/Fx9+J6a2I3PU/0qp5Wwt
n1PCyQ8fq4xgLQXRuuqXe0pSeGOXZxqtee/u8azJTA4k7qZtjrB7H+q9qem9j6KX
X5xcSwtnUaTz2ToNu7HmNmBZE0w22qxZyRVk5izCvlAb/4qw6Dj52zMuAHFSIcgM
7QZ3OvAMJt7BtTOChgL0BkCkyEWq2hmangbOPDC+Wz40ke9x4Obuxgyn4KzSmQHB
dLKHffcza2FYQyGSWLpOFRP6osJDuCo+1PHEaT/P91FO+rRvDg8IZRYN2qSMot37
BMy9Nbo9VKrDNDGMfN6G3NrsXPSUdqberaznHrSLMQtFi+EhjrHE7ou1yhxlgqWF
pr7bVBML2AmdikY3nHGtX+2WaN/63n3n3VPcA1YRuztJI3KIK/QRf9ogaFO1hYdw
UuMQCiDmPTpi6AbX2Qay/yQ/twyU4zX9lrbgNDBIpV2yBnRj2CN4Jp/UA1at16uR
/+KIBufmwl3alBbrHMOOuAJSZxyNXEqSpjNrjCPrBpf7Ne0DZjxsVLK0/byoGOm0
Wjb19rgtr1P1HmcR6DSOtOKO9d4tCsZvjIGkslR31xTLgMC99shV6pKRSu/k0vSp
C0JPVrOdMsgkf/J0/b1z1dQVPw2hqKU3F8rYyXYRlFUWRgZEc3ZOd6gYWGlJvGWa
fM+kSCgNWkXoAR/jvuA8i8mocselz4iP7YYiwKPeMnvZgznirn4Q9M4gH5EZ7Tgq
yYzu7vxw8w+GBMXw2El7j7hV4qipBfG0Y/wLlA35ox3DD5yUGrPHfQr7iWNr90S+
yT8/FONpPn61WcZZtCpTny6qOqJnWrlG2ROIU75izY5f3YkhFCeYe+UzTMtL5n+U
Xbclm9OeHJjtSkUDamTW2r7YRy595W/zhjqu/ZE/7Cy/6bW6+1YyQaL7sTeFYP0h
7fZcaqD8iiEr1GdxI0z0j9sxnbPyf4HCGI5o/K+2aitovv4jmY8iYnc0+0VEfPBq
wNZGjQd8NHD44ICLExZvgUVZqg1el4Cgx+yvpGiiGmxZnlffZhSNLULUPqRms5Dz
w0tjADzMVJPibO4AEWry7XDrWld3sMWS2aKbXevoq0i2LEaIsex6wvsSLkBaO4ZW
OXboU8UNp3YIdN9UAC5uNHLyWsuuHnlQj9vR+zUx8g32OHKOVevWjnoBilK4bPYo
BdLWrBQRhYEUaQ+vXPgdZ1dzL96FnTF+UEU1iXFu/GRrH+p33WaXJTVffVRSxn1P
ErHHEoFu2cH8h1JJ5hU+lh4zNswflRlNsxcS/kviSo/aFNXYCL69RJgMx2DnNS36
2VpkQaYV7Vxg7QRxgfDdSk5vaUsYw+S6HU7Dm+wl7N8AtftWS/c+/+C+iCnt/rcs
cE0TkLXTZWHGjko7t7upFryoEvah4L74vhf8lqG7Q+NFxzkufLfuNRdCzLRQX4uA
qhLYpynT4KKmiG/DWtCGQv9ybJdKZmWULYNsz7/B7PvP0rmiT202ph0JuSfelbmM
XLAR5MhMEMhhaZPrCoRB+96F1QE/20ia11MxYUFXjvMO3qLE0ixNqqIehdj2Sjgb
O50DAAchtuI2Hj5PpANzj/NyAyFc87AcfahxRDv6Ow3L9jQ7N2+ZOQNIc/YctSXg
iNRDZhc4ZR1MBOJQBlZ+zNvZkdyuF/4dUejN0VTvD2E6madM2Sld6274RsT5P+pM
dqsMghTM6IAn0canz6Bqp+6ZPA/XW5NhLyrYxrDCAAqzBPwaDOtQmX4cClZHaQbo
+oJtY/kLxxh+p4JSbofmQegmHf7+c5QKVqfinkA6lwCYI/ilXHITeKxbgqWl6m8a
0x1idmngU3KIQd8qwiFLCUd7kvvbM5FkxOxZNvVwn3o5CXO4tBUiNZCxOoVyoRlT
3ZRXnWRGDPrrIhMG4yy8uobdEpr5/kc5nHdI3WhB/HnidiT+O1dB5+ivcwikC5ma
DfhEQNwGYhaRrvi9WBytOagnqB0qhbB5nsoKx1ILK6bwR93lCV7MXPxaYSBseT1A
L0D9gH8yUN6D/YloReCxZJ6PtmKqkaTvDMN8swRBfvMDcFUxUE6+8WSVOYDVtMEa
fr5rMmEWGf2kHAWgqAAT3USieffh29SaVL1fvmQ3nRHCRo+nZAcA8CyMXVsxyu6Z
SiUMDZFeaJM1b7fX1Z3HGwRq9nOLuC2HbXvuio03gx+ooA5PlvsloC0O7VayfZ2C
GzQPNvWAaIxFm1FUnptgHSOAIFiVuVIQrSoFYJ/H8qGvkZR+rfE9KUI/Ok2g72XM
rJI/0iV5OwkB3K67i7fPOrzuS7d/cIYl3JumrBtdJ3O7vgRl5ZfFBlWOIyNYD35W
enuMf+MgElTThXt92/sLMN2S6lk9HwJaqv9UnswPIcV+2utwBaiwXCuKe6gMUEsJ
2VxRSQrUR3kXZetILQQHlfhUq8vftiIamzMYwfF1XExMbx43ji/H8Rd2dQ2qSVUo
DISXlvQJx44ioWIoxyWzDOfVQjkHwI9k7GUNFxw2dxZcil3Mzykude2FcPILvHJS
XQqvOzXmUUMIb1/AwUXYhxuEAVWwLudwXEuoSMy9kOGV9VNEZXTJSXf7n5WAX8oN
QsB2WfcRZN9sp+gr2aRMnQQ49wl99yWi7At8ZizZN6hg7KvycVCy72h+tuaLR/4b
W74JdVnLuwMdohjj3vBfqD5voi6cM/6rfYj/ABXDlfTkwAaYxeIw343B1BYz9ReN
QVmg7vHWDQ9dnTrgXqmDlSsTDmYCylPGgek0mPlCyBHr4zcBRet8TSmMBJrdP8oY
ytuKWtCcYZTIFwDP0QiiWR8joHRPRtxc//5ex4p13LqCvD+esjB7Ax9IiM12ebtF
f1ViBNiVlarEIyvPYAXkJdgPNDN/pNoEoiKABYWUw4fs0yHVLIhzQoP5Ge3g0vY5
QuB+t/2cQo2cuF6m9hyPVSbF+Cvneuic+jIPjiHj3M2aJcrnTe3xJrK/ZAjQQSFH
wEhxU8RUYzpWIDr8WqmxREHIgZ1+4IniXEw6iBQEUyPdOSPveqLUJSa/cGrbOIiG
ibCk+Euwh2FnmGhI/mi8EF1I7FIyH8qEYXX3PViWHUw1vA9NYYguStJRKPkCIji+
F6NGBZD1drIfDRepvbzuxoEbu3TX2fpKE5RBEVuE98adm4AueZT+O/kNFvpAwy4t
MgvHufEAg0rRUKv/Pw/J0VJlFVP+blcloiV8c3izwY+aFoLfFzK3Hs24P0WRbHjT
SIISOd8wv07B+Awwx+b11yTvJ8ibvUERDPbsZyV3PVIDLalKzCGy5RYk0Cvm1HeJ
ZI6bflyytedULsE3qZFGbaltnYLN49W/3JAZM3MRJPkafG1fCRGqytGnQpBjH44F
BhtST+hDqRQTF0wdDwnP+1W4Rlr50NK+fcQw9tsZoui74SZR+KiwkBtB57nnmQim
N7irgrRT4WRCvzEqkPSWQ3ezuLWuyM6sakfA8P9fju0KN9vFeo7pG57ZZpifaNZR
ViQPiYZNyln8+0VShWkC25U5go9P9Md00RzDS/E3PBS0N8brN75RtIX22f/ZaE7n
8TgUggNFJU0usRhyKdZYzGhAbDchzLk8tMm2Dlet8S7eiHlRVC5ET6krrK8jjQkc
t9ajrv7/3TAKUpeCuuYePn8uiaUJB74CTK8Sx1yjBbxObu3u8nloWgNSXuraJhGO
+d9Dk1o4LsZ+cfQpFWeL0mCMDmckP2n4HQ1licMucR2ZuCmZjXYsjIonWPzbdqF/
ShXtuR4lHZjX5Z2n3qddY9J2gK9N/NBiCPAl/Ca44DXBGDy0gda+OhTx8imSt4NV
VdCOzs7u2hOiy8RQtiubDdTWHmkGJyN+BMZDuh2y09NL1VV3gy7OYvaEGGRU25XZ
hTsRLbTbW0pI+vyKNloD4C+rwsOm+DYqw23nR8Q5icBGr+HYTjksIvl/THZN8+8F
wPmSqX9zd6bG/VTVWHdvSGOZEWOfQVpeRfnidhpJiKjWQX/g6EvOuLTzJZrDJvXn
AWblQsgRfuTr9O5pijz926YLK2DeUrLW568LoohLkoFM/54JlJJI+G1q/nYS4B8b
Ktj/0AJK/MboXePgKVp0U7tMz6WX5ejCMD1oNGDYERwk1Ic+Z0cxMBSYzYuGmVFX
Q9wD955sS3AmDDuc+Zb0wFF+DEo8T+Q6bROA0FokyMyDM/2Qy4Yoin4rjHCeQk9V
JfQ0BuH7vvCC5MotawTN+d80bbubZyabrFvwa466EN56tIucflTPwwLdTdHCz1la
bd9IE7FkmjjbY5l0hN3EeyKyOnao6G5lOCL7zOv9JFfnl246c5ZYlnOb2QSZCgvg
b0SRALSNdMiwYWCMxeE/MMWyy0GiYpGDQMMDao5D5FTSJ3H5TVQ74v4WpgOIdpnQ
6jhCESibBcTy+8cw3fD3CNyKb1UqJPbquZZrSFj7Uhdv8rS8prLAgPMyHLyFhPhG
Ov31Pojt3+/Mn6trBaH8kvjtNxNycoXNckltvYiPGWSAdlo575s643GE5pyn9M5N
UOGcOgMjxDRPj3nhusashLGsTByZt/ymwcPuxjUMLcA5bCIdSD0EUjjtzGI6ObHz
aPVxJ2/dABJPX0jh0EE0ZAc4yMapWgFYhX3T9JaKokyepqlHihSpGLot2XqzN1VA
jQjEYFhVfO0fxLFnPhT3SZ0rFNLhOZHhifrgMwP0Gh0lnqC1rFCS7L0WHVLALcWL
7ow+/JPYwF2HqPG2RdJXgoPlW3LGJkjkqI9Oj4HCvF2RiZm/edqzbgiRWwMPMozj
4a2iHHvvLtTx9pawnk92PF2K4U3+Zmk7GsGvu2xkhA9MpM6SzC+Hx9fqW8LiKH8p
59B8mCZz1/4desFdBjRUyBWB08JUSDJmRTC/0FJ5DFDv+/nHfYceEv2FoE9zGrkF
WDbMCcK+dqg97ql6x/5QE95eW2BTL4d0sDMtBjuj/7SuBiO0ygVAwEv+dpYOroF5
+rGZANMbS+m27Sgar8PosPf72anRswbgqHbBsYC/dUW66QGjHAWFDVBwl23XX6U1
9TocXh+SCGt1sRqe762ySSo4TfYQZ5b+o3trt+Eje93g4yJ5NfEFxpfZlq66krlK
y4UieVJyPj9o3oNIwenO4D868vAUzd71IbO8jDcM9SNinIgLxoFQ5lH/L4wWgNi8
OA5nEHdrL3aXoJtaFKELbzwY1UVBu+zzmByGGy2+fNMZin83dXgchy8rh9A9CTXZ
cylkCbGHsTL/mvf3qvJqeY8GZuJUM6SZk37wwkuZMDtv+Xp8vtjfKkUZQzouFukt
L2xe/oMEuGS9giHCX/3om/ubzOfVHFB4USY/5DftFZ2Vu1JqMGN8WkWalQ00jmja
OrSrC++agDslPUINXLYey+DldSE8SnGw1v4fk9b7t7FniIUqWsUsKpq4vkwdkihw
9fqUYMNoarAxEkBUIf6cTSB7k+M+0Nb/j4VkgX4LurT7TaWBpitT2lx+bgb6MuQs
nceT9ltwx/wlXq3meK24XUbMr4Gn2cKBiRtNEaIOdLb/3J7hEhfV+5UKJIJYhYKR
jw5Uf4JpNx6v+omDgCzlnhBU1Baf2SDIgcVXvXMQHNl5KVGcm9EvZGF2e6SLIHaQ
4wUSau6SSu33keIqQ88gG/6geysSt28T8Mwp4FgX0FmwZCLOAhhX9tyaeVwFpnE2
0RTcvj/StqWK1Gg0x/4tK06sn82iOmJkw8gvZM+FCjab8P7qCodKgXgcWRb7JxmI
18Ix+pqN0XGuFuOY1tEkn7Un0rRRN7RZAETS7/OI7KdSnZUhcyF+sVK7jyZAUMby
wRE+iIeU7kZOO8IsrZCQgF+hAX+jWmIg9Yl4oSOvJOjhrUDG2PR1VWVrlaAOyFBg
uzeZGD6sKBpgA3nmvYwXGdOQBpIsTVcHpDqRJJ4arQaT/JtMzih72XoYuWhCzbzN
ZHZqQ+rV7dGZBqS5dN1bClVEFFeFKxyHJheeTjxooVUp00hUdv7B0NilgXoQYFvf
vb4cB8dIpWtKZ+2dwXLh+/pqMJuWUBMQxODhn1ohIJ4diGFVozzwptkaa8N2zifh
clPWv8iObOlr/f6dzG8zwj0COpclstdClThsMqdz7z+y5bpnYvnCzgpvJIA2ZCi3
0KJVuAIfAoAXKBZ0FQij4LV5CO1xsFGW/h1xg0MAkLna6JyX13WMTZJHS/lvgvFZ
BrLoaOk5rKjNsXmxJ0TyxpDivgvC+749wF+U7TPyr06fvNPxEC2EEJ0zZbo/Fb/M
7nhBliVweMeRdoixRv69eZx7MYzoZIzZKCWDTNhpemnoJNW+AEKNGDVdwj7S3F17
ctYAzFjOybpGx0Yjf+j36eakjDKzDlN80mt09lfD43C4k7ADkJcUR3sR0+ofCvtA
IWevLa90+ou0T0myvaaBkVxrfSvSCJza4G0CVYOCwKQEUbaIhD2fHiiFMK7ia9wE
eOUBdlyhngLDn7wHxLxaR7KEDHxhezk0xV3JDZi5HfFQ8eG/oCZP8ybG7C5c4Ri7
uBj8HQOZQ/ZRbKw50FhgfhmCkKIJ0ZBSl1bkoHYs4S4k9aBcaRAdxCa7wYXYN0tX
LInaT9TROPNY6fLimhKG9f0fKlUDdv4bwNqZW4uTQfWjMY/GpyWXqZBYIjreLqVn
VJOJLNUAREiIKgraAm+BfJskjS6rbyOzwg2XSC7KBLoC6cT9kCc4QCf2d3HoXdSA
YTwO4Lby4M07BKGQ5UeboKHbmTMl9MfE2en/z7kshI7mwM0a2EiUvA6aR1cAVPwP
wLtyyV6iCc/s+GTVQW65RTJ5uKmwmZAbZA6kt+12Rv0xY5jqDjd1W+DG0LPQu5SN
O4tFnSb4c8RinnOI5a6OBuaw5SUuuGKUC0cr3wsAO3v9q4qyd22KI96ez6C/R99i
DIoQKoWlCQURErMmq0zLSvDUaRLpBIOwxrOQkW2y/DYT0AA+lvpHDB7w7J3qeNAq
W+3rSWEv8igVGyzFcpLTyxG1/D7P9+Q61otsDFZjfCYeBI3B8XwyTmziSORy6r8f
BLqbFgHZXvDWBGuGmLIjAWeBlu3J+0lHQJQJEr9RYxIRZM9x/gdC/t2nFms1jWVc
Zh2qoNeos6mCXgwys9PeftrE+Jc2sXZmV2tNMYKwKBYWUvuQHyocg3B+AAJa65h4
2lmUQ9XuR5ykpJLTx+loI1aJ1+h7Hy8qTsqeJOYt2QDBNxo8xfnSeBx/30IMI1yE
prDWpBI3cpbQ3FxGoRwof9eTKsFeC51euDwc9fjCFXO9KlHw3bwgsM5RZ0sLXAj6
CkdMt/naqFfikBNXyOENTuHOB4JuqCUWtQ6zRYTomAjIsKBPCuIbgLsp//nZg4We
EVs2i+pEo0rHQJ94RaFx0l46IZo8ldQPAKIPxg40ZpAHxW8WV3WWvlIVLgmrc2SB
ovaUb6UvBZBKBT4pwhbMzvOFZ11dWzopRC7grEJllyWL1ojb4lIHXPRd3o1DPvMD
5uz5ObeEijnFxQA9xKlGXX85g1irW+iumhjwyKyXBoPKlIgPykota1E/KwmUykA5
hhReQFHqde22qCQNnt8gte86+gGEEP+mNDIg5ehSEUsjwUQ3LLIZn/J+gb2NBOKI
YriyOW+qLDuEyRg2zSsJjKFlk7iaE4iKN5uCPXKddhF081B6kcvlfHuvlte+QcKS
qx15MzbmIr2o+E34FZtIUXeV2DU6vh1UdAkVd3HHMhbRa92PCkvRy1f6Q1KpH9Rg
0fH7FDK0fBQDvnl+RHqwZlRI6F2K4uAli8gHydsGtqKrfdlzMffs4a0xwqKWYvi+
TnfhMM+rchwrn4be8naK3kKfxweK4Za0XKgCXKJ+1iPwnZB6wzHtI9uHGAv2En2n
hXyET/qw2TQGjOM3mR8Pshb3Qi9H97C9hrB9F2NhYQEaanPCcINoZvyd5cbdRRr7
OUrZnUMyeww2RudtjcPSnQKvvvUbYd/CKpQtQG2OM/DqBRc91YTvoWe0RIYvqvB5
6fDjEG3vo7/QaSEwGH7FPtXiJ/wPaf7iu1WQybAgEScRjR1N3y8Fw0DELXpiPn7F
bEqfLbbCbF/p47NtOTpSqrn+73ZJ2vEEo0FLrWyngdVqa9PeOUsC92CzJN4uSO5E
ZkfFdQG7TbWPY71yyJkRkSi+Nn1af9pkan9A6zEWYouC6X5k6ihmScJYw3KoopNr
2V6TwFRpSHiIoZpIboU7Fdbbor5P1ofJT1zcQdZl6j2Eu99q7dXF72s+7yT4bxam
ZJlgRtZPz8uqXXXd5UyFLeOAfQuHUB4YcSPTvWZpn3bq4owtSsH9B7fxwm6/+6CO
2e3SHgWvuUIzMsEDhax5/6MuJBPpswQq8MqXIIEFlOZmRHOPvPlVcuNs+IOygAsA
zKzoA6lUkkO0yVA7buexSFFZG5470fksmtVI362A9eF8ZtSi5Y9bphDBqqOZ73PY
rEqrMMO2dTXsnZU0n9rEcMyoWJYJno3fcIzDB3eBn4I/PAADNQ8M4jjzsIvm3uFC
3D/bwvTPTET9bWmTpxmGlct0VCm8lLC8DL5/pOYM0GCFKL3Qg9s/Fk0MN9OPc2lK
Iyfle2vFKdtY+6vbteZ4YFkt0Tdjbola4D5of5OXkWPyvF6Q2JvDJa2JkH0UYHg+
qy2isIAaKJhgTxMo7L7CZuK3FbhSoiNQKsQETtBf9Y4B3vKODUQVH2scA5GMjjOK
EmE5OSIr54kYt7anyLxlNVxXlqqF0LouImtvLLURtq9XtP5fC/JeYC6kd/VJC+HZ
wpriGf2YzFSn1WtNJPqcSU5Uhz+2VH3JIVNhMoyz2/ui1z9RprIqiJbLq5FF2yT3
oz3yrVpAIfcIGUUsjHqPBVfmIkTWx+6D+IIVf+UpNSVfqzTot6hqyBDLrdS+4eM3
JXoTsoNv8psqn6AJQwelV7SndlrvrTAHjFv4Oy7mz0tO2uV7C8F0FR4eQ4ui35Ah
TdLbSdG7HDd9Rlgi9TTOGwi/ZwYYullQ/miA6QIWh2hze7J8tGbf/BW2g8uGxTdc
yOKvfU/TkgJLoXC8a0m4Dd8RbMjSqvEtxNvM9kSHXWfjfpwBLB5UYNDh9twCENW3
0lZh5wvsv6qcFEqMlGEtdmdJUgTdOTkNljp/uvB4fEuXRPQKLgfK9CtTGoJJ178N
Wi6iXs5SkKxu+oFciD2Ihq0VI9MeDAqGmxdOALs3o0KUAb5IiAXbY3zq6yVmJ8Al
lBaNhUWJnKTSwTLz22kaiD/lCFpJmo7HpwcCw93oraeNwZwHcrn0rrWI1kupZy0e
VnJwpjO7QN5Ru05HtZLsenF1sx4fTF3D9D3auN62JECwWz5hFid7ZBE+CYlDH+bW
3Iul3S5eonkYzDLNgTTjHVDqcOEwVRZV4nrV1RCEhcpWG5T+daja0VHHCtBgWZfK
5fL8aAeHEyK8Agm4JGgUaOmvnkmCgfu8G0csJmeKntyjblVDGD8HyRL8yOWtsWW0
/0jeVLq9aAbtJaKC+h2+0c7coY68b8t2WlNo573IPDiNpNpYLfvkxl+FFjbXIvE8
jktinxNtI0lKBS0fvxHBqq9NGbRtpVlwsh6QA/mnm+EsjDir5TJmuzq6zQvVkDvg
vdBGzPtr0GSqZi81FLT9w/RSbU6v5i3Zt8rrytM46rt8xlQwtPgPuMdUfU/kmXp1
+JQ3a1c47GvC6bJQkLanQepB7F8NTAP3crk2JJFew+vO3TZL03FupcBcOuKn8eOG
3OSgAQIZWev7+THEjnmjwSQcgS8XkymQp2DmwnnyFo5mD+HBrgADxLXGhuMwm6qB
+83YcTIcHT/w9CExVqScXQvpRDhkinp8fwfBd4kwXhDS4AWV3/cJO+lQDwHH2FFP
1aV8dffEy2DF3bHCeDvWiSehi71YlHWPBPd4Euk1rjjUlnODGNtvZo9NzbLhmHBn
nvZi5TEeyzf7D8N1fNZ8cqxSImcE1FuLGa2Hn7fwIN/Qx2JieCO6uGdydoJsiPru
fSs2WdbN6C0ODZOWPgwsiDvg4Lj4TTIYaXs38RBNxyhkZXgmoWimb+7UYooAaY+G
gCM1h2DDKHu6uR17GB3v9bEzNBRaS2gh1trodgBGchtpwq0GlcYc2SUZOk05aZCL
u3GB0yVM2G5m32CWP1Wi4Sl8+So2iucrIxYlFjdgUzdhLtb3ozzfBRXeVyF/aski
yNNAlYK68jEn30G1r/Htx4Ef6RuUahfjDOtZW0VfAdoqC2OI13/vAbEk8qI8Eil4
5rnMYOx5uqIZr9fbtD2AAdUT5OfONsfIEnOVUBOCCD9t5MpejetJpAf3ziIGagZF
raVgLJkKkFCXecfvCAXq+F3dD5nTXaG/3pkFY4jarEkNXITYJoflkag3M5XXjjL9
cXb9AtOmfbGlxHA1ohWKk2PGW+uImH96V7HwEWCisu3ce/hHF587aCnHhf5YV2zr
rfeiZQkXykrMUjrvFaJ9Bzhg5D6p46gzjU0d2JHzWZL6zhTdXirsgDCSk7yIPnq8
vmyv3ALMiVIBrYE38jabPlPwhAkg+MTmSjjPbSjl8D4Y2VLcTA4D4ktizNalcrvF
C66qzk3xkRclnyJZRiCDkNja2Z8+lYNbLurCa73iHrGdjk3BYsDWwvYvN5qQ++RF
VUMkm9juGpkQuK0nrpFZqNhq4YfCtoGBNJilxHlm0IdqxdjBOMlztWcFFKn3likp
E2KUCaFCXeZZyOm13X31i2cHM7OW7mel7oRwDKIjFUd9fcpHp69pc42uwo3Hp9UR
qQLcn66Mq0jwtAJcWsZyFbSo1NjJaZg/n3LKYY6ycZH1Fox5trQ/+GIM05fBaQQj
XER3StYkq05eOYWkJ6TqsqxuFnCaG4DIWCmxThraiEmbn2mUFvR7zvT2ZzUw6Jah
efUpofXMCmZf9j9bSyoeGsOBnYCWkHB/v0NlQULI2Vfg1cvmYH1qLe5OSlfxctAf
t1z1SjpzknYo8Ag4UFj2roaC+SFwsajUEQH3MzH7ZYGTP0wEH1ZO2SSS3om5Y2DM
vgT3hl3uKkejWbF6q1DXpatMGYMpEDNYfLOmypHy2pA2WwwTZpkH9wB83rvM0ucw
3rPxOZ5dGD+9XY9fnmaqC0xkEV98B3T6qfpHvAANgNqYDpUqcB8lb+XjvQ1BNTY2
jOtPEupczyQkI3Sr85OCqnR904hcJQlglZWByC4oBSwVjd5Tqa03Wsjw48ak33P9
cGKBlTGtNVz14lO0byFkoBR9WUwpXzJ+pE/AFiKCLLffzD53zVO6ulZ9jG8xRmhr
Rl+XYaWIXk8aa5Od0deNYGTkO0Lji29b6/bryXVde2dmGitXhIFwZeKXvhTsf0jX
NtvR83OXJXJHvKiQV3DPRYUmcb5wsPbrN5VBWwyB6N7qLKpf066ZjmzvL3MdJU6A
51sG2JHBSsWQzPEJwx2Oa8MqcumAadlgABYHAGYKiBa9s11VX2qVhdVEQu9TvuK7
ftZgqG+4sG2bPT1q/qyAuXBOZ0rBAfovj3vbOyB49FqEs+oYYXqL8GT3R0ZWxOsy
72IRCqDo1n6MxyPiMSI9/IZDXbr6DsP2L0UikqkeLeDG2RmtFyQequZaF08hlT1O
f414ZvPTnTlYcqeXGA3KJBjUp/pVBrKgdFurR7LBWaixSaFyGnrUGA63WvAnKn2X
009hXiEclpPoxb//+Pko2jXGCi9PRxPOPn3CuWfQgN1c41cZjzKCNFqal02o2txS
O1mFzYAAQSDyM8VoGwzAGi+vU5snnLaqOpWtVMMQ6CRZ/2F/YltKZ24sJzPTWoGj
wkS0GgmnEAbIUYIegIQvecTjqniR8xQtPicRoETcqkdxtYeqMwMGXz+u9j4p39lo
pBwYpvYu+1cWU35LRIh++4roVaLRwVaZ86sLXQJqhkjVZjygf/V8Er7JFcY7s3sZ
oVlz56XwW11RPGjUXCMsZgGBi8uBFcz708BTlK3cVJ9pICx/tyUl7bAR+RGCoVNC
xKoGRaoAAAO/HXCP3njlRZb//6M3EWw2KQlYN3lQZajwkc7D6JMfqZDtdFJQDhBF
IEeZSYGC9P4plZCiEksb2+h2D/DWN9LzEulYwtJcSRE47BA84Q7Wo+kVTBqBFBaF
66v/e3NcUvSF/0+g4tJoNy0mkn+FxVVvL82qZkobgfihwRFkQL1TZ5cCaWUCGB0F
xrJ832GoUXnxzw2EHe9xVYtXgfpAeDO3ucf8bUlzELLv+LNSD/9/WvTd946Q8Z4v
KEb5HB26nmrXJA3oLLH4DNvHQdKVovr5gCB7rBL0mBe+9XjHBpRvsHGB9esUlTUm
L9Wdo2kPcO2AaAed3mKyYaNXcs1cnQl6fdltJNbLehzvKditjFNYcnd6Pt3S905H
ddHMVRv5YStmC69dvdtBL1Aqzp054tJ4eAAWShejiifVbdRop6AiFSfdNoTrm1jr
33FvEpb1/BbEaAL9JB6dY6wBkWZTtC482QjUVn8+Owp/zA3LLxGkTbJBpAQGAaFw
7iy3j/6JdqZrKXXE9vp6r4xQoC2w53PVsBY2KmIaFUuIifNyc4lLD3E0LA6Q6cKp
sNxm7qUcaLLa3ANyCP1RLPH4xyXD1Nb5GD3JqTiAAj7rMpxXhtxjV3elj2Wmj3d0
JdimqjYT4n+lpInQ3eHm1Qk0fD9Vg+KaNQRSV2Z/umehUtE9Y/5FVAHXVBFpH4Hp
qkcHHN6RAfrEkK627bwxBTDuB+pFX7P7/h45ZhJ+ku23Q50sJR0FoWaj2+T3EK3L
kOD6FGYmkOIvGC1YpFOKY1M3uxubOmNoAVizTvDWBWoHYfXEVJK+KrLvyW8yVipK
rS7KxrIRV2v9AhHCuN/3viIniW1HQEEflN+aQ2DvmmwK/DrW3KQxtMtr6uTGTZbD
XNUWTu8N3Uny02zR0t3lKCdWTe/2nxaz873rMPdYHPBUdCyJnZn/ZKC792nTIsvF
HAPPS4RoQg+KLqGLqwnRA2fo9STf87CoCop3rUdNQgBzhPymdHkSg9+f2lPeXEzt
OlZwfFdip18sfc9cYINKlWMkZUiAhDNUF+rneYdLIiCMPvr/UVVCw8d1aBTZxRv9
fVPSKhSydP+7HHuzZGyrLpkQ2IlZzWQFlD9PIcgQF6sgcZuCTeLi6eNcVoJKjany
/eOCWFqGuFy9eWIVwdo1H5I/QXDF+SCJOtQy2N3d0QOLDJ+IceUzkpockQMwlRmS
ZYgRdFgCamCEizehlqilcspxuD9vDOQZXcpTyHj/fnwbV2RMWCSUSUT2hc8oADDX
3V/9VKgdp94XkTHDCkaYBy4e+xeYw4YCIbizI+VHXBNaEo0IrBi3e8yL1bf3TqUO
Re3XZcm6T2neMF6W8zLT2JfnGKuazV27tIHFfxNLxEOUaUBx4CNjX2cb6+IN5S7b
EDX0cv0+DEH4zVaYKBLKQd/6fAhVJfuDkpyH2z8ScpuEYY12Uwr8RL6XeRQIh16W
hsCdqzQyew87/RWZlfeePveN2Wf20Dbwi/JgLVQ95Ri4N4Yz62hXpCQyyulS5/Gt
PM2h8R6fIwO/IC4Bl79PxnKj/L6BWbIOr4wsoY3snM6a33DLem+UWiPphXYqrQNL
yIE9Aj+ZFuXC7pYT3v1WpEPN/iuQV2oUYM8VUbMl4KdvLoXOBvgCz1rpyryd02ZE
DfJMWaoIej+0wl2yZCpp+AlgweeGA7M6vK9Vw3FtB4ObU/aQURxJ5M2IC5Oa9S9o
39ENT1MutGR7SrTBQpQZzlSZvzM1KI8Qrj6XYR5GmVgRyoTe4LbNp3rUU+wwfKwv
8fEI5SSZcqQ+pWXwWVOWW6pCdP6ZIARCS+Jw9YbLketTX9UiGDdK9Zc32yMEN7zr
9kyyXZXuozY1H50qhUOKfca4cSrPNtWAJeaF6cDZovA8NI2wuPpyx9r4F6YemjqI
gQb7+zWXk9+T4VsfKGhjYSqEe3NPFpcrgT1djMZ4PwSJQz7g1TvkDTYDJVJbcIga
9AMDvq7WjyVrJnzq1qcXtmfD+2R5GA8oZQBwMo1v/GQ/VW+HOtQ1GXR2hHVQyd1z
izI7Ik+0XNugC25r0kEJG55DRLTYcrCtjYvdJsDCPpcrUu3YWVU8IfNGQgy51GA9
ErJVYwcIodfCQdko3NC3dmw/4Jg/VWofF9+Os5+xvTMmfUbMy/YR4spYQJ+50R/r
AssUkC4eaT1hwbrGc0X+wkxsYG+XT1pSH7Y5XN1oMveSJElIXFODxRZth49wJSKb
uexTuvyGqIZfxWj1syCwGxrK+5EDRTWyQQhsPX7jvrOzQAOKEEBSrcvbqAMWQvOy
pGGkr7zqj4NCSM+y4Tr26jhhzAwuqGj0owW3QV/KiuJncLqwJknb8JRXNL0d5KeT
N37S9wHjp0GiM4EJ0KhDxQVEhsIJbjJmhzdn3icR7kV7MpaII0aG7jWi8+6R1UYR
zF52hV36bU7MHt2uL4xoQRpnRxYILJaLg+t284q8BnBz6FW7RYMl1Lir2xAET2kI
JmeT1ZX+mhHZgJ84OzlswEP/+eeqJaxWoUWB/FPOgax3eosBRcY7pORtEwy8v+eC
r/38/Mt2gEV/2EnBdgfJ7sChnG+gQ9AImIl3dFGEiIvgpy78GH9ct0OzpTBr0NFG
f5z2DAa3QRoieZ00lMpaU1L9kQ56h7sWxeLqjU8WXQFR8oLDJMnoAb2c+xFPj1UB
Lb5BsUxwu/yQ0Nnom4xt+rIv0i3IzqrTWlDbSAvKO1hNzvEYZGZoRAeHEQ4FUQoM
tlHAlLF8sg+Tp5VR6uaQAjpVUlstd+ogH/Lm1x4SOqOvHf8SzhGBsVYEFvDP0qGF
tKrlPce3LDRz24tdQbZEOi69rTDstYCViLDPBkjwvbC/yGFg5cDIKejzCJH16Vxs
A3v9mWBAimDo1D+XT0TgLUq5EzQmAqgEy3qF3RWNxZzlur3PEr9yV0Q3pBRvhSQB
0KLgp//6N+vIyTMQNagKLeGhcxaj3fiDfVBve+NW9/OxXViMYCTTbd6hx7IB4whl
VS9I8ZUJfKJJWsTv1EWrIBdCsyFda0y0AUa54a8U0diS8j8fC9C3vtMWnAN0zZ1I
XxVSYER93M4UYVlk+So/sdN7vkVdkHDMHyDmv2VTDyx2dJe0YAcsxBfZQPQNCvRw
qXPAanQHHr5SsS6FkOrAPMLvEjxIJMVMVtS1NKFsmAJbl9eA6vvw52Dxx0Fgg6vD
ufXMFob5uEvNpWwx+WOJT5Pe4YVsUZuFfv2tFr7M14tGFmAc1Qk8K6ASK80B8Kyb
zlmUFYEfAC8RMzaTI0rhG3LtipMG6Q69xwPczYroD+BZbnunlpfLbxXAjTDtIROb
9fXT0ToFKAhPVb3/J8rM2RNtS6BGfM6hLJoWi1GvwH70c/La6y8z89lQzs+kpyFo
2KYh3b3IngOGaCdOxEsePfX9LoQbIZiAl5ydVcxsfnqJO+hwy5x78dPDyD+1jGVB
VNb1XR0DBWwaHh6Fqchl3E688QvCy6XiIeKKM5Ixqnk0F+clkaga4IZeXMbFDAus
3y8ylnlAOF37Axy+TIKL1aWGqRiG93iU9PuzkOU+hnM2SfiZRka7fl1ZwEdNlC7T
ldwv1iiGNT0/LDxPI1tXtLu/p6DhH6c0UWGjLQdr6cDg/Zq356//oJdjZNI+RmJ6
WckMPRZiMADq9YYOERI8l4Yj9n4N7RN5cJgJ9yEFUJVuhfeUIKmA2+Z32g6CMf1z
39gZ7QqRJmZaMGaW7jovfrvi5+weJGtrwQMn+T1P6qO6WmzacyWu78oDTo2w2Y2u
XJft+8HicLz4kMEi3fo2XRtC5eIp8eukp6kEnt6FYOK7hE0T6AZb2wY2OV6bTJPH
7Z7TRJZi+s94FB7tHyNcht2xXidg5Es8Sii/5jlzlOgaeRy/p+l5GORx9OpopTXD
ffVYShX88D/uri4Ld/O/bsLBjLuaVk+P+e/4Ie07Q9Jn0hm0Vz5aNtwkAnyqhsho
EBe8I1PIdUGNnxMhaAOIC1mVwJu3ImNedCX9nOXJ8RiZxXHxlSq75SKJ/WI3ieJT
pG8gRGphmNALjhhzmLvzAuMQW7qbsQ1kQLydSIrGZpiw2RS0BuQZ2CWR9J2lr+S0
XH/pHdYiMMU0szAXJaEE9MpIYQsox1d8rp9F+nH/2FMifHQ7kJF2Rc/2rAPpdfPj
h1l/CaZSDAi97cY/BjncGwbY74cWLmkLjumPsOvISJ5sVkiIrcT/T7OMKetl2Io9
uWH+CRNihBhfm/xZ6kMOne6KdormLSJmpcp7+MxJhHZunx5ALa1W3vGZtoZxPSxD
jlo0GhHHRMzi0KCm8FtYA+1ElUj5Yi9jbRv1B90ANRhUA41HFPJx8mIWUMJmSdWf
pgIwCOfrZcoyc7gFmxC4QJWXG8cLL11vEMsnkiVQp6La6KhhhV7muLyoXSXZhOU1
VdnzszoGDA6zG5V2ywFlSzUQ1YIAI8RfZvaN7jMgD//RTp2JSugGHbD5hBYcFI7R
ySBfqo9ZrLDhv+kdSNYNjD+KDc8SXmZhTWs87TebolMAO9o+GwbKbxF+PtfQEa2F
rDLK104SL0uyB6/N8ib9S72TCA0FqMraa/V4zlgc+u4AFbMFbPRiG45sUKv0up84
VGjT/sy49HlBy8/VVxrTteWJHyOZbRdFmg/PjK89NALabaSpBb6vc5gpN1Df+26R
hJLPpgHfQDjDQFo0aAtGVxcIeLY9A12qzavJ6TPtybQfYmq+aknQD4oXSKc3VUvV
Aa0+GcbcEB6dmPEItoDTBS+seTZEfD+9Wk+9NBGNXvRgwgt74gvdjRmloD3rqheW
XT+1/lQuxG0Jci0Fx1R6MMJ7eOBAkyBrvyfK9CmIKuJtXm1UI+P9euveJkJ7ENam
gjX8CM0wuMtFLbJuzdVOTOKMNpCfsMwLNgqNBog0B4q6onCVHA3N8WXmlOB3eBnw
Ao1RJYytTnSnGQ+pt04HGdde9/cwTn9B5UTr4q6VIj7Tl5yFhhFnIWqmcuRz5xyj
qSrbD6AB2MkxWd3sLiPaz6O2My1nFZQJF57qNnyzE0uUiTNw97QsUw7Z49zy3srh
ELlEDXNelOTKEs9TEYk8Av7wEJjE06k7nB/fLtiBUs07c9WarJB7mHf4TxDhgfgY
zPZ5lQWLApa/yW8PqP7WSggkwEjVYpeK0ATUnMOciK1rCWItipi8UNS6QMWDYTNv
aSs1Piau4/hPCWppKXxBos783ovUYkV8ppCdt7fXlym0mEPD3547iFmqm24j6gc6
3Ys2xrA1GafPeqEtEpY0TvaM2dMHuPV2xodnkh/VHzY+gZ+HbsHILAdcneI9AvcD
WxN9ONFahHBaXdD6cUfui+COUyMLVi+DQguzqkhIGEwyQyvmqQ9I2TGVRNdPxkOG
HF6doOHotVz76iTxWurhulmC9HimxAWYZWduCdYEcZGf1PzL3cwhduf98PIOnupL
CWGln57O4nhWSnyvEysUXdRCUi7BQc1ZJq69rNdAjgtyMtU/k6fbpLlVueM4GZvz
7P+YygpNRvhRqtOwd3ApKT14heNraoB5bPv7hh6f73Gy5SCZ9TZQfnEjG9tQTxz7
neCG2IvSh/WWY2CSTLYlR9iUgvz1oxbqZxYoiewfmmjvyPOULDXdRXgBzBoJGxxm
NLe934txmc1VP5hVVVcLoF9NqsPkmxIjIH3ztzPsIdrBBjLuwZKr0qETdtrd5npT
oY1SrA7Hj8r1tAY8iSYi6c631d3ZK4BZq4DAQpwO2w6TyjcnzB69EmMBGBcEmhsv
phUsIxxK2EskXLZGZPiNOaOgTCpX7CJbdj/NuxKq3ouuFeVZya2rOEy3glvNteI1
+lHNReqg8dDLvs66tnEnPvHDRjtg4dX13fIJUEh5R6MDeAJt9DSPo7rH08uWO+IU
nSWau17i1nwsZSh5/z4CmJl2G6iyweqfIRWpKt3S3EIad5fstiPc6LMOPV9motbJ
98LPIg94RfE1BOev7fKtqfpyFNOxQCY8u4ALUtNTzZ62um0nDz+1nI8T8ncfV8Zt
sKtrfpMQalZ45W+YPudq60jnFUwzPaLfbSXfRWhzzAmXUoSpuEVbIJqrPSTeg9Il
6nzLyiNOxK0jsDPb0Dkmt+7gsxv3Ir34F5BPeQOgtKWCi8qT8viUFUEaWYZ6q8TX
ByIlNnB5moqHM43jiyRCB4MnZsVrFVIcuzc6SpK/7nsCPfvU8GSa5snYYpEK5bzc
AGtjxznq6UFOZoxi0U1XuF6Wk5qK6yUqNI3ZHd2gHREShT5ri5E1n6xH1eG179Ou
kX5yCy+2bmMSwIvo1tU6Qyl4ffx0qeTsa9L4YVnOe0SReLpziRRArAKVmhnKxmPv
4YXDPnaCARysPVuzziJHlE+meMTmMDR24KXflI9+JCLqaLAV0kfjdgyeMKadNBRr
zHgQk1WI+faNNR/ss38fGsDPZko6vKdvQkXWTtz0fITwohj7/hWCptEvc3SgPEUF
XTokALGy1zU0y5CLjHHOtKchOBIjcg+O5UK2hbROgNC5zA3DftjdwoNU90fXcvon
wFOW9hHc9+O3mUBKMXrQavxoqee2tpWXzMWFVDcN25EtbViuJ5R4/JO4enW58+IG
dDMN+1OJx6zX7yAJYfLcVaRbo+t0pql6iJVIxNHg16b1SMhbD+7if3CW3TzSTNx+
hrh0MY5XCPjyHAyIjbyXWHGJmaz7ivW8SMjSGpgcwa5RbdC9U76pdva7cncnD60/
VZMTOFVOzeunKDvOjFmXbSDe5Ji4p85v2RY40AhN0EQ7o+L9sMDPPVXStOPzd7op
TrLVZVf2HBlMft7q9VJPTFZiolDYCtwnSqcSpThdnkG9Lq+/XHvgt39fiSwon23C
O13W00MpvqvQsklCV9mzvg8oY4Rns4E/uQCsCAh8deWwng4oNjIapBekK1a9WPIn
rNuFIeeYD8GwW878IOH/OqBnEZPRHhv8M2378cu6yLa8RuDnjfHGSUPox2oHdR/J
H2NlyhMUGBCDxxYA3mHKLkMBEutN8l47QvWHomKXsoPIJLepsJSeeZYckybm4zSu
TvfI407z6SYH8GwuSKbKFuQUmItqh+3KMfyq1beKE+GS6iHBZsuIMgcMoMofsdy2
hIsq/7hOPj8zYPmwZrmwPqRpJhYgyrA3Pzkc9Po65tEoOaSGDlGJymdB8p9SgMWL
33wd/rJ8lg0J2biCn3NnuOes/kuO0I5U3eOx8693hs7pRCOO5457W1j4GDPMt9AS
i6n8ODag0JSklfZJr0fwum66lwNl0yYIADqjyixCGXnGtGBRDpTo332LTrvyUHan
dvnIzsHO9WzIqxPMJCaIYyVqateT6RHT8nGJqu+HS9LxT1rl9Lqb+KxCZCgQR8Yr
HnMRs4B2AlHAMJhn3cWNarqGeS3vmePVQ7CrWR81NxnRQk6nrfqlJaJ5RiuRMcWm
zHQ+Nqijip7B3dUfKsDgQNNDL6xhvrn58ge25789nhvnxNvUq7k/KpoM/SYRVGD0
J7SnNBMMxxH1yI5krSrWzcwig28m/P7UuA5vG+rSYCmbiLjJmP0QQmkY9An6ysF3
6UHTKu96hj3lRa5IXAPnUpXS8fpsYCW2Zbncqqx++qPFuI5f8DFlUxGmmEixD80x
Ru6QSvdc6KysAWTb5EnjWT7Yh9aYn826Y4KoORgrSKmqw4ol4KheL7iAkP28zvq7
Ojqjvdj1t7v+pS70o8oJi+Zq7MQbP2NqlJb/B0evjh6QFRG2ezgrqWA4gA6fHxwo
9e4xTJPpijGbAaD38eU96XDx5/Y4YCG/yLB/aGPhfqmqM8wvyS+JK7LBh0PX6uF0
tv9i5fso6FPu685ROOhSqKNkiFUTbTBc5h1vQ6nrpTTdmSRSgMqrBnpEntH6OgRo
bRc5wxvUcz5oOTnrnr5lV2PcYtUNqreo3IAsVDv95AK/dnICOsMH+4gK+BJFugQP
LqDSABiB28mTqqXIQOOJSA/GaLtXYEhp/g+IOFPFyKXKk11nhh1b7g6bQ8EpwBo2
XmX/iczOHobnDUp9B9v79tPMfbPP5WNNh/YtbqBQK3xXwliU/lkoyMBBIMKRCL9j
hyRnDrnBCXdIS37sFX3xFLOXRJUOBOrB03ZBgN/GLBsTXDZfnArwAZLZuNcO2h7h
7gJQADS5W2Tm859X3uUtz+x1ScNp3kgv67C3Pmy1qDsVKuR9nYS1SxU21FS/Ep57
b08m0cr/DhpB/wEFMlxn2FI/4W5qUrvZAS3KgaKoGvscz7dpgVBBJ3k+QnQvGguS
crbNmZvBdR3FFk1LTi3/1IH2UGbWGpEoOtQom6C5HlKKbw4GyqgBaBDiqMY0UqS4
iHeLJxZ7Ug2FD88ZYJ62OVwkGmI7R8IkitmUejYtw/kJMu+//jDxXIVGJY8IGV8S
dkwnPxnAGTCXbQ9qYx4zOyUoQpYn/23+hX/XdCZz+aa2pLsY+cPvNNA3UK8o3ihG
4R6DiygTJpG/SR8IWLB6T2oIcgRhegyfgBDKKHpsmk8G/Ol5ejMPW3VnW0Y1me1I
51IikvkO603eKznp4QPWSkRxD0HADbzzXb6eF1KaeO2ESMrz8h8Q9lRPTyezdqbq
NqYeivHRtf0sBmWuV5se5K1HHbp+nN/Rk9+4teOfEJVvOIH/TPjBbrg0hvcIueSb
R56aEQXoVQPs5/tf+vRMRSObMUKGanzfFs1atvFC2bfxGaqMfmBKDW0kSO1FQRh3
6MgjXDZ8+pQCK58eHsNjLuowylFVqiY1VCJ1RNfR9uimoLCnawwqu3kmKZC+t14n
8lAr+lgMcpvYI0io+7Rwt0RQ/hCCNIDCwmkNc92mpaje9VWgesWn2uVTqEFTdQq/
ARdEn0GYxKQRa2rVvl2fxnfvGCGNndF5YM90CMFGR0gZDauVCLnfBRbIsHvLIn/g
9XWf+TZy43M0tmpQDiBgXZ+NKyyhg+qDfUftc6+TZ1Yn1u04hSZUeUFmgOr7H3tA
y9uZrB28MQmdKIR/wxu381hrZCC3e4psOc+NF/nQtCMOZg1ZAp0V0sndxFyVsP1a
8DdhJrR9Kzkefn8v+VEsUGiOSQZrVE0L1KI5g9o3ZrfshXuSozoBVbqLG1GFgSRi
UCh4rZdU50Z7hR4vN57Qk8k7dfhbhR2LX/h09c4O5hYEcKylY794kH6lfiJXLGxw
pemYjx0lvODrYAsk53tHRBWhUKGXUgxzEIwFSS7zAxPhr4mRH5pRnKrAxCVVgTTO
Z+4zW/0Sx8wA0qdRH/boMib2eBpnBF0NAXUuxJtw7MvEXB0M6j6tyEh9/dUykem6
E0NHs6EeXmd4RSGD4a3pOiuVmyINrnEwcxB5jMStX2O2mljPmGUUA4/JUEPQYip8
8Ztf3QtYI9d9J8JKMmYuDJ05cqHSiFOOYiFzzGj9Sha7/v8LVredZcvA28txnpqe
khgIcKwvej08yYWsw0m6ZKV8WmQWtyAEun/1nWS9/o/a5H8JF8Js6s8KDBbYMPWA
WsNiMQpOLnigUQILVZsqRW9sGL1RI+3FK62vXv3Hsusy33zsE5YwpoER3LKpuz4R
sT3PHGQP82Ltm1pN+KanQbnydUnsyFefK89m3PQRCvNegGfOY8MUeeKjsaR/q9S1
FQBemCp2hmivVgOBMhODQTUXhj5+Tb7Y6KR4gJ2Gm561A04Td/GygRg6DvcjslWX
UNX7wIikxknDnbzPNYVzCdIg13D41YiizLNMDvKgBUFeqZvGfUA78D/YP6bl2C1T
5luYitSfWSXSOGKFJODOZfsBnq00VaiJ9KfxfJ/hnRJ5AULxPi5eNQsG1V0QPR58
URg7Gc4JSQTnLxfTY2lHGStDVGcG0l4Y+rOL8EtlW29h3EGBI5vF/mUYw16sZAAN
ESchuFLIMRjopbayzfMnvIyRQ8Ds+U8mml5K48NEoV/GIQP0fwUxE6ijA0BoukP3
6qFf8YXcISt6OxnALhQ57uBA+JTE+1l/bkkU5LLGk6IlVxQQ0r9R1xc9ni8lsISP
942ZidCF7ZLFDcTsKpIQnONnZQeJ63BlbCqkei1J/1r+qqkB8Ox8r9RRJI7ik/Dz
YUuSqxwX0B+t03bthpJaDT0Mx8J8ktKUd8ZLYqyvaLjoAGXvMXwT3l45n+YE9bLp
aupxyTwt68zRe6p18t4ArYQdlBMOJCBMxYb92sQ4eVnf3R6NFcBVqXpoKUGdD5pK
Vvbv8NVVPQRzZ8y96BqqqRPQrZalHlpenO//0kKdfwTEt+nkJaEb9G/rVmHQrzj8
0DDvPWqBvKvsr7GSGXS5MnyhRJB77nbkvn/6EsBQvHT/Fzjczz/GzL9/7fYp0sdK
cfcq0NacKEc/+m6IMV9kFXk3VxHjPj4IksiC+AR5juwJnZTOe2xhsCW1igJlUBO4
AW6wP7c0ryfmu5WC+YrS6dMimgFVUIH/46+71AeosgIiVpm7YFbu5nKReN4H7D56
R2KzWBlXdbQQIXBJJPLDT3dHA8dmO6E9WvBk8Xeyy0OTTlIBTHJbvUWZr/hEvFpm
2wLL6byH4t8Brir120TKBvR+8iHkN1bt7U9dg3qfqYybYPVJRDqRMEeupZP8vWr6
L1TSnZw7ZMjN7qgxS4UYcAVZEDcVadCL3aEapgQct3duU09gK1njPY+NktA459P5
2gcdiUCQERM9JNMnjnpeOSJEDlZRX6QYrI7bqTsgLaoxw/sO9lM/MhEineRFFFkb
bZE9mlCrOsywO2xrGemuaJXPD5EpefA0lxmt90pJ4RQERghwDlCcYUlgSEZ7NsjG
tSzt9wNMhAi3I+PeRYxUhHtVIiQkkqqVcCncBQl1WxOyXHlZg2b9YLtsgyCvxKb5
penl6jPjdJNHGSnBQF911qQhCm/+hvW1GNbAxeFNaV9vbylF7QSYxDcrIzLmGtEO
CxE+oM7syLDA2K51PfasOJseSJkxR+O2NEtB7/3oqSOt4mtCNj5YNa4qUf24cCm5
++JEi6WuRa9E/6HdySwIWrUwsgAGNkXXU7QGPFQG/k/HlUjdDzb7otQXNRixjHF+
H7DntaIODFz/vHUrhf/d9mKLRj7Qs7YtRIDnnNk/q5T0kIj/mzcZYpiClKSuO9Cr
DbJcil7la5Ix3c83Iv1e5Nt5oTH9f9lAkEE8jNq3VjJlNy5cgzeUvthXrk0namUa
6ogp5/86AIUB1l7aiaf2vVp2LW7a8Iu+Mf5kxKwk/xVTmnWAyoea5LKNOLR8+vDE
0RYFvYECRHJDhbmybabP4SW7b8rafMnwb1/EvwIF1DXN91FvaphJY8hmIqSj2HKU
odnze8jut8hbRVj5DvaHtsN2yBOAlM9o1eaEe49NAbUR/UV16z0KgzyftmqoCMLz
cxFb0jWJijqPGb62rGDBtkUakPQwRXj8+x8iAaXc1tS6Lgnitt9QmllstuXaTENw
itb5YJWW3aYepv/cHsOSPtITa9WDkeGtJ3HDYzd90XPqUF/oBz9hcUzj03Ps96zg
zE57odARJAg55dYr17F97iC2gEZon0NsYNq4HNGc6xM1v7t+iXYNHgMq+2K3fZK8
hyJuQXx4AGbs2y5GPfnaIScL/riWEVOYsYZiJjafvglIFPGUOupymz5Xni2FKc+E
zi76W/C3lstDvGh8DmR02rZty2mozVtHwSXUupK0Yv+ZMoINknZFV9jW1Ux7gtLw
vDtYChAloT36lUPNVHSSpt7rep/uRZy0PS3uSgUFK2OJ3+MYduXBwZ2mM8yWTPyN
s5hn1CuZFGYO5Zl0Qpuq3dee+kaX45QSmyM8H0T7Nl6LkkiQmNLWM/KxB0y9pcko
z4NdUqAfu6RGfN8Sl0bnkalKOprRvfV8dRyx6uF0cKyLoRH7qoMypDXueZ2ZWdCf
zIVB7ExFwykyJ28lZSAknzZXTHlAN1lss7QNyuZAUpt48e7rV12vvS0H6JVKFRHE
Xieqs3OZij5BlqFyBKMKWh8stOyH+Q2ms9ZNTIzckeK5/zonsx1wnmRoiuT6vP+Z
pGNZoQ2n6aauNncx9u+HSmr7p4xDWxDBg9EadtE16gE/j6+1Hgn83UZ95Yv9vIdm
8oCbymnukmrCR04xxlCITSWZud5TFXdSFQ+RDFtlnP9u5moWcCzdCCVmQ6fN5g2B
v8D78pexxDNgqyWGAzNuldhyIInZmppaft2CVCAFzaJBeEX9MxfvOSSBMLmVG8hx
7uPhyLrfAhHGsNPOmtxb6hYRBJBt6DwGJ6RGfzDfkWwh17pAoBrLKVWdb/bFUjOi
wdbSGHo6N+gxvUx6JcdrIwfVMz0dULbXMEaHAED0O22A4YIKj8I21qznz81Gnu8M
0dDE/uT+EfDF5oml8XUFuD+iDHHzme5xr8tcHM8D+2HDFyIQETAJqNbqwOd4Nmne
Gkju/j+RgFFjBVUMVpgTBjSg124d9xJrt3J4VpE2vxpoCBE7MMOS6p9rvjYzoA3v
GaCR6bfJQueUruoPJxRT9J8R+L/goAAVGN0gX4DqF4rNWZ9ThnyevL3ROHHk4Qpi
byEkvDHqJ4kgmd1cnRr4tWMJKsBgcY2VZQU+8S113r8FzoNKje+o4zfPdI2Ad2uB
U0aUC3jo+hlQ3lrmvSeeQhs7fL9f+NqBeInibHdsstkvx53mIhOyWSJB1mowV1m8
agTTZQWNPL9krgVsMR9hw1WWqccpOSyZ5segcRQqzbZ4cmvat3fBjKF+N8L0ujxG
anSoSwxD8GsQW3xGVAXZELN1heylZ84aVqQ7d6IMjyA6kCqq4Q7zBxzeguExqrq7
0z//XvPyRWtHMVmIbtwBB9WidVWyMqqOkFMZgDal/hIHZYsVoZwhgbF5tKyxG2DC
uCM0c3E0EEYcwpk5PH3l0www/QI2JeN37dq1AeSRBU81wtwFQGE9SoSSVuVZ/Qof
lH+jvJP6V9KRmA9nZ2xniGhkqCm7mre8Lz/f98bxE0h5qE8J5m+6JVwDc4gKOURu
GEVrmztxlowQ5Rz+LQs7UfpDRVKf+mwUqqUwZBaM0WyO6lC9XoBQR6g5p+CuWreS
2w8J0nizWqzRNlzCZQCb06XHOCJtOCd0Ic2GlxKltbAodcR4ttPzpfemgxLCrgzo
Tebn7JTz76PJW/tFbJXins5keo/9KG/NYcGlC3bAJM4+KUaGS70p3TCCv0dNI8dr
hvfuvGR9kO/hEGG3LtxuI5Cqrh9Llvlrg2ZUhnd6u5bWrUGC9f3/VmQ2rzONR++Q
OHpBWo6y7NCJiAU17IoKzEHdmrYwmfkiZAuCr4SK4GCnLldHjzJlwTzBgsWoNdRD
zh7HJulGX0C1lbq5VFN4WOl1i25UNGrzwGrXFtdC2sVwpxJrbhvYNhly5wnvYVyU
KhIXhZDjZhkdaUw7mdGAZvp6uwEObew8Q6A4GWyiSOCDUs9nkal6vA725AupiCMs
xOfHx/pJf592TG7H0P5AdvPvYs2ATB0M9OCYkJz2y9NaxdEE6W2IKm282cS723Ql
vZ/Q5Hlyhl8KdLuaB5UW4RFmX8ExyN9iA/bgtq0rHX65+2l8nAbw//Q5MlkcSjf0
Uw+i76/li9gXAmTZFl07wUz4FayalRem7UW3ZSY2vPIe4A9oVEqzFo0679KiX/Ll
Npx6VGkpdt76TYzx2tP1A47VC0MONU62rRNjYN4/eseAvd/FazvJ3C1jZWtznrHR
PI0sbdvrWrZZz+V0ebaqdJHFpes7nAv2YXxLU8DXdPHX0ckVegfhpfXygTV3R3+N
Hs6d3fKigUeXWRqumhBfEZeJ0zeYNQ5bx/acg5vvzSAJYxOfgTe4WxTMIPW4HbMz
hK2A8nOtbdQOere16eX9zMdlITCTVrqzM1aPNYA726urO4v9Z8O+TdUSZ2zPg47y
y3jQWeQvB0VsPZlr8tDnBf5aHlIYo/51NJzefPVszVIOz2fwFdp2pG5N3vV6hKGl
44/Wn/LdkNr4t82NHfVPBuyFsj08cf3Qx1N+Wf6LOblAZ182o8F0TNh7zvhv0iPc
Y9sKe07absadDgQVDf2afWSrq9sceDTk51lkTYFSecPc9tKbyI/wXkAnx8xbv5eR
m3KH5tOvRNQoHvDGfTJX75hENB0Nags+X698hSuw1cYTA005n+MqluJRlMqh55Px
SCQIlysKKkxZHR20IqzQxGGhmQ83urrrDKT3P9U0+wa0Jv4JvwfSq8UFM/VMX4fN
Ko1l8Lf2fampB3aT3dzXUuUD9s7544dvV1KYdaRbvgQG/11AKQWJrKBayK8AvOK2
RNwTIP7VJFEX1GjuZg2VRR5iEFm/tqkjhmEmsJ82wTjLf5/ehS+fKADQRq3mrCtg
PncWNT+oY3H/NiTuvuzqahd+FMHJ2Es1huBqoA5uarjqqJeAcfOw76EaAJ6MdvCd
RB4VfwZhqShN9c8Jvqcmj1owgMpNMxs+Y6kyHSKTYt334xa681A4hsjOKaDhWPPj
uxke4ZnYtZHKLk6OjeHZXfftSV6nvYEiBfPFxn3r1HGiDH2T8jX8DGn2Z9Ziw5H6
j7J90+rnfln4W0MQNyhmA9S4PO4Ibdmbt4HnCd6lDPAwXkb/798bGuzguBw4QMv7
rH4mL0yyKYZhD0fvr29Im1xmaB5Kk7TqkMNSxOdNyxbIj8sbxAUha/2m5jOXr4aE
7lxEZw5nFkAcvlKuvJGx/PIsrviguU2pbgqTMS24oVSNpMSbrmzphRauxpC9iWij
65rmBOPdDTZfo3x9apXxy/zmEUlCbv4E78HPlSk42G9U9lTORzhK5bz8ZYl3K4wM
d8TEHUxCHVYCetkuAhit38w5spqQu9FuZRHvMfaga9lXYlrA2BhXeIMkECD6G7gG
hKw82tjlAiF6AvmQ/wWoaOnEYLeVWTEyjOi7JgHaE1Ba+G2e4D8wFWSLsEjIiRkU
eaFgTlJjInyQdG1/+9z78hB+KYcfRmJ7OEDnl8ucItO5JYWvoE1oz28o3UWiMFbR
DGji10w/A2yZbKxco/70XjIl3lYyKB/CI7OLCLY8lI0VNwvkz7x0/kv7pCsQ9oYz
zBF+/pVKlI4B22oS9j53V+NLVI2f26XvLS5bs4HGnpLx3XbtH/GKp/3yZgEP0vQS
wlO1IBy5iOMrM9mo1jszmsegqxcU3HMLgfO4Qx0qwaYigwranBGVbiUunOs5zzo5
AyJLAqV7JdYG8ORVYVkSgi8ubaeqAh432MU/lCSag5vKniyK39lAb6wbDTiK1oi4
nvPjKsaLCySSrP98GP+HBh2qFkExf66e/SeYGjsDDf4p5WaeeuojIIU+y/uaF39F
zjdrA97D4mxgOTJEwPprYvAkVBCEUa2175JrYnmQGuuEPYPEpPF1kbMP1fo5Y8OX
aYo5xM/RwNeE2DPd7kjZvskAWMMj5gPlZNu4JEZ51nXeugykaD5VgLlRteNuIlof
PFQ3NfvE+0q3aNp0elVlknWudxavNGRtYkL26zxDqyFOyUbw2cXu56qZ3rp2a/YZ
kPn47ScTYd0yE+/y6G7yIPKF6DOyPmtzX6CJDwAmWHWagsNJzESrFnDUTYaKSp70
Pbwq0LSg6eG0PDhhO8NqJLR8EjgO3o3yZbuoLwiKeNX1V6hJLtt8zo742uhA1GSz
GrLq43nZZ8hpkel+1F87UR+0MqKOXGgjr/F+bhgQnD4bRZOtH3OUSO880MlfA77j
LwqLDOwDf2eRilBgWFe+wcLL9Gt57K/ApAwrZof47FmGh10rTaXZYWXu9vnGmXV6
4iwtoy/WKCmsJCCwPjaiKyzVUAXqmrIt6kQqkAJhsTHoNsiezS18qBGy7xV7A55H
XyRZQocd+vzH/gXU3D8Zck8kqTMWqM17ZaIPxoHBwVoBiudQEkqc4hy4oFxrfpGt
iA6sIL3DMyS8mdzC63SYnbo4o4nyiew59CdpfZJOOUjOML3twauT0FA1cqb7Pi9W
ulaMlrl0PrM/IxavZOrSZ2MT2ybN6V352y2rZu8ATRINTnLW9jU5mzjGO2RQYSTn
qQMhGP2YIa1D//3S1dfs9YerD7hrxTPwJpEHAs8Aeefn+KnQfmhlDGIOlTh+LFFT
iSHnpAzh87XB72pF8Go/NnDGFi+kR2jfn7K4jNz7U93IfyeOq99n0Q/r57iRf+Fo
CRGc82CVHHpFC524VvvWG+km6q18iOvHgehg+m2MFauc5J6LR29yiPY7krThzX0X
QI+8/7PeNJNtu6eJ3HOu8FOTuNEwv7O5jEkNGavN0Mpgrkn0BE6pTPtJU6iLVHSi
0ZNtWcc8aIKLXzyWpnbes9gCYQtcejkdx+ICx2W3vT5U30xNqQrh7JQspQ6bDprN
j/Vkk64vyW6h6VTLLlCikWCg8kIfZXULFnLq6+bqAgIKm6A86kVMi01Bz2ya9l2q
T+Y8dispk0XFhObrtoRc5KrZZKfERzrnlhGnH1LePGCEWevMiWwztH0kgu5/eQ2m
erSxuMPu9vqPm7M3QLthiQUgLfErf9cf25c9Lqzla2saf7Px6dLbMmESiMdZYiMV
RU6IvlW+xKQ+jgF4qJMFem77Qjn/FfWW4Z9VSjqprytnSoGGZjmIORZjztjdYSVj
OoQ3dGWU3N/H8l99UUg3QpNKxtmeUHHqb2NtA2P0fe99Vwbo7RUW9UmGP/XN8idN
XizTna/4KyQWo7jECCMXlgRCAPyIYdBClPDQZp7121VXCf39Mk51GrHqijeQZSe/
JcbCmboUlruY/5J2RQ/XtdcLsNdX0GEMRz5tgeqKNZ8jyuM68Cg1HjY51JyNWCLm
33NWT+vjBfhKhqZwHbkUAR+FuCH8zw9ufwJ1pW9Lmj/grId9QlullXim1g+nFNwn
9PnNgqmIqoh/HeewoXDEMZu+uUmgW6do+sO0Rw0k036Tl2W57Mag/aBhYvX2C1fU
IQpfUZMWOBw4GACcfAu4Rfu/CCJyvhK89VlkeDa/YT6K2le+7oTGUolnlzmkHvE1
CwX+Tsihtlf8/OoJfTTSR7UWY8qyDy8VwyYtljqlUP/2hcpNFL1sWCM06VLBlsOl
8KsMw6Lbban6nNsmjFt/UE8i2y7j65ue172GLgpVvdyrEqF1tWboZYGD6jxBZB13
cU+Bg+CgNgxDnT37D74mkU87ORZX1IzrEB6jrnV4xDNDWx6bL6OQmbvBnKHjDYEE
jEg1h5YeGWaiSwun5RZWFdDEwfpVkQ3fuh/v3kP3mBolXIJ24lnIWSHE/YGpNgVi
JXIN77Vp7R3syWbyMKxNXFKQt+BQHxz1TP1qP0H4nl3Cd8Lt0Thp35qhyrQPSrZZ
cRkyWQpgl2ACwC3/Uhz0o0APp2uhAaG5GlwMmGPRzPZQiHh0A2Pw4DwkyuUYcHkc
hYF+Tczr5y2kESD1uV+M3yx5TSkp1J6Ay5Ju1zMUOhMkLoyZJm60WN+Oo8GMMISz
47qQbPTdxFT3H25jA4AnOkrMJOYFiR6RMg8AHAiwk66Y4zzmM+8OcuGs7XOLAr9J
w8zWaGqBi8bOCzRvDduwREQqLenaA4lwSYvrQY58Sjo4hUVvajtUZIwx1Gnbbd7Z
/6qptdeyrS02m3LpqTLRNyY5Q0k/ofgJeefbwZL9Cuz63WnJaX0Glf2nQ9/ReiWs
fFGIZKfYaCXe/uui6Qe+RKJOoneG/aoo8NWyAAinPiKUtquicGJse8fM7b4u/5au
YLfcBPg5ONug3nyt34JBFx0OLFzAT3Hzd4SY7wWSwL5LNoP0pADwkrFprP6BrHCu
Ywtou9G8s5ZsDE3IxyOIHDVSTQ2zI4R8JPl5Gz1kVk7j3QWz0C18Vz6nPRJsgMS5
JiWVcByJLH90XYK+vusny4dGyPaJmyVYF1Y8+0rsnvJR93tnlOpIFuF1m1RwGZ4K
omTHySGiap85XInkfVn5tLbuWmL3P4veMxgLuOO6DTyuXmk9nAhbMZbLdYoa4rwW
P9++Ph+RZxte8KkO7OQ9K8ybS2blDhk0f6S1mWf8I5K553ZoqnpSccW369uPYRLX
3XisRys/Ak29LlG8baCoScALqnYJ4POdbReYSbS7vORdLXhALrnR+eJiEvlke8qe
qjI7z43CYVLzfhgG6V0Z1Mpj+H+R10dTU4EhsVCQdd3+6HLlut8A5y8Gz8oSwEil
vIamDYwwcE6iNjGSCL6h11JKMMjKVjqlSuM3piq0hx9Kg4/mSz+4uNEn4ZUX4tEd
3hmVWODtQCHEM5ZTexEdZsXji9RI8IqmBr2otWBoN6CBtM0pM4FV+nK1VXL61IzC
1rZ9CBB34j51WoUnNQd5XIjz34tYSErDzn7ZeU5fcy8SEY3kOD3v7Uf7Idf+mG+A
Z6JjEMsls9vWkdfGVfvjG1ChlhfUBq6NkWY7qA+hZ2cG2VcdZN0EhwrsnGGFgS9h
hqCbcao//pn3EDTsWjxiVyq3i58QmxG9hSdZts3yhGRjYrmFIlH5+GRYiTJpL4PJ
Cl1PYvdVV2kfRlMDyovITeD9hp0VlxSZXSd3Y+YYrTruiFlARfif9FsrFmk+MTnN
7bR9QBXYMxMaJLTaTqcWSzRIXlRmPvMyYvjnRjemVuB97uzZ0GeDmtOZJdKoEt1Y
yKiZ0BNMQbqTX9sE6vcOYVzJRYXSFl2E3sq3rP08OSk8ptKzGj7+aJK2qmkNIQqd
anDCN6MWYXLrDHXyKdquG6ulc/eRFhvI+fEebB3PgdoCODK6llTd4qKJO0nk9Pz1
VP8gJCxzKNGL3olX+6wIW9m2k2WALrltopnJ6faZieG2Fn6f5hB4oH9MNgDOxVT4
DM6sm63fFUmOe39tX9TT2ja4METdwy1D8XLaVkw5HylXNsLrTWPV01Qxg8bWlA6C
ekkzApRRTiqO5j0UQ8xYhNW9TNmwrPhX06H9+WCoL2y+Hr+gJDOd5LuaBgVSMldn
95VZiPo2PijtbqdcR/yIXeao9BpPvmWRcuh34+HqnPnlClg8Ew1Kmm7hEHlQrrUB
tj1p4BivNosZq+p2tsa7Hj8ZbHWjMmGSimKBsPpITwjcCbPiJHyvZrRhC/wRHQcN
UWsf6ZCelVcP5Z4FC/yzbI+c5DYxqAE+AhWtpgXRe6FISo9i8V9rsXJ56tF8NKZC
KCbwj4GPPRBoqxw4gmlunwyjyPHhnlMlo4lNZTLV/5nE1DXQUKIaTVyA3YsyzFdO
vmxUIOaWDQpzZBYR5DLXHIOMRONhYzcLOHPqHN5xYu1g9EB0S2Znjsqt6P6CUyu8
44dV01ZRSCrMBFs6dMUQ6De8H3XBPhOALW6LbL51HDZQElUGmjR0YCP7VIg5MEEz
B+dBcnSDFD8kiOVnvZj8kfABtYdre1pMMvgDWoyKzgare1hiK2SGbmakWGtUmwEO
bHnLqD6twGx5osxPSUETcfzybhZ8Fn3gaDhbvro8ZilgtdJfuEt1OUrCKYuNfiJy
Yjwmh0w/q4IDInpIVjNUL50SdO4mxz/BRBZgoJ/hbyzIBDLFx+Q9HewyfoOVFy93
u+Jc8CgtCzsqbWEI4Y+8l2odEbSfxKZLHG/X29U2QXaJK3A960kedEhbKbeB2Xns
lsWEcED2Lz6FqCvhaa+gGLgQ9RiUN8/t4jr5Szsqflfe0JGA7meif4euzi9kFkRJ
U8JjquQjPusCvI9ioqGTnyUv980ANBkjim+kqGPSgy/rs0ALknYmcJKz/eC5H56c
r8BX5INMXAMzTuCEOwQSzehiY7t5KuSkr1akCnhb4FePbYuX20zyLyEwfqgZFZ4r
hnMnJT0S348+8FaYXrk+Xq7zZoxEotRYukZCZNUhkjvyRfl3dvwVQYp09dVK9p32
LVYP2O8v+QP9zs3yqyftqnGZvnN0HS559fpFyA/AqQ9uE/0pLh+S2YaAsru5DZRi
pQYrXzwYioZ6Y7NH3LIorNU1aCSpsXbbubkOGIU9P6mzl475lpiXEZ+slwZVTl4g
DSODjdLCyVYYQW1Q14be7xMsLKrxJAUGl1Q6BK0072DjTGZnhE74GyzEMM39wvmK
KfOQBUn0rTNt8gQ8/zHIB/ZhlKgOPEX4iV/ZNjj1tOzRxHXbqa7tC8sfL4n7GESt
MQJfNUQzv27CUVSpFggUvae/7/tCamyNBBbExP99Q5n2OrDXesVMnZjjVGy8P3VF
QUQhLBZwqH8yj1d/g2WU/+nDazbOtvapcIf4igUxD0bValSyi6kFVZJ3ur0Gh9IB
nBi1k1dwCJ/mDwjmJQHn7gJTG3RWSdvghEebXcQot7/P6CJJz9RiTUEoZJlX+OuP
r96D3OmuhaVFF+t/2e7W44KnbOnFSze0/ctgT7PLbF4LUm2mGBoqA2hLNlf+mpUI
vbm/lPLnSUistQxuGOINbPb15IvpomxgA2jdnQVWRnH0Awf71yfu4qiz8gX5q8X9
Sb6JggLaPL+9diKGIp7m1Gbq+vG0KnjPDsDpTlgtblks1IRQK5v3MgZC3Fb+t91w
1uL5MoNZ2R4sgst2SC+z7p+9LmqCIaZGActi0/ObUzVPbPs/gqxw66GNm8lQ1fEh
43ZcfCXZT6mjwur5PpTmWLLTV7DQr4dXnMmrgdr+ND4m2ImdNdUdYncJUmpuE47Q
7im/uUKpTWRGn8gOiLwLErNyYQFN4kDoQMUvvx/ZnkaO+PYfRdLnt5/8cnd62iSs
1YXg8zPTS99YYkTb1F02Bp7AVtFgLC7kt2QGvU4OYF12Ym1TEuOGw1xF1ES3CyxI
OCokn9YsXHJ9jQwIJArzJ0g/jF/ksG5g1h5ZSKnexjUjDYqBqNeMTeR5ggA0r0QY
V6vJJFiaf9iXT70TIiMLFycyRiXCJnJbcyVydfGA1CeJChtZPkDU6FWlTkigd+5A
fJExn0h+zgaUsrCi51iInxWVZ0kcuFMrNyuuMVkHMEEVxTAuRhQZfEksaV18SrDf
mSM/5peVqrmKT9CwvjRZxlzO9xnS3XA+QRG2tX+k2zY1l/1pi3YWD5pqDUJC7La0
ZKYKvggcOzrhf88Nrx0hsXdF1cRyxIIUeCOGIZm2SMhirvY9sg1tHfhiGQvND/UF
WfXt7bFBjalL0ROZzNeXXGANFUW32/THanBWHmda4T+JwxW66BO4slkyYugVOHMp
j8ZHK6eD4mOtptkc4BnzTMcmYAScNh3rbeCTyFSJdyNRuMKzKp8iR6yjxgdnp11T
YgmGyxo6RLNdnijO1ItfeU5rrDDEbLTBFd2RdjH9kktm9pzgRdpwKGzH1E6wqkm2
qTMBL05izPklpdOG4dV20i6wadoF1Km4zQKJocSosQtRyl3hp1ooHLivlp9w7rWT
GZhUNcTmpHKU50sGjBrtY9qCCyumwT/swDGicPmmnpONK0AuUsh5HevVRpELmIKZ
ItHF1hmm94cJU0NrFgGdvpPkqJtYxzvPL3v+tB0MqYf8ESXxKOGpmYNx9aZE/djJ
ZjJs1tu4NdA2bf8NtZ/bX8b7A/Mw69nvYmZve/eOWuDJ199Jvdoutfl0ydUAA+ig
h05HO1UcGnwVJM2lhJm3wgR8CsLSj44GFaONpYB73J9EtFzAmI7tuxfARnqPO5Lp
F1PTdVfAvS/OwajRmN7W+Qrzi3I80VnlGTueV+pcr79CNA/eeeuoNkdAfQJbRO0H
F2wZ2m/YHhlW/N7+39D1X8+A16Crpc7v88Czpe6NqfV85b/rtNU5hcnh4l8yvE1P
GO6RjRLHzwEMsOecjztRwTOuYt5Fkd1N6DVCWTFrA5JrjrA1DyC7vlZMQ5h+B9DG
b+8btPSwvYtHIQCi8gI8KBGHcSaqqhqoW+B2ylVb/d4+Toa1ObW/SNrgqA6Lhy1C
CzkXBF2MJ/+ZfhT8bIJ/F/fqEGwIEpAxDBVBBoa25X8m4kROScezdLevkLAq7Wn1
JB0aX1qPatZJoFELFs3aL6qclVRJp63l0F9ZUfpB4fgAwBolwM2XR/YmTIs4KSC2
x2heVf7HF9+6ijbn3Wfhq/Pfnn1cvj/aUBmoncUv0QEsKb+XJPPzDiKpRNZAGXwz
e8rZN/qJ+YmiIe4khZtgCg4bYjntb6QQ+WXRNyD3cywtCPU/0TpqufRd6ot/HqUu
PJPSBMAFKn0VSZbc3+XSSP7OKOxTnKrnBwKGVbwCWOqrZSldIbVB3rjI4zjrbNjK
aeHG+6x4B0dadEk79NGDcTv46t1mfvgcibYRCEOmXo9FQ7K9d3CqM77KF3llWv6H
GeINSMy7ZUGU5YZyJchQKBAVVtu++FNyCMpVQZHyYB2RLaC03ZRXrwyqH1hsXAFt
PcP9si6T4n3KLa1FyWFqyrhXbp/cD9eNSSNknfSBcf4m099ighrIOGJCbiOFBfYk
DUuNFVBaWAM/D6XPTFQaBGz9bK2BH73d7SRN33vkwdPDDkhtdGKPwLxTE8y3opap
RtJ2YR24sVCqGOwxVJC5hGUpWS0WsXQr0JJIytzH4bhG8xsYYXV/FwDF3PxGqXHx
it/hToIeVMQOF5ZynwnQa+oQHntVwjp059vJ55MtCPg79KzhL71EBMo/8S8H+X8i
vOkRdy5bnO+rHykPu7aM5eNRuAQ141Nd+pGQtEKtGfjgHFV+7lS/DpHMyLLW6uGb
W3nyJ2c/3n0zKuq3+G1APERWeXtggXOA/S16u2PJL+t+Sadh+NPYR+BJ7Pq7aa1l
v5FrugMFnotJqvzVKvZCJWMsX/62rVM5qp0mzu9T+11kT0ZNrKA3wdBQ7Yn65Tpc
W4oCJOMybYh1aTmbLpJlaP8R2HMnQPH6kdVT73C9CmnWiKfeL2hhg8LKsM75Jtwn
9cbTPL5eVR8Dhd1aZ6vfrC7cC/OVK3DdXsSuxs0nT3MRHvqGrSPOgBSMcfqLZLHb
2HHHl0Brd2t6q6oiBotBOpP/9bAo53m74l7MHDrzzTfhtrxuQuxubG1KRJ+E0y4S
272Xo99D26uI3HSwGFRtbKzmMZoG/Ih2hJ1H63wdK9zEgiiRUFgjsmqE+LIzddEV
AG0mvi8bFHiJ6HNhkY1B/1M4C24Hyz2/uTjBxD2lezI0o3EjdyJ6ov2kqRo2N9qx
C0SnREM7/QZXjh2QklFWybASFmwjytJPQ5MN3Keqh15rUHCKbGLXV9sBw4p6Dq8V
NaSScCwGSbh51tDSWHbtopiNC4O+v9EdNH/08N8mAXaQI0R3Wa/FvKJf7/FUSFtr
qK37Jf7GxP5gkmJaokRZlWbwwHg32W4ITvTjAnxeNIrL+A8X5FhZVKen18KA6fmE
QNelFaEHeD9sjOtgJrMiqZU284/3YeTpXVRMHMnNJLzutdL0nk/iqEGAvRsL5g28
z32nqRAIclRpas12ur81fQVgGvVko65lgEdGJGhKA3lNCgQnuE7jlHh1WE3ORXlj
VnsqUsIQHVCWH9jRIeuBEQlvcV5V5agzsxesd1aLvxHxc6X0r6YHG/F7wYKJ91ZW
S81U6artF7nLwWLd1GhJ/GoQta5GgAVq8uby38Sk/ERq00V/FDPvbh9ezGO6bZbI
M/PoJepi6w3l5d6VHo1jA6P6TRABt4eL5vllFAcEHmQRVH7nOilZVTfZN8so9z8X
mzJtFPDmJTQZasGK3DB8WA7HzyPsyeZigneXzGU7jXuHq8FAxulDDejDbwWzJCSA
Ln0aea+bF1MyIUPzZDiQNFD/efFOzqnlDvfqD8qKs+0MyuvO6qxekr6OLN6LsaRs
Tkz0JfIYzW2P5ShANA9ASPYXF+Z063g4GRcNdGXOjtBg0fvVzTfskQ4FzH3bbB+M
ik0hgSbEjrY00jQTpfFDkas1SV7UDgY01HC5TA1sB3k2EP/j89m8o0ICdfCvSTx1
VWqbEazarff6qneY/jUZVOQMqYAujEIysBGMPGpZBDvnj+qami2IJTGU8SDvMNiE
/q2vfhIyi0E/Gp4CCc04cFdmLjsezsEw7U33htPP8osQgCeZenuESscwTYcriw+0
HCEvaTIVwBHr0FwgMPAEZsIQ/rkeoHoX26IF/gx60+mNwPJssL+XPyGU4Elv7oZK
zp+5bbcVQd0YpwtzIwViFrxd3l02ovVR/kkCVmsDrNOqueqWk+64qGXu255rYWgM
nQI9pNO+tsg8PF9NZI5mDCcYUZkQTixAEyGHeAtNtP6vqGrfBUiRrBJT1Ax0ukBu
t04jEp7lze0KQjVbj+jFvani7XKOBeRV4I28uXXQT/XkVxvPC1JKYwIO9TZxYMfO
95apHZedo+4KVwMVOvIZUvf4ExdOpnec656u6+RBSUQWl1xaBwhMkBo2DLpJiYJJ
vJQQ3XSH9Mu6ib1USd1Usj4qIF3VHe7AKRQGulto+yPXTl30XcIP2g7FO6l264NK
e8AjyMyLPLLf+MHY/7iNzMiGQepECx6+vNClcIFDobsiPlXeWgYSo5cQmPAoxpBu
d0hAoJsw1/d6XdTdHa8sLOH2ZJwvV/3O+hxvY/v+nXm2wP1ZwBlyVb5gAxvy7t8C
IyYt8SQq/ZfwDB7/pJdNiLKjWMwBFuRgHUDyNaE+9FGSUd9W7wNrlq7WMke5cEHw
qyNloWOBPjgTzqFekj+eOVLQ/3JaL/ViWgaSuc8scIBeBTVXVOfdjWOLrug8agKG
KznSXizimLJP4kJtLl0GXq7MtwR/X5neyhaxqsHPmRKxdM0drIwuUS9EpVhcC/wM
YI6r+99+D2shU8FYb+omartqPR+atrnpas6RMf4C/G8AkUpfY0QWbagTp98kPEAY
VT2Vhkei5KCoA/FDwKOFn5br5/2OWAU9wu45Ng8++hz9jUKLnliLj7Ox4gwQxWNe
MUY69cR+REi3wqhuGO093SDAuuXk+YYjAOStYGPYSvTBTH1iYRtk3vgkBOadwRlA
wjHLClA01Ww7Ihkng31ZVDMsddQp6Z9vNtCiS/FIaVAGERByHOM7lBYWeSztY5Xg
+fqBJsBp8quPK8mVr3+8NXl48Q4mln9M+zHy97+rYV2gftKTLzV56dH4rwW9ib8r
BmX5IyiDxDJ2pa5u/cxO2mktyf39KNyRhbQ+628WmWs3c2ckVj/VkRgww0DmgoHD
S0TTV7/+yPYb1R5NHF5N0VyD9wozMzan7EaqLDzTcT2K+NH6ZWisPfzxTfbGHoxY
fKAmeA9hGucv1DYB9y0mBVdyQsa2wOtXIOXb0PJhZRkV6zjqRw43+KJLyZ4E6klV
ktqyOZLyJqawe272IYYoDO72Wt53DAjF4oKgVjz2VKD2Yu+n0wea99CPcVLgxD41
N4z54VUFB21yZ3zvu6tUphN1TQS72jRbqm18ZTdtECBWZ5V6w+v0psJsC1FmIJ+H
kdC2soPfuXDjVSTfwl+Rw16+LnsYTwG3Wxe4BswqOyLGWONkwAMCrcQHhJKqv8cv
F4A1vu3BpDIB6HbkrKtG99rPtZJLUI5VrK1AZZNQw31vx6k3R3dvBQopGDdKjkLQ
ZorSixsyor2BuaGEqZo3gvcAz09v5Vzh+RHiUTufmTu6OeOv3w4TEJRltkKtS7JW
YS45ubjxY6QcfcC6GQjz0PtPmq2n0j6s6po4b//PzH93ZNKqFMyyldRHebQjedlN
fjyjjUSFqS9u8VZtNJ+VUQBusHvKgUdVKjZAEgVElZEMrRzYQlGVjRQUF1KeXwH0
FTkmk4nHTw1z+JT9v2EWdtbkGAIhtVmDpy4i8VXpgQrGZ1BrrYcsB2cWyjjfbUWL
5ZebP38VFrZhRvtG9otuLm5gqs6B7VIh9bsDtWSN4F7il2xfRMQ3FILktstGIF6r
+hozaX4FR356zEtmNERw1slIPYMsbvIE6dK0Gvf+em4HgQ60Vuj3R93DqFJNYTJK
kzv6/Ag4v4I8KZMPEvTQIKQcRMpdpNnWpfmTm/m/CmAmFo45paqXwJhUH3imuA7o
e000evnq6gTfoYE8Saoi1AisvxmV0SrJPA9J35EcLfh6PqSWCyl2GlMhFOfghxgU
FyZ/I9V/5lZs5kmy90+dDZyDNpvuCH90Cw6DCYDWRgzc3hET6gECGu3myK6CLy91
jG2hszU/n8zLve4O+OPdOIrMQ/V5eWkVG8CO0fo+Ua/1JyJLSDCL8GeFl8J38vq+
j6XN+uqsPUgvWKgMD0ZqqBxHTZk2USS2nSGzRjv3SPdRCH73tz6Y77KtTXEXxmP8
uYqMaYP1f24oN/NLchIhJSBxeWnvKkVJhBQzGDaLF/2g+jhkjtK8sycS+jIOR1k6
F68hfp9QRb1rrm8SFkJKKRwazWQ4msAPD7csgdwqJFgMNcf0pYB1QsmHOf5wk94S
teZdAe7OtvGhFDEYYtljIU9LbDRcfKTq4Feqt0vRusNqEYrBcn5P/WYjCd43xf/C
LenUa7gXVhs6VSvTV0zx0TeahwVjGgCkw2unoEAqXKbKLKyvr5o27GyDUvE1D8JL
54Ttj8HIP4wbFHY+MUBjbPTDXmd4dRJdG413awhqq/54DLEchvExz+P4WkXue/7Q
dYE+LJ8Ib7Eme/GrfNoLhITNM285Ta952btl3WlU0ahBKVyXVpbAq5nsw+oJo8/z
4VE03Yfjk7qqZiEDfM3fHLbPP7i0Xhivt+OTJXVkOL0+IiBR2/Beg2u8Cakn9uAf
/rn57hfZQ9PlXqy5XNGi7JBvVD56/dsS+Af7s3KlBdC4D2+95J4nDpL//EkwZqaw
h01uO5COodOD+7DMxybLcQBpc/nMe1qN4PbbYBVMAMVVhm64InMKTnjWam/Y55JQ
S0EmujBV7xMKq9I/Ktp905gN/1hfHzEsTaw2pN1zjtRgjaqwuQMLTWy/B9wKIjAF
DvyOqWR7kc3CqMkanSd0CbPYOSF8brBwu8To9nVTgAkYZe3rJNTOUH+uNyDG+4bD
iXPlX9ObBaH0jiVZ6DI0A6OEKsNRqVY3pNZcnkDJcKH7gIGForXHcY3dQ3rUXn2A
3lXbv7w7kVEJZFleYluzKeVHnsOKs1lRu84TypzFx664hTyC9q4H4ZG33cLrRAs5
zdEH79Ix2FxxuPqAlVFvTpoM17RTsC6Z7VvlGJeILJ+AYi+Svoha3KOVbC1M2y9s
v8hdDkwbdDASdPsSsDyJ2YRxu829i5qYVnxmUs8vy58xL7xz5ENYNLlqyPIbFxHj
8XjpVwmMjYLMwUmtQCn7dUvz3J7rl8XWWDoSo0k2mkE/ZGFtFTToPO6xOqJ1JIjQ
6trIC1mAX+sHJsqYAzH5MxgbnIT/4T1Ms06pDJWFR0ztVOw5zOEUK6gMpGZrYcXc
QoEaek1a0dkgYM4bLtOzkzkMWuVs7uMT6vHUhUlTl/s9aDAHroOHScodQy5BRjAA
5qjWqNdcly+oUxmEc+VTca72iVkjt/AJaGYzgNUuAEOLtNuDECY8E8tMHphjuaMv
yk4kJYynNS+89ap7zz8KKyga38kWmJ3eL3Ks+HwGdf9jvSvJykUYQmUWlxpdmzCy
Lec9iXe/GSarWnw/TPbgPvyq/li6cJDcW9YRg6XaJW7AxrdSIfL8h7yRX2T/iiBX
9zmRfE7n4YWeXMWqSFgklWX9wxSjx6U1yGqkoAVgS6rVubvTJ6RUR0ZxeEFqzykP
7+7vukJMN0UsTcBXh2q1GwrpSPYkU1M0TYN2STP9s+KImx2HLWAj6lNBB0yDO2q1
WNDZKs1NGt8Yriw79HUA/Y2uyBDwuBmf5CAPyzf5VWLSVyyV5D8ub5y35eBcaYcD
uuTtJI10EJ/PdS4tI+kqpF748z354XtV9/qEUwJkBS030UIZBOYVlFqukSX0mjLc
vQwnMkczROZyKZjV0dQWq7ts2sq268gHSAO8LqW0JEE8VRXvsimn0yLGwRsJLvOh
+WBizRGVMu1RjZ9srQGsZXVpms5Ds4Z3RpV7RXnWpl1TcuIMusRgvYCga2lthDdc
t9kGAbyfMnXooP9eC7Y8MLk2L9tdusK5g5c7CnO8aBDhCyR45DTZoArTQQBT/Fnz
5SvklwdTxfayW3F/1b66qGClGcs2g+Z82z08o5iWXxUcUOHveBS9ZHRmYvnAFeir
lU6h8wWSC45zWkWhJAfh0205u/F0WsET9CZ63XCXK7PpfQWMVRG/ZMdgaY+T/1sC
+iRY2O+jXlq3ssYuZNnd0HinxJoQLYXLpxlbdqQ9rMlaoUDCO0SbhKeSaLYM2u1z
S1lZGrUmpTm64iGrA8/xGMjMBwR82wPwAF+pU6PWlWk2QekkSXTuEM70YSgPQiYu
Vb23E5fLCKiYqU58dcicfFvLG2mFpjm9Pzsxfk+WvhZJNNKhZizwp6JkI22U80Xa
s8qxOPxft39tQ8fE0/zpHD/IUlGI4KBsXqbJAbP7qOXOk8CytufPe1DtvHJJAeg4
HSomQaY553reXJE5vnkJJ8oB/Q1WESNgM1PuMzk4n0uELcU4UIivQvVBu1Ze59jx
s907zdezE7K3nyoeTVFchByq6yZTAVxOD1RjCNNmE8QLkajghZCRR8WGXUelP3yZ
9hrFoH8U4DYctsQvuIFLWfgdDj4jrL9cveaxYMIIVQahvIrX3mMyhItk++nBoAHJ
D/1dbCaDD0LvBA/LffKaihISTKnaD6fX1vw/kIzKLjRhvbyOwGRsLhGyAf1BJyco
qk/mj7c3vCvvL8Zy+G5AhifZcu8n41M5AGxtuCLCMMwfnzy4A5FQJ9lAzsixk1Wk
1N7FCQiYVhP57W6ejq/sK5yIPHcrliWK9orE87/yuMl7wKTpf4ViZ4upxrqWF/SH
KUZK8XuVZ47ymObexF9gP3g/wtfHnX8WeTLes4O1FbyxC2mXEW7k/Ix4E3to8IIt
HaqPKdulH0zjTz+/V09bfKNMVKQAJJ4Y13wDjdTPkmTrNi/N0uHTJQkn2W1m+xu7
sTp+ogDydT3jk/ps1D0jPXuXiKVIc7mct0P9rKSOMiaMu/iXtzT5H/7CeXSfFMbz
AdFlUde6dOnuJZ3CAvLOImjL85llOXzjwfAAuuE43Wk9Y5cnRr1W/49Jnrop2tBK
JXCyz5j9e1jwLVzL+FqlbX7gJ0dKyLJR5BAjC7tk528XGEkawlwM0PwmU6wOzpIu
505zrwOnHTh382FM0qrG6E7QcVhL1+qz6rdrNW75yIOFhmoXFoNZr4KIPz8TI6ep
BIt9h4Otl/QXaT1pTCqeh/575p2hntJoXo5rE+yB/9zXQ3PA7BEJ8H5HHqkCWdQv
S2ftL8iFvh8rvOvdUMVeYJVvsdHQ9skyFDUvGZi0veq1XcNl6YwfhrNJ5raqdJiU
oigEe9TxB/Eie1IEoRtULAh/JZ/0NHtw4IXkPwP7hciyMys3f0KkhTKOlLNuQC+C
C+Wa98r2LDedFGwmAnnpukK5mrvrLokBr4KtwHduT1FieCw5xsrZMS8qpLbgm2LA
fqZWoDh4yZ9C2TDI8mjlIxKbWwFvZ2vn09w/q8yUXfXWogyY5cKwB/zmDLymisoa
6/roe1OY5WS0La99dYNzxXsFg4yTIHqTiHY/1VCuIf6bzJploYkApuSvUuzbTJAD
tnwieP0kKP28qSnl/1xWOVxapUFunxTDkiahVpvT6UIFs7T/Y8VGEKVyA968vxid
ppBNkNimVQG1nFIw1j0mgLTGDumt4ArV2ouvYJvqNW6HJ5+VjyWyMZ/iV3F2cs5p
GGRTxiUkHjaPOeCmkU4BAxdFMDDAVUWp2xjtdZ4B7n7+Hwm72kVtLF+BeVFGbsS4
4BAfHXF4pWzInFuni2y+FhMTZqtn+AjKy8Qec0JQJQ+psgTcIkaMwWjT118iCwqU
hnAG4McKZrpPpCbFijO3kl3wr1YLrfEbQ3oqRZo7pBbVuOj2JBC3Zxy1BQrNMgz2
CxZuWWH0OzEg/sXvUu6yXTnmLgel6jNm3VPzpRPvQuWHCWlXcW7XsYvpGUxHzWr8
r2FMr8X4Vow7xNle3s3s/7nJqMtb/ghzdd68jIdrES+MFBrh2+0SVlS2brZqyueC
VUwGFMMb3nF+L40Ji2mB3yLIvtPpPC37DZvAzVcL5SiS1Sf9huzGAZsccDTF6Fxf
P42bATiUcluSjwiusYKOONQyBZLc8HCGCdnFmt2BF0LUj/Z8yyecFiuvNVBlgpXV
+Lq4+ZBBAYbH8vgMctdKYyTy8BNxxj+ZmyzcqaSm3MYED1XZOxQWwsjd3tlnaqhh
vXHeVgZjC2NGLtBaZplFLHW8FDT8bt/ga4gtOpuuGbJtE0rp3JvQqnc2ReutdCsZ
BN5dn2SHUHqOICLpNkjdB1d1i61CD1tbaEJ0AukRKZ+CAihrIuRMVXdxQQxtEJ7h
9K9vWl7oTWBaiWFvdFZvJVkf6cjuwschOfTui8NAYWMtQgo0HQ1rA2H27pEf1BR5
+5+ct18/9GeHqgIcN0rSc1xxhluP5TiDdtkLodvzIUpr+5V1L3CuDoj6iuNbUMBe
a4W4kaeqJ9lFErUb4HCfrRsrZp5ylP0gxz2KuDiN8OkUhYio0tDq8h3CfiEPH+SM
aVr1guKLr1hkhCGx5z7Y4agKviO+7b0DqODblD0qHDilvh2jj/vcA5vbDGJ1EeWX
fua2c0QSqBfM6unTrns5C7kWiepoVX06IgtN1jwwf1mHYEWBHGBp1cfKiYfq1hJr
PaZQ/0yexafYRZgl6X1/BMpkgtazWoCnlyijDoV17F4IFqva9J+iOw9o7qPxkMUR
VdUQF19XFD14EG6VyWxiFODmaAzawzzccUEciakJXPQpsPeDpdkIT6rO07/Eedya
SOexSUgUoytb3/qw1xILHtnLYBGTCLpazvB7MmOLJUJ2Gq7c/SlJzRsdmUybd0aM
TSj+zZRbMiLDB4Cg4zXwrJx8Jmf757IyL2Bsk5R+5fq4YKVW38HFycbtbON7KE6G
otoCKVgclwfHT0gQ7au9x5MdfxQUIKgqUd3jA9Fzs7lxEMeqrNdB5JObayfPOuk+
fOl9W2D9CS60quUyrO3sRZumv7pKnigDDxMnHUVx0jS50qoESkiI1U8W+Xw8MyQH
kNnPCZIm/Xvkw8pwYnWbNdTS62FdLknqn46Hck1itfIKzNi7ZKe5hbXbjJgGUWzi
Pg+FUYlEO3qeTR22bxR8jCw7pRve/LWrkvii5MUjzVi3x1fRLksEbb2jNtaPhrQc
vru6cj5heZ5uYD9ifNAS+PsZzC4dtAgaS1yiM/tJEzGQ81Mqa6+7GKdE3QpJfj7+
QiP8Lald1i3p/+A0fNGQ1hvFqKKgwfJqbHVJ/4Bk1PFnq5xwo2rl2Xesg+RanLEy
+d86SJ+0/G3HvWGcBLVTBS4NiFoswKeu9qarFyypKEJrkl6QmVeYCTMpLLDVIP1t
sUKt3FA4/o//NiCdPHtxOr0cqiRwAwZUZSZmmDAmS79U3fcidmVjPm6uB/c0NlR5
O0FrFhRKRn6UXUxtHFt/iXuiIG3nDOgUg0HSvlZiZOGMqYyscFoH5d/zz72o+2jm
0hUJ8vuABxKEXAUyS733lvyq7/VCurxicGzLQYkYY/7vf4JJ0wuz71+whSGEultN
rvHzTee/S0Kgl7wDBy90Fd+vdDdFREPfVcJ6poDN5xDHMSmyo0xnZGvwRCXksf5u
6pZ+K/l39vacd72Xj5lvee++7uRrtq6aBayMsMPo05t7OU5mNVZPtybPd535ZTeP
wPvPu8uy4JAzekxHCCZ9xez/Xp/NRsY0oMieYFuUAg/zRRv/BHlDn4q9n5qFrylT
I5SmIOx95C4TNlWr4Ux66p+OP70G+To/Mr4dPWzQTZM8mhjDvdqgIr24v4VsQryo
O3ioX156QnUCq1gdqEpDRRTvjanvmHv0D4sh/f92gMylqVVyUQzzicusLykn77i3
ydFdpWMZln7q3n00+ToJkQKlv41EU8WraIXkcNvfl+6vtmMHbdcQ6v9luSvnkisB
hwdu2qD1gXeUrqcGioC/lINTngfmk0TzaKhVLV4sGkGgeFUipJ1kAnC1/+2szhZj
irDEcteoKcKf5DDT8ga92pN+epxX/tYDydBIy6FyqOytZKT3swvLVovwVNQk6Tjv
al68U5U7U7g8nIdKVq1QUbDzoUvL9g9ifZcFM9wfY0b8E7GXvidMaOUJ3NUpTUbV
IdODx3M1oZhx86UWIwQ9gGy3Eyh8AVAfdE2Hrg2gF7GLq+/G5wQQleFEJm8T2as8
9FgLQgEnuA+TetIzYeCGaYlGqMkmt62eoaf8et7e0bpVLSf6DeEIX0yO+dwEW6FJ
qtIFCIvZa8/SDX1igI3qE+s1R/N+9Z2VRkl+4QCHEUHpIOYkToTnkjQ8n1D94CuU
POn36Qq292SfbCe+9f+4dmQ+jfqOZXniXwqNYzSsNDlRGLzSVzGlWHF8jT90+tcn
FXrINDOCS02gJnDgBNLxIwoMseZ2qeXKxCP0SUTsPYYQ/BJ4QAIK4GWNKLV5dll1
dCwDl2QQGRFeUZiuiQKpY+CkPfKQZQLyRssf6SOio808qJAE/wYTtaq2cbIM18o8
+W2ExfttUydiiu/XpBdUubOJ+kISX9dDC7x8n6Go7VtPqF2+NjCZeBmWyCeWBTJl
4/+y6+49Om/+r3BUIAeVbGTtLRPcDLPSSHA9xKZoqCupHFmlva1p73EDATXO3ooE
qc4yUdf69sQ5QUpSSuJhIVXRe7dXw9Wn7vBmSh07z0pQ1S9H6Yx5dJpFfiqqBcc0
7LifVt68gDa+JpbFkoGfstNvRhvyF+x+X9PQvwimS+Z/PaSjgmh3gu+EJrXK60fg
2aN45r61Ol4YFTIDWUeIaWyu+e727aFDvTUqLCNAtC435iqWZUwTbP7YYzWA+wC4
5MluUWw9DsgMEy/UbIfsSnCuHpKL4cIOObnZBdCmVF8JAJgm4Hi2NnyvYk3LzRPZ
gMnc/33hUF+Qu7+lDqxERAjL1g4iekHe8k3ESVawUR6QKJn+tBgMIAwHPFipBegn
79rQOLlHZp8qrx5qboewvKVn2B3w97IXOCk1A3TB8MNQt/dso588YMO6Htpsy4GK
HpWZfvTC70q9oJzLrj54S1DRdlg4eVdnO8HdUyJWjyJKYdKL6XKBk8lVJWVsBRg0
zaGtJzqz773rJnG1wHB6bhsRYAKLcfboBAvI6gGoqNVh+wKkAHsGcq3JdmVYTPBs
YpkFx0wER3gs2SAoa/fY9P9BIzHgIw/907+Dbk/i9FEuWWcV6CCd89DrcsTnszAe
FuD25kCk2JDnlCQU3VYKc0xLE/2uZQaoeLPghBfN+VTJ1SMIIfPO17AGPz3Z5jp8
IoRLCIUp+fqdlzVvGYFPNgTXXg9oYVi+OhI4b91xix96BnPXCTs631gFOfhna7Pw
vkcL8rDHbTaeMLd6xePtrC3i/JW2qZZ0hU/K1f1rdF1M0oobJiLKbp+xfqAhChUi
760Qc6+l4Wuz6UclCZntzAy2rLPEvsex+whl10OvO3waO+2ukH53Jv8EGvZuo8SK
OZS2X7+RzEvqZtSUX3JbxQlbA6zdoHqN+xO7exCS1YY45a53KLZR+RaobMpvCyBA
tdd+DVZu/47pREZFm50BHN26fq3ty+73K1FvHaLiVDSaR2YBKz7ycSDiJDsaN7y2
3u2R3Q9UcS1agASWPZbnmzarNv0H/bAug7x2GFTBzTDpq+c/xBUu/RVT/DsOXu0s
1k89T1OiyASWjh/H0ZrQyz+yl6trg9hJMXu5PDc7C3oSzdWMqyItzNxZQNCXb6SG
hSgUxpRpatI4cPqVmbZ9TpXh15MnfWZMRoRrJ/7MRtTxSICTJ9vGTOO5SbjUHV11
B2I7GtjlWkIUjw+kiaPhQ/3Wc3OlLgBSOEYJC2PXZPhVPsKlRDlY/UUzZOXiiYig
aUsABNV2/8xWsSOrzFSO1fHf2jwczMB2ClIi7+0W4nQ99F5U+5PwCqyRWxKChJRn
r+izlwgHZ7G+dPHqlDgydDOtJlbJUO8lT/RwPZDIGjtKc0DOeFTuhT7HKlpT4cAn
2DXsmK+P7wakgtJNqmmuS09sZzmqixk2jUuvP381MxbtyI/ITR85c4kGyeqCGCfp
YYE5EaMF924pgEzot+pFbnPL+KS1PnAzrW2L1PuQoI9Y2/uvDOHc2gsTc/tryNSn
WR22GI/GsX5DViI+bn77vyLLCo8llfJLwwtcgIkJ8qdo0OPvbmPcmfd1FKI5HqXD
FtQvWnyTcUPXHYOqZJLGkabMqqWXTFLjJQ3aRb0vFzyIBgL7MCnH+NedusoIxCq0
fnlQ1ljA1Q6nxZqB8Wy8NeFt7T8YxKy+nLU0NeSa+k3ohdkoqDCuFoXMyAY5PkiC
5Dn5tEwQADbf0RnpIqy9mqo3HQilyw4qs1oRN8VJ5zgmvJRVUqg/2lBaD/uIW3gb
2E/UshSlJ3L99RyFyqUAj7y2Gsa8Y0PzfKeYtYPR2NWf4DmhH3r9vfCC7JinmS5z
8LhpoXnQii/YyDECjSWab8iAKZAK3ojsOGS9BaStjhe1xd7yRsT4Qe894DuppSsk
/2z2QUG7Atu/GT/dmYb+XvjvBZ5gTf4WQR+N6zKL1eEraS2PUvny7RLI5wdAN/dl
EaFiSiSebbtrUgaOIH6aqoDHyNyFVcfwolFhLh51a3e79yaBJh4LXb/ItyDYeONr
Emx39IVzHwnNO3eFaO1Fc7H/ltMhYFvJooau2Zxkcty+aILeG0Yn8wxaq23oh9UR
WP9ZBxl+9uFksOVWRMaNPUFLDbnUlxLdCU07v7obHMFo327VQ/CELSYeze82SUXg
8R/lyBO+vSf59zvhLXSt+hMk2ZqwMYehlG5wZZBOkjVw6ur13sIBMetACs30jGtl
o80st/lcs6x3sjEMX/yzFkL32zc57caAzwYYGm+sQMvJnjJBE9W3Ah0MoNctpLsW
iackm8NC7NctcITUtiK1+DxGDwEd9sLgb2J5v5KS9KMKFTV7/LnXtWZy8CD49Dp5
4I+IfUWGZX1pymYnDGVadd3b/GGbmbxJfbbZP/lui1V7FAoLSpMJfUbYfFFgx628
u3f5kt/tzaVB8aBBI9NiOXNYLWsQMzVD9inJn2dvJuMC4eHnql6uu5Tcgb2SMnXg
CmrHdqGzcWUU7hsO42J5oEKeNyBE/4NMB0ayNMHd+/qtv+eH2V8XjyEs2oPNVSaK
Ibs5hG6Y0YcKX3ahUStl2e7tRM3JWh0Z/BHWWWLTLP6oUM8AYLKnZ+iSlYtIUVwi
+6OzHwROk3nIlMJqGPKHAyj9nAs3sbnLP/dONA+GYGTVPhdgr/80vNGsVKRXAjec
MvggB8JeaUoAjlIH4OuU9UGc1u28/REeq6IgmcyRGosSlj8TNEViqMy9EYBPJaIl
5wg9fUb19QdIC0OJAi8HxLtoHy2uvjCIwn3AwUloOV4iRpUXMkK98NVdE+7JxsQD
NO7iH+cpu2RZx1aJCqlZXd5TqmzpKv5EpPD83ATZethCvaTQwX6PfsuVqTgnzpJ5
mnCQktKiqY2uQIO4oHE8XuaNjxSriRUFyFT1M8vqVFpGMvaaKlEAAJyJ6LSED+OU
HhSewrPwcb2ytK6vMZZ+TaeyQayVU0CzNLUdZI4nyFY6CjIYyFLGQ2e6/ltOKBS7
Mlu8YjBCwcGqDqMae9MocHGzpyvud8DwhV/MvFk5RVxz1dzJFcox8EHFyzpM06H+
7rC8YWUuiN4gMhVTX1wQjKv3Q/Q80nVJbTwOeJzkkdFXACN6llwGhZXRTYo1qssO
wNidsfl6zIfKFarnDjrUpVTIA2kZFnKZd/7jKzh47b68KARk7Ywud31JsW0ZiPT2
VE/I/lA5HZDqpeY6g6B9K1AkLv8H4HFBbKhXO102ATXvjISHmtVfyLTQXM34WOjh
WvI/WL94MvCVmX+hX95b7e/vLH6GngS2uOeXlxi6nyj3i9upYvTpLufPGvJoDs5Q
7NXOD174rN0KOypm2FcFOT/jWyYWdqDQc8jWVSgSchQI08V+yj8GK+5vJUVDKD0v
yHNYaitFKQo8OTFFgrutUzb/G02sLe8v36zjjuy9MMiAe5lSfUvKBbp8Jxa4gIeY
J+kkLccbW0IwDADYCQIPsDd4OX8VSAXzg7d6pqOcckmt57BawlKH2bWed8W7cXLh
GeY9GtkKERnU5NPJ5GlPfJRGHsDWdvaa+ReLEKHJj5+J0PyhJ4w0o5ZzaUFglo6G
Qh+JAvJl0NILtSClGa/CaOVuCwhGIgIj97O+yBl4EFTnGDvpmEb9Y/4ZW7WhtChA
j4Iqp0MILwf1AMAYeo0BdkAxsgIiYGe9bQNZECFoQN5jWrMFZyH3d6NCg+K4+E3c
aPQe9BZwvcj9RdjGBbXNTfx/U077vly2dODRwR+nPzomKsr+LcHDL9ehsuy3g3Lg
/bbm8YOot97+/9oalPCb8hxOdrPNrJNm0SaePcjoUhdbxa2c3QLvMniR6a13IwF7
nTWQTUbyll0oZkJIECaqkQlqCty2hAXZAocY9sGMsuhUty8/0FnJzH/8eKXnCDi8
gzhPwfcLNOuUpof1o+DkU74UIlWvvUgFg4Z2vtgLjlWrri6EYlrhycgH7Hpf2nmL
99FMhu06KvGsRqODO/59QpSI8yB/ohpfUO0Gf3MK8W013TuDSRKQL8EpNCLQN4Vz
Hb9MAutueSDimQcdPzNwrfPOmljfXQKuJvihJzXMaO0e/xkcpTBsGGONEudwylSX
QIhrr11A8xbnkJtg1M3Zg7Nia/dTBsJW+cBYUZl7+IRqHNNL7pCX6E6wyDMcl9L4
W7f0BhYu9XSsIySxk2X9xZTYhiEOV/NFNahu1iN2KmJK68RNAVdrMVCaIEL6Xj5W
u+uAvVFUy9h4DZ6EBmAi+s5ZdwQ3UBb9pnJcOt5rN1ayiM0bguUDocuJIn8gQBwS
1ahDlkBoP/f1pVEa5Ey1nMC6aDXsiVmgV/465KmfISLOCkGOq8KdlJHswJ5lQfBd
2SPpg6MZeJakrGnQOlGQSdJOFlIf23Q9mwf0kPV1sPDl85li/Q38BR3J7sU2ZObQ
f7n2XahFyl8cUzrE4RydxFyNDXkkIAUmo/x0PGSnfgu3uLCpgjWIGrKg1qgbFewb
JOwyBo+4KxUUKu6SY2iTlc+rSlBaK5lcA8cPU0SZ6FGlRf1G+aIrdGroNXQUDZr8
12zuSGKCZ8xwcJN2I8OUS8giyFQ6RFctF4UZNc4vz9+CLLxc/WsMSEMMgZRcfYBS
xmjyHIbmBFRA5kAqr3QlwcVR+JzU4j6/p7pGCqCNBbYhAKP0S/Q8qH3icvxi8Oxo
3QTAMkK1yWY4ss1QeMp8fEkUm/P+ADO7y+XGT6mc1thQSHAnrbWATjcjGjXC5swl
Vsl7CyPB9zrQbYg0AhZtBNhTuYza2rtAOR27M6n5wTwQyGw8OatFGc8IN9eWdcwv
kFFHMsgqEOyBbQm+uZnAx7/in60XRHffJ19/TCKU/OvtUJpzKmbP9D8d7oAy6nH7
UCv67T92Vsv9bYA0A0vT43jDhwgF02hJw6UURthi31KOYSn1AyzwuCTTkQBJvIOn
YphEVSm5TYOsxtfvhfVXPRizTLou3Cm097SQNzrITs/ncKkwZR1pVYeJKQcxcd3L
MzHWW5ofnPT1+obzE7U7rfTm+SOA6E27MvwKJ95y0L7lzsfE7GOYBKLjJOhOFzD7
tuBQlpPzUd0on1rcQX21Rqoms4FvsrPxe+amy0OpAZAd780qRwVGReW5zSU3KVLR
hbjoLE1Uxgy6xFbsC5An5aqvTidrqr87glYU2zAV8M9T3PwexHJsTm5LNg+f34Vf
wBcGsQdp/SNW9POLHchzLiY7suWDW2xe4SlvreALKtP96xR8qVpxEtpfqE3UQC/i
CHnX2FjXkN5b2jeF/toSrZQDT+rwQSXPB/TstE/LbWPosipDf3cRTjKl3ZzbF7rN
2MFmgHyyQbXrxYyOBwrWU/fWmSspZ6vZXEq9FO5w9vw55/+1k2ncXXwjnNRvp02t
uNDo0frCmefvPDhFon6n8aStu3IyUepOvO/gcWZDlvkKzrHrDhE3WHByuNPOrwsM
IF3ACo+EctwAz7PVSYYS6i3irNyr0lrQ3l90hwbxDEdjE2ftB1I/wP2nAQ+NLDW4
7h7QV6xwSAMWf6jHD727DvazkNZ4g48zJ0QcEtcjrxdx+2JiwD5aDViaPm2E9ZtT
YKw8x/4w6HFFQXUKi0/un1RMTqTS0kNGLn1amWA+IAhPeF3ZlovkrnLPnC3Vf8a7
9AUxR3+HN6jDHLmXWn0EwJqbFag3P+DT3YJcUvoCRM0XmtzKwX380v9MiaRYDyX+
uWRAMr2AqJmAMXXHhDBB3ezFOIV4pplKR+wBVVaY0n19ei2BMVF+91f0sR28xc2l
m1yDwOqLjlvbF6JPyJityxnUHNUWdi4DHRWwDJD+E+efLgeotJO3041C8e0p0qLj
o7j8ZTksIObSZV45DFPCXfJ3rfKVwSZ/eWcubMMIJCkPtiSok3o51atgIkmnkwQb
r9iaC5k3whBzoDt9Ei0U6vtxbqzku5mhD0X8YYtQQon4mSjvubqwB/CydmZlIz++
XxGtbLsYAcAdAZcl86OUHax4yZ8AG8sV3hW2H9pfOmy1z3l16roOPTLwxU//pZQp
f7GKo+PL4jiFlOSzyAtr18WsjYBsWrbNj/2d8yIcl7CTFtVvJMfpSFoG4Cvfy6lr
P+/j2a7NPUlMgEmC9EeCei/AGDtLPzZlmvh1RDjGPjSekReyk7Nj4nPB2SnxqJ5W
n2DqKs6kg8O+zhyB2Z+hB8BNr87OcWj5GV2aNbgxTwAFnqt3lA0yF3TLYdbHcm5w
PmbLp9aekRrKTGPcCQ6kRtYRVQydJadMCa5D9RZWF9jV5dn1ERH8kjNylqbecwIu
0Rfq7EJ+KJ34c4ozZS7l75EklczHRCM54C0BkgCc0h4iEGSGvNTm0nhVIdO2w1ge
eOPQXlqui6Nx6QpBAIqbtP8u8nXKBfMsvkc0VXLKVc2pdBuY9f+wxbG2o4Mah0D5
Q6t58Bzc6C46c9sb/Mw0pJH4/wrYUHqE/jOEOj8RweBEgxwiRGqEAhYGu7wYW9Bw
Nir9E471YR65qCAoUphp3Tc8/CX0GSIBfCIerDEsWfHmAzMETCVg5LbAPtcGnFEr
GgDO6OqN1PTI+IJo01mrKv0MSq7uuVTwdwz2hZUDvKVycwHJ8D7RGBuTqa5JG9vz
1BT5UqkZWj2Se10LH8y/lIetlBgIOwA3R7rPsKJ3VN+4wEWwJC1Zqla8KeYOUbgS
5czIrgUvqqr4AiMAJAFqG0FpjklSY1eL7EhWjuFcsD5VSabvZdvp9O3pTiCBt2l1
Rlvb5M+QDkkQGQSDTpNSn6CQHNZFefWwM8GN8lYb/ZUqyt6fkoCDIKavDrRbhaLV
Rm+1QwBEHrou81r5inElJffEI84cGTfubtN9C/HFHOWf5DmIzHjCpjQVoPb6jBqb
WyE74aCShYw0hLSFjh+IPluGmnN86YSurDP8bkfeM+WmKOMedoinQJp78u/0HodS
EFdkbH89nuyN3hl9WhmsS/AoRnYI7l9BewfAY90IyecKyPGL3zJ/NYXBT0YzA3RX
Xr06DLfyYDxDDRFbqyDoc6tNj5h25LSVtSqU3F5jx7slOKpPH8k4VLr2PZJLzIk5
0CAmKPnSDSUDTdjsIW+60vemNH3EOe4G35Lt0sgx03TxGmVQRj/veDEfceL6bUw5
aGYA47Mc/c2WRRW3t/ejrT74hcYZkM3X41x4J1T5xqSDBzL+bfYzoZP7naWapKxh
LEy7aKZ6kCgc0MjV7L8t6CWfWCsOO3PqY33O4YkcZQZOoY+2B3rQm+WtGCelHsMr
gwl7YXIhArLRoP/xlaLLHu3cjIW9ozBAHj8osYd0/bR0MQqthS+na60S2mvoHbR5
/R3IEtnbTL4hc3FGJP5n6LjCasReTgjbSHFhCvhTZeIvQfmCDggDbgPZpEug3BRX
iIkaF7hRGr3Llt21QtKCv7b+fVEunibdDttTB+jbX52lYi2/x1EJ92fHfvnz6q1Y
O8YwPF/geMOL7d6fLJG010kZA6Yp0de7MjYgjbXHrcEZBTYU7F10R67UNMDxslnQ
YrOf46FyewiNvdF3UipK13ozan9n/4Kf+eFCEhP9qBj8AQCFM0KAXMYm7omGqMRM
2BJKZkoXzyVoAF8+lgu2gQoIKGcqtZ3kLWsaNolD6GhIE62EYK+kHktrvmKJt0In
IkVicetwC0uYdUbYDe5m6FKQAq/pkQ+AlNoh/DIvJ8Tqwc4dmNn+wIdx8aqfAvF4
BoqgZmS+dd1pUc2GMEnyN7fDSVCuLHbq0in4nvHzYueTqQMmoCpdLnlIZStFpBCE
rXZr0RHWuJS5ZKda6a2L1hsWg0QIE9MYYL4bJB+RLC8nziLkJ5hwud++9YSqCp8Q
aKaOYyrcZTenOIKgcx8n6r8FDQgnRO4LbryfYHUJnAyyFo2vwIa+988tpjwkh4M9
J570BQnmI1jmDG43s+PhdSucfLwknNWcxzUJm+QEdmpLu5nelo3Qt+rJyVXCFpG4
aQB2wn+GecuMvt/KsmCz7nG8p5bA7ues6fQLuIPQ5RAc0aoIguz6QA/VmdqYDafv
dOBdSd1Dc8Kvmb3AKDDO/eQdMxFpxQI9hYFSARS2uTLua5hSRCbBnTANGUxBPsXR
YN76levmj+jW/EWNmp4g/mjYNxD0NlP6n0ZYsNPlw5Ewn358MIRoL3sODR78LFK6
OfM7HLVsxtLqoQX/XBIaI2D+6QGXjCJazYki4YSjJVcuN/S8oQ48EybnGDMM87bT
SdtoRFHCGsa71TspIFK7F5zfXcHg2+ZXHAsIu0IcMGOWpzaC1HRmobWpWK6Yd3jh
m1zMtV8y9V+Gc7UzKRw2yRX5Yi+Weaf5BC27QYI4TA6LZwAyJU83KroXzmNCo1jF
TofpLvxg0B+wJFwxqsmRjXEqpI1yrdYpvR3b/c0/G5uMdzQMr5+Oo9hWLXbUTIXv
EinD1u7DnCqdwgavpMhVWmhNS3iZnAKjNEbV36godV17F31fZddg7nlSwUcwelQd
ubHg2jPQVdytZC0Z/pOLERnEcv9fRUcyefsSDBA9nUuPGlyvIgy9Uu82SEw5ToXG
T3ygm9DIp/+cGgOfZnRpQMfL8u5aeMfUk7Br5kRI1c1+AJXOwuo1k1ry7F7gqtOS
lIY1XYuqR41l9Z334Z8q/mzyxgOeHzzJ4Ng0PO5yC/ug8nsuZrYhB2Fad0XtrrOL
ZC7WiFQQXv3jv+DEKIEj44HUE/kVncyxg0euFKzpV9bYr01wkVgIUer2VjlNiqso
Zud3CW4KIf0CcOp9Q9CE6ZLMi5IWtGEkfh54uqDxVnchePbn0fIls/9ZciHjsoOB
wZ4sUkoV+d25mL/rBa4z2cA8n8vxahj2/9x5OVpho/scfBNjrjsHu/BC8E5cGY59
TwjAe+lB1EMJEVrEfY5GR6cLB0CvSFSLSkcrI4Ccn3EusI1kIVyu67pegLz3vJb/
QI9wWxWY/lczH4J9JjkJVIy6IFdsBN7O3TIR2lKODQRbTLuyRcnQ1R6ByuToluu4
zISppX/fQXlCHga1nx/y2KgFhsPwYaHs3EpM5OGJJXtIWlyUohpjcsyNfKNuWXYS
Y6E0A8gfRI1J/L98eDJFwN8Lcz+yDgS7Bg2UUq03tR0QxhM8qrhsYtTpiIzcnpIJ
ndGD9NC1NHKw3kUNHRhVZ0nPk0w0WUheC5ZrpPc/WiE2VuopCdwr237ChA/D4hLy
80n23HmXBrYMb2Y8DHoMBCNNVPwQL378xThyyc8A/JhlU8l6OI/gsVlYQPUWRiCC
o0lNsmPMPs485guz6D6sIwm9ClU5cjEiC8y4z4LuUo4Et8QDscuuzoZVpWGVRXz5
izxt1O9ROnAl0UZ2uztMwJE9PkeXKykZ/+XAb7YprXBhDoq8gcckH7NS/xLJ+KpY
nO963hDuV+QTzUQzk1z2RO7Q6s6XDPb3XRULnnPn+3MCqN2t/lJqeciVgam6B7MV
mLhH0Ej71PuLprkFQMGLQGPGBqnUGdmRK0mjKO+VPNvj2duZtEJrhCdo00lRPjCW
wOBo72COQ1MaynYjRygicfFEsAhGt/bU1wUpAuMlU14gNaxIwRjNRDIbQUGXsnUF
7rSqMuLS7Kzu2MNalpRHB8Ig8wzXjcVeMbgeVrFR2dq15XBQo+XT9pnie20fryLS
JhfjRcoMHF08Xl4Ju5jxeH+fCYWvVTiqqP4K8hDIeZWrLSC2aKYNbBH1FLme3WH5
L7elvLvwAHmpzrGhXJS2ZWrxczn+B6ujzjV6TL/SlFD49Kzc2gLm3wbGQB6IgNU+
jjbNkz3FoGnSrciOSwzAkELahcAiklnEgyc4X+mLTRqh3d95tm8YnGVsakt2w+91
Y/dkkfpWUGHsgYxntIobl0aUJUtDpDts5L/72i/elI5ToZBqxlYdTgzKuUOdSaub
kw2NxTWF0S4TebbM87J/1BdGDNn5jrDUjIbmSxQo+E6wBSh03w2lOE3rlyYLIWrH
ToIlAAj3IrAh2rUbTZ54lPTyx8gFxMJMNodDmrOTUVmbU/0L969Rp/g6cQCCqGiJ
GnnN6waWR2dOLhnKNm4XM1QPhdnBNExnjH4NZZH2oZKuDI9Y+sH7b4BFPkgw1zkj
DWEdJqNJmMStlD4uhdQlQMC82BbTB+n+IZcrynfuQJ9brOy0Gueg+wUBkim/I5OY
GaX2TDMzIgWR/Jj39SlYOJAaJWj3zq9kiMXR57m7TBx6akf8ZV97y9z1nYCT1luE
4qXqY79qgSr6zqKDYzZ+Q8BJEP2s8CKWg2Y6Zn+OMF+FkrV07OR6h7/xx7lOJuC4
NeXMVTFYOEmcvwo9pA2nxvQ4ZYa77Yhmvj6nXKYDjp8K4SE0lZkVQAodGXQ4NtBB
GQH1L4aav3FHJfgN1sKC1bfoapUA2F7dWJf0AjmDjhalKNKibIvf/DPI04GCx+8X
j4VjS0899Zk4OlnFpVxtAu65aGQdRCuBengaOxDKOBuAY04LQryRY5Z9RaWD4ddA
8AKRzaI6uqO48bw1JwgY24e2gq4/wkV6o6WHGaR8mWRBus2p3s95drxQXERpG+MM
EblyxHPl79+4o5z5iT7M1c3gX/HRe+zgVruyhPtKRovKDoW/WTwUS0UOOKpjUUWR
0jh9nz8cxpLTbuAt8DRcPUT9E6k0CcT2N+oslLvDSpfC+jq00/V1mVQnZn0bgyUP
kLBVMxAQAeZok91ASp6Vcx37aa3xLivl4Cbl1ERP5poetSRjC2fGNYorZiNtIJn3
38jtYxebvwwFlQLRhN9U1cZGAyJE3FETED5qMBCNPNdIalbIknCfvwESl8zRxhAy
BvT4ELh5nHwO930cRoK7XhD3QBxxiEd4QfvfMsvrIf4g7O3KxGZFlDt24mQH0qj+
ZUOkhHTPN8FiiCj/AecbX0eGFmCwXBBZRx4LTInFkYG76gBBHFWxgaGfpln2Yews
4Ntt+k2N8UVdUq+ygsN/iv4DwQz6/PyohS0LN+ZhGo9EXcdqnJLhR4t3+/d4dmRz
dUp0f96+/pEil1Dt+PzfSTj9BXvnWC8s7ir+EOSErrdiAHJZONG9iZcMdc+Sd7dH
+yJm3M0D/4N8YZw7rQRRSll3p8HgQkXeKBrbY5Sqq5UbYSE5+17T+V8r2HP3GGSu
tNA8rMylweL3KTXWurMZsvbUs1gzIY6ThPo/+hziikwuDSGu9bzSG1YmYlOIPF5w
08Bbdndb/6NaivLp4GBN4eE9C08sPjs6zKaOWMuYQ1nmvbHAIGg5DroOSAvPsaQK
v/FA+J9kSF6tHyl3n4VZgEKdGj7G9le1fA7qprTMbgkEA0ARO2HfQH0YwWXrR5nY
wX8HykhA9Uk4JgsDDb+5AJ7Qc7THkkvD387MnrkP0B31BtjHz1Fm4wDQZZscUDu4
MOgpFkraBokFy2vpgjY+UsJIrVPPAEUKuJZqKaLQmb/rGaIE+SB2fI5ssAm/RP0O
VBP3Gk/cvZj3hZVa1NOJZfFo4ZApjj4b3UcT86cdBWA30ABrlZL3b7Wf5b6Vipy/
jWTcRTnRbpbfFO4/PNaoa0siUz1becC1+CxSFohQCiiy3gH3aQzXekwUlQH803CJ
4HxlKPit5w3IsmVCte+FsF9PUyb9KKbnpAKPxPDIUyoEKjhUHii93PGAlN6Pn06l
dWZZ6xLKdqKYrwy6ythI4/jp8BJ7RD+3U+mEMCn1VXO85iO7DPLPApbCEWdzD5AN
sdE8P3tcvnwsWcG9O2M3ojo7IvAh24T2KaSBP93rnuBuR7LDNc8cuKFq680cWdIv
CWqaKrtWFLTrtSSE4Lo6mqP5CC6M3+iTuhc0dG+s49gOem5jQxiAXMJAy3qosOOX
z9+jZj4cIUmCJcMDHoYYgc7x+HGbNtQUeEEq9AaZn6BhD1Bjemxkal/TUa0AZQX/
wdGpIlyvDMjq2jowXotK3jhic4ouo/DyGjsIcv45PUk1rRRCTXvVDSxD98b05lxc
4TBfCvNO0UZO/5ZLv72b6GW0CFQqyVqYpVUtaSrqwH+cKaVRYzYyFuzELVKW/WSE
zy8OR7+zylMPZXA23DaGVhTZSYtK67TGJrfXzDX82eAFZaGAr4MH4s88qGaLTajW
B0i77MRVrAen4QgP/4POFt68vAHS8h4lutGBj5RNWZpsVQQssTHZwV2JakJ0dvW0
uplQdvTvUyrlor10f59d+EXzLpS3Wi1bM5ei7gMSikOUDxeh2S63ILp2fIuyykLo
26DaESjmlD7qwjO6oiYYV3sBPfqhhBuO3sgA/NxrnwINOsZWT+7JFS4OqdDiHniE
4AmS5S9wapr/1F79HUZhiAi+X/ZYrWexZo7l+itMg/rTLVhkUxS5DL2QkFDUjUG+
8TTLDFUcLUnVFgLAxjdOgi9VguJY/zlJt2c3DATe0CKQSXLH3gYULLv3+gJhiPYZ
OLq2hcPTKlFWAAmhxzOCIYysObFUZMdfE5BCjU92BbWGkQo1i5Z67lGBf46jMFum
FoItnHoECx6LolK6fAyclvRu75sOM99nBSfGDsTY/tzGxAJwskncUJkxgOGQGW5x
fVC0m3m5QctOJeBfsj6XWSscQmSBd+6SDHem67rb2a5ZEWrLlFnHerc+IDjZPvPd
z/DOIWI7ZifTSbG70lk0hecV5oa5+yqiwE+V2YaNKeda+pWUF2yDEOFhgEnWFHOw
C1yoUS0x0xSSEN9wlr89R9AuWip8HfMZ7VEv+yYIuGIoxoN7ka5yokbdcMbHi/N4
aKZzREFfDuyHAdE+dZ72omdmoyHI30dN+fK2hePHLvZaD71GRNH4izOW3BuJWMUL
yEcymAbAIJPVJxbAPzXLdU5FqZ9Czz+cBkRA4k/DLLkrSy9Zka262xrYPsUsbPuZ
rX84rhncvTX3bsmLZP0VAKOBmgcjrGEoyas46s5kvkyc+jta9ODlNou1pc3F6u4t
dWTDylBolScbnWixIpJA2rYaHQ6MkdjvrJYJP+9qIdjmaZDGJDrqK5oNXMATTcJ5
7YLuwtrqU1WxlmkX7mj8okrYrMUHEGT1fXDzqJu9KYLBr9RBYfaPyhLW2x/pseuQ
iWgL3CtsgIu7Gd+H02o0JtgYlxsXcS2pMFSGGcD0MCBAzMk2/GmfrYPj9ybBOHrn
qxVC1i9bcIxpDFtuj5JTOc9ktvDRLU8ufMgeXLQF+0WrdJUZanIf2wNR7Fy9V0/4
9bavppobK1wMtCSIQSlZ8ZqlDJmaNi8hAY6fwpW07c+SP1HuSQOeT3e6odmmN1Md
DVbmvBS192AEN1DbNT1YLEE6IfM1ynuKwzrqCh7JS1q1ZdT4gnz1PR1pdAX25s8H
0IUWj9GNCYgQzCqGM0oUpDfzwslKQDGpQ5db8fJHH/cD2r0iFhFBS+vBX/c9OXqF
SwOFpi00c2CwUKYThTFU2/qTw5Hf45niIwAt6w9V/19PxcGA82CiUTvJ8lmChODZ
q6x6YUwp4dhtTMQq/Xwg13wdpXN110Mgn8KSB79JOsCERqxyCKw5APwEJfGZG5cJ
PTOQu4FdjTpHCYbxkttw6zS5yELtgV5TKVgFY7z1fo8jGC3FuLS7cISNJMxlc3zr
CogoarrPx0+Bu+iUieB/UnyMLkKptxhJlQMocHVpvmKKfje4Y8RcMc73UQR3ihMI
PQvbZQdi57YyyPlBwUdMzngx7R1EzOPsSzcRcWfQQ/c8QC17HurUIMFVF9bOsF+Y
3h4qZTR/wM2Gb1SQjW7/++vhqOwLs0+lY6tzq/5p1JRq3OZ5/jvCFp6KbuhhRx9c
qMieLa4YCDYd+TiP8z9LKUItz8ySUeNvyFO0QRishfGOWLXfqTU7VhvpSSkeXw+k
giGofKvNq57rBDB1rqtWxvPdSBKR8We+lo5YkbxxEKSWvdDX9OlKiKORTPj7+EP3
+Hhnaq9SwSF3WsezZVNtlQ+ZLBm9Qn53ns5Yfij2LgRoNQupZpgihdcPEvOP2qE7
nfg4yMPUPN+T4IIULvOyqAANHqyhTHwGtI3JuJB8B/VcYbTncCs6ht2s36R1XhTC
mzPGko5C3lW7iQHWE5izG/6A2nV9zsSu8e4ZAI8Sj4szZp/yjUqzLhX86V7Mch0T
Xu2DtTiSwskvlh369sAVHsT3qVx9Xm7wjQBmexfWpJy1eOKaOtSFmqnNnKCMIyfE
5axOHcaNV9Sm4GGsuelKfpNFbx6uDtW/jyZjT/X7c/WNPA4gwte6o/ZXeBCu+SXS
GQbSlzHY+dTuPN+ln5Ci6lwjOSAMT9kJ+nXdkjlRcpA5flkTVkDmHWd/q1VtmjSa
ONMEYvuSmXeQUW4kjQCMFTxcpYFMBUPl/JZBtzW8Bg6Maky8vdwbpP7E43wM2skP
COqDjKj7Am3qHJ7x1uMd/eLS7gHLj4Mhw7iFXrcojT91Yt+FW8Qgz9mkhiNm7vQm
ZwSXo9LBCTOxP7PcwjUPbq5rKwFjACU/vD65qzgtyPkpLHQ9EMBDFsy8Hr1BKSnU
2RoYkpop5BQcir05rmTmrgFOFJuKDUYho3EWgwyZqJ5jBdwohPTLt7PZHnS6KAIN
Eqhc7UcFFq7XnowlYdpBzKWBP8x3GzrrAjjm5rvCxxvQNd3USM42aLAeYg/wWFHY
GETc41nvy+UP1VftUACqfyNFDfX00aZgwMDEiwvE41XCqEli8ZIdpn5/xSXtAtss
IY66LI22EAS+2xljdhpDMK5MPqT5YGUbxAC5As/ohXI3OdBqmPAe+GREHR1U2IdF
n0RDeAIqxTeziq+C5EdxkkBazNymhFAFSlSYE5pDv1RTDIYNW4f9YFDAsu6PiJ2F
l6SswHjFvINmIBAZ3ryIPjELNMhC21zx5erm5VfV6gxvqL0+ULlBhyseU4E6Yujf
NdWZs/Zela26eWIYv6ztVo2Md48p9OK5QkzwwYAfnhG5bEpLIywk132yNar9v9Ut
ZIVl/OoocFDygqjyUWdeE0kdKJTbWfnPP42ojbcHAIAPJzieDswhfxG6c9Ty3Qmt
FUrMS+ZjWiERGGbprQU6VdOoFval9W28ywOMDarVW1S6rJyn2DniQy7tY3VARvbm
oRf5J6G1bigykc11HGYwpxvDaKEMO9cf+GexXjplAsVl80kXnilzIYT7Wa8KT9nU
7pcd7SV5e+T+aNSfDdYCzCkp186tPxiExyXe6s2wNfkVLGyYLzhmq9d35EHL33Ex
ksPorFMag/rTnDYaaoyL6rQrQ4qRJ0HiT5tkDS6lluJHpZvPe3WBk8KPfY9bI8dZ
ZJFK4kBfOFBlfePfG1bClRkdiZgGhoZC1sMIyPiyNIDEnDtmehpsgDJxH6SbSM38
dcDcYienx+I0bR4SPNPCqfEGTwCQGqpyUsPN4UeucrcSO8YDTL1FoHPJm2hg4sQc
0SgQhHdcKZFqitK677k6rstEqQwey4QyQ3MC4U4r1MpIgy/7x32pVfHLbUaMysxU
sftuVmwkWDs0A9diLX97fmPx8LQNgvfcuz6iAAYl7Czcub0hyiFpfSAgQAiGBjwt
dOsZLGUd78NUpvtAW5h8YqQzZHfYZ6SXmjrpp4h1juxiRP2ce2uevOBfB/hwdu/Y
9fONkK6ULkY1skBJLQ4UwtXo9lntHl/8WHJYKvhIsuOamcAGQTTPi25jcKoN54Y3
ymuTSyzOXPgH+e46lLrZ9438pEwqkN/YNzW/UyD+Kpab9zxbmdv3PIbTbgB8ae8F
l8vxEZ20zEQhM4XUwzJgxGMBSeLLTwUZfSOGm3hVgUIQzRo8US2iHxUbqFvzigKr
11T/pYLAXak4jpMfEhjiZVJV3hzpkenX7y69Hm3Qs8WUYHA9nebST2sx8JyrKrQD
NbJ1JB7IU4Do0BmYxDT3omepE7wF59qflciKZE1YUs9QxC033Zi1JJZES6huaKSu
GNDEhtf6QYzcq+ROO3CKL0D/hcaBDV3J3BJgYXSOUGTRyAIqP5OalQJevzhx/7h+
UztTdsIf0PtK0kzQ9NOVBPdDOAwh7pbEMljLjc41KB2eYxbXHaH6AEQe3Ezp9qWL
4mvB9hSQJGXzRp6FME3dOxKvfnVMSCcsrydd2QXm1JqraPDTYchtFgZWyP48yUyD
0m1xr/OdlEyhm7xEdccjdPPtM7bdABJmhkQuLewS879+fpM0xEX4d94yYiQ25Ium
CQWY/+QlpcQqiVwpko1diW2vBn/ovDlWKA8B97olT0q957nbBl8eWFsjhTYbmBRg
vMe8SHL3k0aTE6bYBaRSe3NyWnaGyf0PPg/iLE7Mqu7yk7q3RxPL3wlwX6qlPsue
/ZsMBSjBb6FJtR2AqUMO3mWSEbhL4RGztvZ9FLdxa22Us2hEiHT+k1UqnzwdgXx0
KTG1L4NlQ8t5zmPTd2i4ycH6PQXECtDWGcu96nZ630m4dK6Lviz0mkU96IXLHmgY
+2VL/443vF/B8SDWZcIFBO0u7oFdRND9tp+VxDiMI58q0pl7pfiHUi5TyyhT8xev
NlvOmptFms5n3MQ7yQp3YJe8OBLYLIMRdWP2f9t3ScL99gLX3bU9BKhNqljscTC5
/sg1G6JngXyUJtH1K5f7eXxp+HvDzI7cffSfVrA5tP40cFf8OZ9FJjb9lhl1Cpnd
hl9ygCJ55NzO9bkCQqtMbtHEqPgqT6tkLrEESdmuxBquiB2jQnp8ocEPGf1rhFtG
9QADTjJrtpOSNEwyx6deuy7q+e0oFYldydLMj/yc14PUYPDDhG8j1MZMYb/eDlUv
akirFeCgnydkayxwYBDjXA7dpF79yxFTqiui1RL+5S6HDHKlq4MLMmsJdLb6JECo
fUd1dCqZ//f9HLZhLFaPl7xKD9dwdXmtiFoaVIoNNc5jCm7s1zZtQEKbGoDvwoXr
RMbLf8FvKjD2IaH02UtEGqMf29yP/UXtuQ2slcV4QWskbJ65CoO06TxAjCpkG4WX
d4kkowvyQPDI8t6YUMnpyMn7k7hCYcqpQv72mu+7Z8fIssXvW187pVimiiy+uI5M
jhOD478aMTtZa47uAq75KNyNE7pboERtfsjd+6oK3QyWSdKfDcz2rHtrwp+OuMz8
JUwP4HZ8UUOmoqyaONCQWzpGUyU37v/lMpJgwMDWRf/gglUS2+nlYAMjkzDRhyFP
NDm6TTcuTYompFJqE5ppV4HAHJ2laDMgEDKn2BsnbyegvRCnFVgRVNDWJVnBjFkt
YLnQ2V842CJPp776qOfaXo8X29k3u00BKCKyDe85LoJqnocn4KUzIw+OPy5ppovf
z+CBjNdfuIWMeYFa9L8YBe9+IjcuJzoxPouFu3b23FLyPn2ghvy73L4GihvFAjKX
eoU//6sqZU6OJ9VhTqlsSGENRyeKHU95Juj3Kg8xuj85u4Jp/KMFA/+BWsGgjnAO
T08lbtcTEdslgp9NyminJ4NyKJHgdKihSLM1pXMSC432g9OMbNhenX1XSx3JKkC7
C8iOR5v8riQ5j6Oan0+wcfeM/jilwkPG3lGxZVRyWNEO/Rq6WgF7/LYtZoUX5CX2
aEWVvrKxRy7kYwu/RouYiFxtfC03NegCskBZLAZhr1R6SgI9l6UsKCAvAmV5vhYl
qrZFFo3Xa97xTOXlG7nAWO7OoXbGOLhyZDYGYzVmdGZoje6hsrkTp67t77kCJCpj
yKmN2p85ojtNz3bTHv2r3nc2NidJihwY35uGDhZfUXUNvqEsTT+XCEUAlvtFJRGZ
Tw7eck667WBrYsyC+Se/0AVpvN2Jg4+QuH8BewUGiNlfhPSetmnnCydHmueH9hON
OEouCFNTWkJlRg6XMVo3poHXu9uPrJ0D7sSI1chphbAm3JP67Wt4x3VfLfLusJ8q
FYPXaOP/OrSWoTJ0Kwd99yEJ8XNBOnxsXJDjkLMhQ7hX3RHPOQotkSOrqSlLQcxm
4i7d7x4vnr/dub31x4QNV2OZx/1qsQpDiMpqQR0UJvde5vgqiadeqtV2yyfORlKQ
LlcsECBFjGwNnDKuzxG6tWeAZnDLvdN6mwmn4IfVbXuStp72C3YTyaRm5YPuKsco
FrHrb58JxE1EOJHDD9u7dexPOhkHCrScradQeEsJjM2936Dg8TaR6gGV1sXs1f+/
dN99bbnyqlXh2sxmMaV8oyoH0Yu6yL7XDbONEe5H+M2unEX1S0FFF19Nz65UJUnD
nhkv+mtEkhZ68TkRu2z9m28nEj9x1PTepzVV6BeNXo7sz6IiH6V3AAIezqJEfrII
sMAqR+TjjV8oXtSR1x0bpPrFAXGepk3w7JgRRmmCpbDC5HuK8/06Rr57I2um7pU2
440wm5myJ8SwS5ECzo1JOW41LLK0vlhUQ3K084NdqxiZ996HUcuChUoU9CSlhWRi
tj4RmI1IuQ4NXWNS4I7LqCj1nxnIRMQJlBWnhtCDifbWKN0Be+EsyGU9HAXaXdsT
qvo2QXOdnQr+XFP8miDbjC/hi2sC5aXbfpBXLBg7NewIEyhP38mAluyXesXAwm3n
ESjev/qTOu7BxPYBAG4M6mluXlNp0QnSihmXiQjbZB36Ut1OAnxnEgwtvoqWiS4B
hnIeafZqw2RVNg03nFteOFAzf5oXzPjc0fmQKtwPJbdk1r4nMgXYWYLLeOe13eW/
fuS4ZzRmdLHlULmiGqO7BDwIERB26lldgahE3ywk/MpUuyuxQaxo1jJxMVYnYwLP
iq7ukhxu85HN4SHXjzpGhOiUuUw7Jd1Tq/cP5vNlccUfcEbtQxyvhxgXjziQNcwf
/5t67lvdNeC7ssGrlQF253jsTTd0t8v+lZxPbKGFtp9o5pIfwWFnmRAOAmJnq9lj
N5S6AVJ9IMMSjaJK8T3NCFZmaPBFekpB75BZlvKL8r/5HY2NN5R2hDw7PZHm0OlD
mtlFU1A7mmulJDt0zRIA9iq3QRu+ddIahSf27jI2QVAb0j7MO1CVc86brYS08Jid
r5faL+cnDKImGFwcBbcKn6gVNARvm0D0NquIw69l7O+TuZ28q8/oLNSc+udrdhpq
nATZwDAngVUi8nY2lawG2Gw6gAatJuBHHcLmGzaDLnB3l64iibJSihyXc6DCszVH
rmAwgsOoyzWpyzw/tFR+3JC+ONe/FMiQuGNIvjj5CoGqX0py3aXHAlMzzVbucYc0
xtSiKEjQ+Y+XVe0D2pdqKniel/OHHB4t2wIb5wWSBsL168bVl8VP5/64DcUp0RBs
lLxZ38tgZZ0dxJNWNZqhetV3zhVrDj/TALplWmtHh1QbqL0mNuZaV+0EyLN5IXvI
FPgDuYI7a89nZgUYbuycq75RPqN0n7Uon+GV/smfu0SadruINDCSjJhFoQAWZMfa
nEqNpV4Roo4PX1wYMr+fyfn2wWi69RUIgdfIul1WY6XhMFAuYP+LpLmBWar6axBD
SUxM/lVQ/c264WkXQOTLDbxcgwMVTqe2OPvouqlSYGEQyBWVoHLpju9W1bHZFODu
S770FG4rKznQrfAiweAS+OQiTJjoz8zyN9IJsuomcLhybaar8yjS7jsQLfrtP66j
0dxA9BjukRC0gaqqMWW6Ctk3RvbpCJPP1A094AxIF1ffImyUDVmJnn58Uw4ckdKk
bSwzxDM8YHLdetB4guZyVfX8Or/bVDKtPOIcx0XZ4stLXIN5GenQ7tlFLyUYYhW7
HsrMVj75+zjUTCqAU9XIa9q1ph3UhZlYB+/COki1/BYwhpBgFJcVCyOqjuTl0UvH
Y7Xu1C9h+SeSoxvHcJDMwm09wUVl2VlmenYloLbQVbTqE+LYXdkj6SjKetvOmujr
r+1x5rGDyNJ1YKf496C5jq6tNAd0yTnDoudcKIcVB965Bh4AuAARdAbLWgSYCmGZ
8oymfGleSAZYnHAB+a99dSyfPLCRoJH430TkBlQHNaLlXiIj/lEcvPzbvaAIzSAA
Bj30hNdbZengLJ9zvqaWsEd42S0sSNYMeWQlAWgG20a8dej8On9EPWt7fqzs2ngP
l7v+JknbhMcTT2u4PzU3zijs1ygQBc2+qoSsOoWtpttLdwHEnzf+ZNLUNYHLC464
XGTn95Kx6BVdpKJQ21y9Dha+wbjzpQEGyAt2y4rTTmArAk1BPL7VH1dIi6gGyWp9
BkqJHjF9fPuDlPRrdnMU/Q2yzK3DX1SUgq4NrC9ESWGtzATXTPiYR8heiq0RHQh6
LXkQWJoM1MGhj8BRoX48VNLElkz5fIiEbnCqkh/uQzMQ1faDYyx5ePdZmN3Pnkra
Q/7VGTKy83KJ3AYCBd7/RchzKFpRcvaw/uoOlAdch7wMe82VkG0hMtaClP01YYCy
X0XIG0ugW9i59Zao5IxzvGufL9HJ/g+x+aehYG8y8RPZFR0b2RBOlfVokx8/0hmX
Z2mLJhMHJEbodJIPYaH+6EExUthXYS1tAeXTLgUbhKpdzDTPoQAXQ7t9ghtneByh
wFa0Xbfb/0KNpn0jnEiwLeUDN8/VijxbIX+3pSChyTdWHpXK1nsces66gF5lnRbH
tnOtieiHOpKskO4u0/LbwSzveC3Ze/7o4cGbdYxNa7bf2J4Qf5ZpmtT3sDFUOmnv
wX+YeViggqnRK7u1dKmfU4z2M6L8JXxsn9iQzu4v7Waf44s/bbeAudBGRGtmHJ1t
UyVgRKhav8N1Gq14uUQrdHf+wdMS7KMKKytuaNIpyv89L1HuGaCKQanWYA2UXNhP
i5xOjzSxaygoQPvxAgbRFWoVIHJ4OThNw1xPd4gDx8v0NODYmgYpQl/zirhT92vt
7976uvVtl7Y9/HBgQ0/poAkr+PCGUm2LSf6q6BeKSMGWxhC9UYd1U8gKtzIhr7zE
x0Wbg6fY5eE4sGziLCTdYUIkMF/EN0vMs3IQgf4dXcWbrflO7bm1KIZAN7cSIYoG
4qy4u5Z004rz4Uh/JLmwamKKy8WNGvctABxKtTNfb4O/uYm/RDP15qYpWd/T3r6U
t1qLNuFwlPb287skGGiwSqYhrXn2Sxj7ou1r/O7hplLbPXUw6Pk/44AfpFPu44Dy
qdajUji219GVczDgcgNhtMFVum0lFVwIov/kArCLKr8WWrmWY9OxlBWQQOrrfZor
35ak1wxbGj6DgJN1t5tgPkl4q8tsPMK0DnQATMYQOeROEmXNGI0BANGAJ2qqXbjm
L+MwJc4F1paXfN8U6PRfy6JTL2gnUi2e6/xVUY9MC44Cy46mVrp9rYS4KtFgdM36
EXw2nna5SMGiALp08DrQQkCkibvktHivYE6szKH88hJYdcO61rhz6oOgXlPgOJZb
i3wWZ0DC5Ezq8J3uwn+gjZ+9sFssEdgla4rCu3P4ngzfQKCwkCdDXuobz1YkZuNf
EG6KypyJWnc2nr0Qfx9rqbyc0Czq5GOo95rOqUWcNKo04lI2qYIGO/RdTwDkTbKy
B48RNzA79EH3ZVnlysidP/l5B7nWK4GpCb3XJuFMga9X8TVXLgt8uctBwMeoRSt2
6WaARDMkuUP6WQlfMZnPjickMK9WRQ1vB6pinp6JWo4IfXNj9NEAJYSiLGWLsI0Y
vnDEwtuf5MteDLidw/8S+QUo/+X8BW4gXTLBJJO+h2p2s1FPq2cJl/8+oN+IL7sL
wBQO5SdsNTG1E56yUlyos4C9DqaoWrX2uG+LiLLH733ud8KsQJwsNrc3L6EUcsjo
MqnKqhDbmiUH0otgwenrySzrjBClU3BjntztnXNclIYSgiJSnXB6ohZlgkaLEz9x
vqdskg0OYSrFsrJ/H30tDLNozW4FBUXEt1zJY+tPSnJOVn7BI/yCWF2p1KwRr33h
OqVFwZkTGE3l9RuBgQAu08O8+bBvb6ESrwVcwE2f0fbLCE7RE8iVeDIrhoTSoWHu
s9pNrCmNOxgv5r1odEEaLHwtX84IV/HganzhvykKUuO0/FfRnRw1tyjp5MBhZad+
3TlIIMGCXYg/YSybx+3jpTEq+O0+rojZMMx7hUHDJboANAcBq2KgKU8ov9ZhWWIA
oj3G4RVR0XdTO3bpCSkZWAPT3b6aOmzmC4RLOWyu1ZwGbZ+2a77QL6lRRyRgCN5i
QxMUWrzy0oz/5ae7/ycy7+5nVZvFxuwWPKJ7ChQR504+MwqwAQG7vo+jBidKy7NC
tdVl5smLLa/a8mE8EEvmnBHhf0qZNhKRsi+Bqp2l3lDh2SiKryNKS+yOfItw6zoO
+9RN7DXkIDllnOmCMv3fS7hSaUaIrLC5QQ827o9nTEfLb0qK/GUndIGgjamdTOLj
h5ptSxTzxHkTbUhVg2frE9P/qRHFJfD+RZeKc2ZM295mbpFdFrQ8Cy0IUsuUalDi
z7IywJV3Vr7Ynt3DkYCMDQ2B5B98JMd4TiRZUV2EvCPs6b5tCQ5KCCetsI/OWE4R
uka2WYfhFKoyx2hiNOZO4UmxgrHXLLqDqLcCqBlV+g1ZK6J11CTXPSXWDvjTSu1h
G25LpvzJnIjNsa2A9yCYXQe3iiR05Y8WAMl4YuVYO38nZG8dlmXyDy+oZjMo9/yI
Ay9CC23RQb5xuxsEp7qWGKvvjZ59A/+ETdWlkp7qPSUJ7ciCgdOw1NeTcV45gGNO
3Qw2xY7/3H89kIIX4TB1vJ/lTnyfTBqQ7zUz047hyV5DDyYUB5PLZTduKwbW9Ypi
M9pyh7i63mg7ob3vafKY3twdO+Co0RGcbgLAi83IupPMgxWKt/yVKLBYXCqHOt/+
pgXjo8151xvqsm0c1H7dNKri2fFAnkqLPUH7CQnp3yWxML2p6QxAuzon4LqZ13Av
FuZ3IjPbaovEmjPBjon3Sx/KQVNZCd6x8I7pIW8Rsn+qpxAtnqGwVdgG+ZmcrATg
QxpFDcH2ZotX9MsTUQN+ywy3gkNjW/sPfVhqZTxDIxGt0jrRMbl1SGv+EbvxTy/x
0T6V/DSguJ21+njgDZ3zb/mk9+t5+luKOzrzQwt/LPNPYma5LLdkIE10Dtap7lXN
P75MEM8D6v6sH+B7+uryM5EVmtCm/+xN4x8vzsMfwKBiY+zHZFp/tJ3B9Ap27Ozu
UXy+ZYPfL6Vmv7ZSimZYKQPmJkrstEVuLmmYQgOXWKsdd6RpT2/1PGdChrrGQh3B
qqk3f33D+SUTfXjkxBajehFYHRy7E5HIlWnGbB49Q09SExstraapHJZY6ECreR/7
BfqYjKmwqgSTYOyqIkMiz/Ipus2uuOrMzco/mx8MrhsOWy8XlJiCRfYxCP7Ru3za
S22wxy16aGxmP5F58D/3UOnN3IHjQY++Hur0z0Zk8x9XofXcaM/M9vfS7hZC8qJJ
1Chq65BuNS4gUfYFfUkvxwsxWzd+KlvIiMhM594RcDK+NBoAJv5XAcTDXRoU6WvR
yBVrVZaldTd/d7N80BZw+MUCx36c01ZSJ+Xfw9IpGAfkW5vD6MpeW/lhM+53EJTM
M6kxOdjKfYf6gfNUWlTcMbDTLgJYuKN09BMOTWgIRLIwymalxP5YONE9CpvpWrZO
UDeoVFYxoZ6bI3CpMs/fIyIai9HPHZ/o0mgeaEjXlcJKmz8exD5h514sST3ZpK4z
X9UqiRocGAz1qSqASNOYHwEfHyUD8okyoXVPjigu945EcBf+Kv+dqKz5Ba5Tyiey
ypg8oOyGM1d2bWRxUEoSTLXoKkBRlWDEpQW1Joa80xkyV8sq24F2VwqXeZ02PAti
Hr0qeITlxUC1GTxIlfQMAscYYWRbZzMj0iDOZKh10AWjDMpy2kSOFiE1P2H4QH4+
SYofzLZTOmQjplkInZMilZQlnVS3Rm8CGBgXFD+T9KVxa5PZO/VA8tI0rlfrADoE
+nKUK4f1mtvgV92w2QsnmsJQ9Mk2IefHndplIF+fOIJC/abNOAwSilNX/YRUUqxO
54Litw4WEhMXi9iG9OdpVsK3fjYNxrr2qoe4PDCFniVf3obp8qmnlGwQbOqe/liu
U2nJizkqpm0BCOzcftX3UPgWlpTPlGftTQHbWwDG1DeU0Wuc3sW873rY+m7WcGmN
tvSfr2veufpiA7LX9XBeQnsOPKw14I/OIzgV6Yv+bwKEpIZvu10deRdaMGIY8YID
lGBGFBoibQ86tA+0sLT0JkF03OlR6HHL97lVPkh/CI7ZOrUwnn5irSmqdGeQJPLK
4v8X3B2XhislFtem5hYqJI5xW9ZHoMJ7qIqlFjOErJnAssxkf/n1U5JQ6QR/pLFS
Hp9qgU9sc1SqZ3DbopZKIXaGr8AfrhfjnKeOufWQosyzgsaF765t1DPJzXPoj38J
jPN4JnvyOas70NNowzXKFhEP3S5b+PeXj1VPigpm+B3eUiEuYIpF7LynhElKe/z/
K9NkfsAmahImbZofOPLAOKJb0YLUe16ktw+9/fnxNjyu5tbxbHMd6SsL2kFT3eqk
Js3kRj5qUATWUOhHcr7Yd2lfTsGwJjOfxHlICZKTNpw5CLVPduH4ECFhmt71O5V2
upaj+0evwWwIJe3zPHlRBlJYFc+T5ozq4NEi71O8b9XND39SSxUs6bh2HRYmggpb
u6oVTYJW4xCJQ0Qg8VoYpDMaiDcpGn9ccyaSEd4E/REd7VSQM9Z2+8E+4341oYL2
Q3W2w8Hviywch/dcZCTjivVt6aMacBqjTAkzi84Np4HG8dNQ3L9ioM2BlHQEhjFv
3yOHLm7NUtBSaF45ShmcnJNZCTJgh4JxciFvhLX63avOvYvgLylRXlUmOlJumHN5
wNIvpk6dqF0Zg2X8iO1uADPcJOYWle/nno5xdNd/U9hShWY8+RFB9aRopqOGodty
pPCuE5kGjAu6bvk5NeVH+NrEu3YeVt20374l7x1MKYj6ewCW3tlUXBI+foAETHrz
G3hQfdIcIPe3BwHia5DI1LQ7cGWGlBxjB8CDjWU86ky67uH409urA5baIZgi6eGL
rt7ZyLIdajMBWR/NuSk6SGNB0htDE/EHnzoQr0SYgzSZb1egxiRmB+wT7Hhu4gyW
zwyiS7GNkOeRluxuD9zBUCFryognTW2SfBLoWMoURez5gEE4kxkanQU02IItMCNq
XslI7ybfMqFLel5y+eTys6+iqiSn8N1TErVSP09D0EZNcOTtDX55DTUeX8wnwgA5
oc7b4bsnAqa6+9m+kOtZcs8tes1n/6uSZ3gFg6P1/RwlA15DhvZEe+MgKgoEDHag
ow7qFQLoArpVSHHjL265NNod19I1nk+7lIYviTkpwFdDfWmENvZfJwu25JR1WrYi
DKWGcwIE9QOiBEU7s3ZoRF0uqU8ZFiHN7TGFrS0fe2V+gwmT3dPJ/aldhU5ahwEm
VxxUxN0QrpxBIk1jbC6H51qU86rrHNqCKGLGdMWGUHitgq4lSCUfMaU3JXu4vFwq
HS8C+jSKofQvP9uyy3e3Cq5DGMtscEolD9zOkt8F/QfbiEV3+FO4VXq64MKwkmhw
bAz2R5izTs6BSc1UsT0BAAKZ+NrBs0XRxfiFCU/HNWV5hkFwwMgPw6qBP041qjnY
gI1hQoRA8rBbllIAucown0jISTCZnwhc0wFWqIh6sGxtDVs6moW+4GNJ3TtSGn/b
aA1owG8PQ2XZlZrgdq3fMijSlrzLKWqbExX2V/av3or/BHhyHYE36esP5MTyth8d
Lj3oEujthVz9NGaB8Go/ZHeKgXCnhPtpS/texEtIZYw/XvW151Kqi+KcAb28l11g
fgjblcFZKFVXxDQF2Xr7uYVVAjwdNvwjv7PTImBYNj1VH4LPYqYi0mgUV0dpFQP6
vCdI8dNHuDpVzsssgUsQn4o6yQq49IpweiUn2DSXOreuQVI7CutwAc0oEdiY4Vmz
+A9MmFHaBFYbvaf+0Afps+DouM9IG8LYsMygt9hKj3OkSNw1ttybpQkUS4h7TEPC
Sx8aiGVd9vIgoQ9zGH151GB8IKnfUS9+z7bzosCwwfUM2h1u8SjobG5rJUOC1XNr
p3mlQK5SG2eLTOG0uYinbC/YHPTHQCvuq1iCCfXdhuboTDBsRzb3hRssnuVR2ceU
zTK10vlEi9Djwcg/vv4thHai+Q0xUHRr0EMyy+CUv+ofvo5WqGml3D/0V15/Z5OV
VkAGpwnjdLKu3SO3XtrcbUpu16XqbrajSYD8sQF7WpHN5Z8y8DJVCnfHYeQxDsZ4
QHoRP9dEE/V0iG0Q8wm31JWR7F2fzIvAVOfqbWtc3Y6OwbEIbynEjzhpcoNxwyAe
hjCpLLigQ7g5WklqsEWgCaAeYi+Dgoti0eHSlqozUAwbFHabmTNz6i5bjXbIJc5r
HvyWVbUnx9QMu+hKhr7be1WzK8sN6NgKJ83Y0bIGC55RDfyr6MFAdo6G2qWQLx6x
X5uIv4BuuaWkxBkZFa6bv8tnWB8PsUYc+fBjdcL+D5+OxlFJwMSSaLS9lj4gOyvW
tpUdJ7FYfPw5duyIY1FcRUwfC4mcIstg968yOMPSY6duH8sy95lOB6rTB64dLowy
Ujcu0lRWTpvzBOt0/epAj4QCMaEMiJEi81HcTbcz5Ehm08xEXFWbfZpWr3B7tAtl
twOaIv2T7GW5i73qivnpefiW96yHeN7g6gZOlwFT0qiHeNOaNV3d8RYBkRPMZh2y
cxgat5P7MPayDigBsvfk700ANPWp7UIL9M1U8ijc+UYRK6RVaPA+Aut4CI2BW+yZ
aeAzyiQA609ycjMi7BJA9JTgKdUYIV77tZtWQAR+Yp3cKFcidbT7Iv04DRFiuCIB
PyV+RFll10MkGgPFXXsSBsk4AxhIdjJnM1RryQIrkhuwfrWO6EpXjRzCIw+/ynJF
VvSdECBsyo7R5g4hAvEkukTFSg8Qn+iWoiI01X38GVdmDu2rrnJQmUkmuctUM530
I+RM/FvfHasKmI2+IGZ/UqLalb8vU7ekX42F0ViHYWf5QcNfDzQcOPuDNembhcW3
NpYYjBi6AElZQ+ay2bsd2j+rBL/09BbSwISKk6TkInoNTfE4elFSi5wb3i3pS0WF
7UdnZrzYsKTeQ+o0fpXckZdvY5yOHjcu/uWYlrhul333zPztgsCzBY798DRWzLSG
gfDOXFPIlGzFbXheILYhMOAO89hcbn4ebObJd6+9RpP/0ouzzxyzMqIQIQd/dDxV
RyNaMSSv1/g9SMq6eyIrWUR8STpMRTdCGWlSjxZeeOfdtKpVKGsXrFWqtNsWl6zA
F7GMfpxVaee3qaEe7YioQf0Tyea1KuHap9FheT252uGFdnqe+y0+OJZe5L4yRcN7
dVOlfMuU7hTJxY/tnlvQQEPRtC4p1jGzcC4CLroAv+eTtrpz6P0y5jclDYK5k1PH
lO2B92kPxnxPsbR7T+75N4TwiGKNSAQcp0tOqjk/H6cFVAlmhyAraan/wgz1diVr
xqwaCE+u/P0F++KMxab36WZ/h8aJH3DmQH7uDSLpaCKKSt5yI/uDk1z368X9WPKL
vXplhbBXizOFbrCtI4oM4nfdU8Q6e/PF1ntkrPOOIHaTb/PDt8P8mGf1A/v/uonO
WBYTib90oOcMKXPW+9LkOfBSa3Ab6k25uWbw82ebEW5DTRyyumDymvCT0hl3kOny
hsSpSgoEa+pRCb8RkY5ypxolfu/9v/cgBL1lOWi/xLUTs2JMo8dtiwSAryW2JWmr
4z6FExOFgCzpWFOkka6osa+LLNA1qMmSI3erg2YziwYeb82OffmYocAy5lU8LWmr
9A52CcHETjfKRekDq4tWO9eo5DW1GzGBZvbUsZJhQ1v67B5fKBATFjw7I1lpuN2q
bYgCPtEhRA/iY377IaIYVoNnKtiYLPl5bJdm9bMtqJzuEd/X4UCxed/Ri+tmSzK7
rCruHhX66MuE94kayK8OLzmQglYbm84uaURBn32llFNWHDPR6Pwb0B5Vqvg+Zwi7
7fXGj6NkkM+b9g3qaTx0f9sx3p8q1Cuf/0LU5qHfYzPhz64SVYEBe9/GzXfJPoZA
3EjxAzyYhKORtWjb+087qMLtwC5XWcU3piP3NnmgGNcpGNP0/pk0B06kAGVS2PTi
gASz9I3Y6yuF49xgdel73TssGApTSICzyNV6Osq31z6lyDPOd7O1S8XM+m81HPF/
c4M3Ht68R04sRW0qC9mecOBAkqEOVVkNc0pjPS7eU3RwYuhPzCLwS9HSz0vnyH9A
HR89HrYtF/TIJZMVZHe5sm5ARf1jihqut1vU89RVoggp6SjEoHL1lFHAM8GMRPcq
is+c3/ZXLAJX0BOLXzcq3t+1luuqXELinqlopDDiigfSDU/jQ2uzmuiQE9wesozN
YOsiXZeJERX/w2IOa/meUA0eSCisqHZyHB6ER+/3K1QHhBEYKIICDtxL5QUDhNpu
RxuIlWktYzIwjJTTqHM4xpC95MRPQiZZ5AC0TvtlCNHx3xSShM2XXCuOX8QLC+Bv
6OU4O/hhEP9SwgIls8Y82AIqtSSTAlPmLseHm69kNSdBq5iHwVzLClO+xPuflHyr
9ARdJIeiHuDeqCfGSb+KnUe+Dp6XnhMuVw2YrD9mSOE3/jdB7SMqiJwEvN7OaCTT
jvExhfC5R1/uSHKRxYop+oJ2OV6pyteRLY4w9AnRC4IqCHdzGWttrU50pPDr0DOQ
4QpPlSIuje6e+WT940L5dqRfAuodnaIL0J2rQIxiqNKGVPzv116x2lMW4FV/g/8D
LbKgwfKhCKH49Xm8/+4j/Ks+xZQrq5DKkogTLW3NMX0QskktavLeya7jl1yV/spm
vdR7rbdxZJPh3gS/frIqaZvte6/VYZVyjXmXrxGcKUQj7jptXDKyCJhmmzJ4kzOd
47w0KT9IzUXVZtTskl2ulCTjVO7dvKOtWw3qyL89YMrHg0yd7dY52JC6U+sw6qXh
YSZfiu8e8dSFkf4LlREqb4QZii1RgZAK4hOhm1slgg4rj7Hpi7mpnIb6l8qUdvb8
05LZGsaW4dr+GdI3zaPZpiGC0hT8B7Mfcf4CBsV9Wky4ZNkPDCSbrRfrgfwr9ymc
Yr4I2BGepemqloxWGf+oTQi4dERshmmT5bjo/yax8Vhb8FzOOLyeLR+NVqbCT+bb
Sl2KWSJf66iTfW44XR9VbFMWy22dumtp4KuVqrInHt5UAa1UnR3s8QGQtospbGbs
h+7FEQAi8DWMQ03lXUpYWr7+JaKvzOSHUjePLIMqoo9xaUPTq+sJnKWnF25K4yqm
/YYClSAiNZp8iknEiVreyMKV8oDWOAiS0maZnkAXhb1gz2dRadh+q81j6A/Vp2Rx
4zjw6GBNPVNi0awnHngFaL+DYjUBFrzD+KblRaqDyDOJNSPL6P20THeCfSkSTdkx
HK9rpu+eHhEdBdwx1cNhkuYdVC0ebrVZ8T0bbKdbiySUJV5DQwA4Ish6WZpQf2j1
3jabK/JnDzCcPyevIOwhtFZxFB+aVoga5Sm0o3O9QXOXSRWxV5+XgMNYrR0T18hW
XGHtupNkzMliq0z+xOu7bVrSvCj2s14uGqdZSP7NaQYvx0QInxX54FrEdSb4AUKQ
Dgn5OeWs+RVWghqWst2/9DHZUVhyogsjIwILIe9w3vUvsi8+dXqfP7NIHQun35dI
TI7FbW62qVUdR1AtRLB+5ro2/QxGbj8LSDyYPnxDlngKHbsd5tOy7hQiEp7toDJJ
3Yi1OyD/JTgC4g1t3aRQYY7kyr4/kaajLeyyzr3OH+Ni+Z771LEWw78p3gTsDJN6
/OC4gqeZpPpQERpaKflCvRcLI+rdLY5w6KoCjQAm86ucCo/L8aINI216+oxd6ArW
bXU3Eget067YqmaRiUD1mzp7VxwCLrMOvipWdeUpAf5vEGoZmD4ncIrPhwNpSkMh
y//j/42ZPNzvQa8ZehpFOneSNyBAlBTre4ajiFEVN7JMTrUW6Lq8b5NcRUm/6nVk
/zsnNqrEr2St4VlfNEN0dlO3H9jtLVevsPRcDh3lVhO/SZq92FUo6jCm+SJlctRC
uxUCWGTtrNXRaw7xYkgHxX9URV9GjGI6IQGjXxZzjSReX8Hu9bKjndpmdDUwIKG+
Iozu/XCdyaxj3BdeQUoHzdS8rkk/rmdXNYunFsFAu1l7yEiRqn9oFBfk+91wr3hM
p+RSk9t3pzIESSoYxGRjIPR/tp1j6ZlUxf9nmhrVaBgd0o4a/7J6UD+v3EbAcqO3
XSbTeFLFSDPjUgULo7lDRJelLp6Xac8SDaag7AK7oO76F6gg3a59zxhGtMuQWrdu
ZZJrn8MXpDitF+8TlzT7kQZYCJ4otM05vdSEvw1Rfvy4uo7BwZUS+y5Vpjl160c8
8vLtWJWc5kY1fIuxoKYxEzW9Ng0RfVL45yw++Bv73rAuQic86cpF0S3H6Is+h0pc
1Gaj/iLTOsRLh1LRsqJjAIWk4ej4JV+fTAtmzd9MxbqB7V0oct214NLxeTxgkV1Q
4pZxg6GADn+O17QrKZW+6JSDLW//+p1EV8PiubktIA0JWZX3i4E6ee0j9J8iR5IP
ZxcYKHeQXeM1WwFunZ/2ihHRBB70jeDu/qVk5CzoAXGBTSMk5kTD/B2wEpNQNi7E
+mcjBX17wh+oc7wkJ4z/oh12vT1Gg2+y5GrzVn40Ri2jwe6pl0jhh8e5yEP4DPPy
xF17fLQCUUL0UakcXZyrpAUwjhp6Qpk3vGgW7ahNaClE54OGDBlNtP3in8/Db9yq
j9ptzOgu7gcPCLj37htzmKHLnK8AfAeJLJGiwzclSWWKAGrWf/8o7ix7mB1VcPxI
Eh1VO4m0VlS6h7ImkevbJbBmgMkIUIlu/164OPAfrI5iO1HPPfOEjnfW9cySqwIA
2m6z6An8ZdlS85wrt4fh/+d3SnRUMfEC9VOfQI8H9wETr7mc7mG5LMpiLk4YK1+f
84XvpK7LwV10OAwyG404ujHwBPm2+NmczbjIjb/01NauhGrlMel2wumXWidxfgg/
T2jqwhSIXTefHtO0td+GqqoqnhM6KYrmKIAeZwpC0CPLwFIbj5/S0T35D23u3zim
GawAgN4COtdhJir4GA8U4iQSh3MMuZQQKpuiHl2EE1BBQXvRitVSDFmDgfJh4hyy
9fSUBLdRe8mED0+iuvmPVk6vDJHIMRVaV8zIX/9sfMxHE6mz8ELY53ScNmHpBHBC
uMKtLAp3tdYFbzE3uTtkRUtO3yDei+pbf1Ry3BbhnKXexGjOGJVCKejLUUAdqPJ8
pp/ngdiH0gF8wgx+E9K7oIWYuWTPHWFJ3gyxpUUVe3cuQy22FZNDMEkYMbAN6qh1
ckgIEfUA7pjKsle3LNmbjqC5FIM0/H9EQYWMhmnsDgDo0kmw1fgiSWqSUi5jUaqL
79Oh5qmGQtQGjkwO42JFK5xM7k0JC4YIa/98xOCYY5kRUUkyJ9djkDcBlKidIVU8
0T4gP0j7OpPzv8jj784rNwJ1+XWn3aB+1Fow9CPTsBYhV3x2H6EURsPWdlRHCJCH
IlUcBMmijd/7EeJbiOPwNEiP9JCguutJsjV9o5PYNymjqPl3mb53PQ5BRU7uC4wm
GaMcP5GNIO+ATHQi1OzgtOVDKD2CnwaRIftF6M0eQ43KHe+15QXMeyHUqt8XxigZ
AeD/OwnWuhLImf/bXq1iU8zgYOW2/6qusD1sDpTuzn9xgwEgHssAXMr1220ay6jE
Xv9XpC1Lh2oKStFmAYeCt21MHjDIKakwCSaZ5HVeiQDnxZA2JNLULQ8rRBwqIHtB
GDIKv/FBgBgYAXvc3l3ybXjhw76jXOSoFC80lMhFhDGRqEzHB7Xebx4CK0NsoI9r
agMaY8t998B7mZJqbcobzr/uztqARF7NA2rrMRLnh+2Y94k1nnP8FOIZeydTm+po
X6I0Cj2xZHoymnIBqRVWx6W54nPRHXCPglKjwd7KPv5swv3s2go9Er9BLLN5o9Ek
7AoO++DBtX0KMM79PxvCrJogHYd0GpG7Z0f+Royzwfn6MMRwZKfkmAE9wYIfpzj3
1U078gxrBG/Ce9XUZD1sW8tfN8E7tFTWpbxOTA6qJclfWQPv5MeyIWjMm9YfVDkY
6tRBvtei7c/FzwL8C2psLH4N46ztIWIpwn2sGQw7RivAYliFcwLYdJOMuLq1/A3s
I9b1g1Az+mA8Y1gdby+Y/spRn8iny/8s818CR9LB6rcIiLAQMZWKhA9tmXPUwqNj
9r1I1GlvKPgkG/iNDVJYaxFpPrBOW+yfkhx418l73TwbEtJhu8qNk33X5BsbTrS0
o1jn4WjxRECKoAyXBQo1iecKJbRlEteasHphlipArhGz3HnDrnmNfZ68/bSvY/ad
0nmM9upnTt2hxPYfQrHIAwpSqLm5ofbJnik7bHTQRAZLSwvyBf4GUU0UGKS/LLyE
CZW166IJe6kuyEL0AOrnmg1M9gS/JyTND06q50cSLjFD/iSSqKbd7qqOq/TmC24m
HwMJSDGOv349vTVNhNBET41zFxSPSMycRdFF+DXIdQpi60zBw2ltcQdsIXdZTo3N
M4uAm10G5X1AD3wKLTY18dFKEsfkYmb5pFoDs7OHx1ir0vjv4KNPjeEs2F7MXuYZ
UqtE2CRKB7/2YtaHCh4nexH+3k9k1bSRsI3gVQztUvL5bFNqTNQkhQlgslxeHCJw
9eZ1l8zKX+aLH5SoXsSNWsu3qhzZ29/5U5pTUsXexJ/wy2gC/f0kdB7yJAJPzf/C
CoFYFqXUZ82TP4GItesGQahXZaMrRY/PFSbJG+IGaha+mliUFVUgcb9lkpmGs2P2
DGqB8/NdA9fS7/VaX7sD7nC/uEYP4IUMFAP9j02fWZjFIXj89ubped7zT3001YqI
irSYop8j0MhkGK8Hi/5U2JRHf/k1G6+B1FYJGXetCCv1DXwp88ZhchhiCbK854mL
psjRuiG2xwQU04yLBYUiXLR3kYUOhnYLd5mX2Qh9v2Kw1GZtsgvscWp0Z2+V8IbC
kV7my7jU2ze9cnQDhJApKPMoCVO+7ms9tWriMNWbk0tpJp5kO+krJ668IsUQMvsW
ZBDFOr4i0GTiCxtfYRkvwhJ2R67NjKG5kn1h50Xr4LhADBWb8oWpkX1SCWT3ef7J
1bFR61cw2xOLmCEB9HClgolB4g/BajDTIyKPrHDCTlJduZ4rmtx4RUuPtbC3htVh
IBeoIJrk5GdpLzvBZxlIHSsZvtuc8lhjKRecllPUwqmDlcCMTEVZcK58IO4fmrKp
o0fqHp7zAoV+bYCcZP31BfcT+eJ19Jr5+XuWntNwQR7d9xSjh+XyfOvTrQL2LhJw
ltjbRo+cRxxTCQq9HZdGFwEVLrt+mV4m9vNIK4YWjah2CMP6TzJKJzGe80ysX+zb
rHxSAI9iXEWTBln8FKz974+oMryj2yINeqrA2tr/mWcsP1eSmlLCVRMxCHqx+HiL
6BYLZVeA4xOWopmmj5NvwYpZWzArdUihqJv6U5gyNonmHZ+hU04tyMfmfh6sgnWz
t/QSEg6TEi24FpeeXZviF1MVS01Y2AQOT4qB7SFZWHDw/S4Nf6mHMsPiY1aKgeZs
vHA9jebTaTJnchqeo5QYHYNzJSQ2K911J7ha2g67pZZahZTkXQgOcFVWUZXVBQXd
93XQzEEnRo+cMnGtibWka3IRZVnGhxSl6o3EfgQiEN2eqJUgAVzFAcAtEJllGVPS
LqNxf3LOYbtwrpFO40o5ZfHvf+MggvrDFW5Ebu6kjkJcp+qnuPgQyun+m0SzhU9v
9TGDNlMTZkGTAMBEeJYWJbFrAv0wyKxA8AQUm9K9g/DOYAWqFp7ytHxQMzgONM8N
HweNZeWYT2ftMXeCfBDIoGrXIPTovAFnE7EjiN+tXN0AUSEVrYJ2cF4I2XqySmb8
N6oDkVMCk2rFfFbeEIiSIJTxYE5hsU6AsmXv+L2h5hHutUUFOz2hxW5NH5t/jmI1
1zqTdkznHi5eKkp7NW++Prp5WWado6rnnvO1cCol6vBiyzAln5hcIrimPAzNziPJ
E207UKGClRCO+C/mvJArDeD201IdzM82kg6E3zxn3wvsbprh+WtnKqxy9g2lEfKQ
PNOvVEgF7GIx5rr9RenykHeIAxcwd5fNO8aZv9k3xbFUHE43IvqJUf9PuMkYu921
ETTjL9E46n0uUuQOzyKDVTQv+GvmSydctJv9RcWVEIc9x+HeVJrHgeae1YCT6QxR
1jNYITRXRl1VF+HmVzKOoqkMW5FwhXPH0AnTAlRoIAWD2JUPmU/YdslwP4a8KUp2
08whtjdMizDxzQrvvD+Dm9efPW6oxsq50JFJBWlR5UUwJ0VizUwvu68gzWPVoQVf
1bClxmAcJ4DHCLMIP5RmDWGE1QRwYx2FSJj1UjZc3yqODESuRKcJVfeLLpPwb02u
P6pztH7P4p5JyFxppEPD9qodxKjMKyOsOGqCY76nj6+G8jkHPR4FldoTef3SGKde
oMbwJTuFQCoYE5mZxC16dxZhFsa1+diLVIhqx8O55NoZ7/xuiJvgJF1z7nApryGB
QU61SS6L/laRp5PSmLm7/pcuCSbbJNDXTeE7trFGeXwQV8gR3qPS75NRqx9Xaz4s
NaJhm6Au1P5VJDiQbPNySZhLymHsvIfJNO0z7YWa3CzYyqvKcTuLxMFxm7rxqaod
v+56rey8aGb0pJQlpWTgYPUO0UCxYQb/xw/YuvJO1lU/KhPJeyRl+b8nuRy2OY0f
a+nF85MiAgU5xJTNpL+LSFsO0h3ADoBGLGZeoapWZ2U12O0vjP4h0+QAZqgO7tkR
aj/groYQez7he1hKXU6VOrtJHjrkymjU2fJTrHA4AYoTDS2Lky8/7sbHzPHVDq4e
7xEQ3XcVRS7y9fzwL486Vvf3yF3HIkSZucr1m5m/T0izKpPVztrMcPbxPtN7icKt
ZvEF3ILcnSwCPFN7p/OoLX8gj0QIrEtJznh7jMA7+Fcx2RBmj+OE7IBUKizvxyha
HZg7yBW4PIJK9c3yIUbbymnlQDKc8heK7kOHRbIeZRPWjlQTt9D6igONu2HS97VM
O2r/QpzfRQHXyOjoDcS4ylM2sCzqCU2oV+N4w0/Heklh/FWsyVI2qvifjVvkxCY4
YiYGvXskMmi4H8mn0K4uXGLAp7T5hn29jMtG5nqreUZB7U2oGVc7FljjSWRLy6Vv
Y9VqiWeQ4ZJUWnz5sM7que1znwojaeMwA9IuapPBUYVADRGa3fOEVuhUvxIpVdKw
vsyU52RjHUMKz9nGLYzb1ay5VWRkQsUMjThtlpJ6hGJc5zCOYm/+dUunJdlX0Xxk
ZQUapXVY+sbOr2kGiMeH6TGcdU8zaRGs0IM7DzkcXl0NYJ6fjCfVbcCCsztq6Tg+
6RcAJJoIyLF1poWFMAK9BMpRQSBkwPmKnt/nBcRzmzp/77c3wwomV9Ur/WqXHxXY
EqC4aSvNx1P740PUXJDtSgjLtoorsYZhXf3tqQzAuRvg/Jq/dJohzmZUPgm+SmsA
AhdOgwzBnT1svPWZ1RrlH2mmy02PQX4CHDwb4yjbqrnuO6OyHo91EtdCLBYtmtg8
qPIuscd4HUD63gCYXgnapzmVu6h3zE6R3/WQz3YpHTOv0V4gSsG3bl9b9HBPTQcQ
oylnMivMSRhlxeCqn+yIVLrOw084IWTfem/mal9IorSMZ3eoKMATPdGv6gIT1OQG
MxuXaTtpk5NS8oTKkZ/fSxQ1xszO7RJ4ZoTDGCm55NTQIBHR0wP91E3tUa2j32X5
XtGbrrVHFxUaClbj651A62L88rr/dAN7X62cOFp/yGbeSBQUY7SD/Ukd1L+HJPGt
jCN0iO802ey5MQR5g16RzK7WgYVmnhJRcc2jpP48e7iqmezrXUswDtKFHf5li1aE
lA9eM5Ja+o1YIGqDvDgkRhCj8FvUYmMYPmZ2D3smI4P/wfdeySEvSIwcDycCD4Wt
chPuzkiDE/HqFkcaEClE5BVHcWEPJ8+epgNP8Xnu3+2ausZer6KPKsT8iz5pERHF
BwjTtelwbEb+aSE9hy7ONDCI2jxXiJVh8yyUOXUsVbbOLrQeEG01CINL3fjrt9kV
r8AALm6ZW3sa4NorE6WaeYljlUb5r9n8CU54UxwagUaVp4pW3tQqR2uNZSEsl9i0
8bsmfMhlk9TlMXFKWpmVEcvbuOk3TjWcygqceT1UyeUQBc47JxnewcMLFC42eVZe
Nzfm51iXOWYJKc/XIPdagA/AKFGgw7hmWaxrT1SvSIMn7AvaNooUypp3QNSDSC02
rUwZh8bZdSbit5YFTqwKs7P+hnIXYjJXw/hoVnLZuLccGmlgzh1IZRKL2gjQRSBm
pQsYP4K24ubIwNOYP1aaOZibdmkGmmvLlEpQvekYmks7hl5Pjm3VDaBZexAE3wiO
82wNaPczyF76m0aWuuqm9M/8bCRNhfUZpvcKWr3IzjwCzm9ABArNTmU3QOaueIaE
mkbFIZkgTg8kl7FLvi4wd8Tn6BfNU9BF5WLQQ9IlPrAZ9prCh8caOWMemBYhDUfv
8dPSSkWVopDFxgJvorWhCMLUVZlwzfIKrx6TepldPtQKNcXW1+fQqudBag8cl/8i
IJlmjptvvwidzizZ2V+0TJAllh9APanHbrMaiqkcuFlorkxwWTrzg8nNtytdhChD
rIeI1+qKHdQH3jXt3RGnFEa1sSW0lDn3GcR7kZI3dSBpEmt6irfll+n0v99j1PGW
cPBjbkLqsh+tKGbRYtIgRJFifvrEyh1wUCw6h5B4KYu3E2LVJl7DwPR6Pp0SoaB8
vaNbOAkE6JxYSotDxlICsqqTvHAMN4d/qyJ1RodzQGODKQNle59PrFxpIm0JOHnR
IKCYW9xG7mH/ND1FshLK6feoyw4bdxR8+yvY3pl+0d/t3NVqXg6ZKCUGzWLbbYje
zezwPnR0o7q5G97slz0bbxMJq1Yq8ZgNAJA3jSi3wRcwYN5mz4uVFEvB3VQQ175w
9X/CZQNglpgSr8OpTDXEL4qqwg5wlJZC2bKWtCHJljRxXN704CUwmcNdbFYPe18E
2DOQ4HmaUOAEMjK/JDSQRH4VIl/ihAp9sWyxfD3xn0UlP0yAutF1qJQl2Lj5LNRV
PJyHbfhxk/RCrv5GBoHdPeKgEePFQj1WiNKjW3N+fDh7zY4gan2QPP1Ultb8Zq1M
D6ev9pimwOf6xl6VzPcxTMi/FYSqwby4YIVSBKu+qYlGKVOai0VvbJtsJNXJctGV
hu8AOuF89JY6BEVmguxDQDfI61EhiNk00ZSuD/11oJqbCyI3iPGsINNbSsj2hobx
VSdUPB0b0+13ah4tzeRxoyNXUaruaqZacimWCL+m03tMqw6YdHfrSyhqlXiGNT8S
LwXworxow3sazupJw+kSCu0Gal/z3ov4s2lcAkCC8xhA4Tz4X1Mv8EQH9m79vvdp
8RuP2ezpFhw26c/15S3EfMYmUI+qwiTJuwm488vRS/NabKIGsNtIoV0CWzdJDOQA
1FFDJoCau+xaDM5VEE3UZxG++Uqe51UQisqVy6JUtivVZxM3kGzvZGMGTK6Oj4EE
cnP3uE6knaNdeCwHZFtMz7TQo2D3wyJVu2aJm3pm05a9JNgduAUIj5BAKgCxqicd
ubwRxR4bg1VrRatAXy6T+CcSHFdCy3uPQdH49+/zRAL9ZAxgMERbmu4d/pnb32UK
kexZ9M8AttxP9iDkDKEbJXyknvPYcP++lyfibL+7TeggyZmbK4uPJOHczVFMuuCr
sjNyth7VyoQKIwcEyNBi4gGLnZmWvjDX1lxAeTh/kh1+RksxJRniKvKcoBBc3Vqp
cwGCcXZR6lBQ2Xk5DUECFB+OoQJNE+jJ4hBVoROq0Nq5NJhMY+g1CRjMjCTJ8unX
cVX61THcanCKRORkZ/OXomNqzuBSsNWFA6lW2ayxxCbpALA05/S+de88Dp35CWet
DVZLCCY4QH4fqmWgR5qDIrs3vlOc17uO389bVjCgNDpqmp+bLpSK5KDdPTWIziuX
fR+IHvxWAaLrUZe0k97k5747UgPbC4s0kWbn6pA+v5wvtFWsX6RdAtofW6cILPnv
Dj3DS9SlWcz1wn1erOmfSunh/XYDyO3ebpGOm+oBYhkppANITv5nnHTfHrb5eZz3
0WE1V7gjJiAnS7ym0q/o8JE8sXIeb4aHMyqVpBnbqv1XN8UfW0/nyuOhw+7uBCzc
lwbB7BJW3JuPK09SbQCoqyUPFqpVA681UhMYp1IA6u5OZ1wFu0L8KjtMnEBQxt2Y
+kxqqIwCVsywX8u1Duh8FHUEaM9BqNVG49JijH4vop7Mh6pISpW9zAbL3M10DWFN
ieuPTVsr6I9jqv4x1FxsmL8a+wfybndcP0z1f8mGRc4b8qwRLLjkiXKwveK67dyc
KTa6Lrj2qDpmfMVOhp331OOWmL243+gPGc/g6UmXzb5DoCh5S73nyIU/onQuSjPd
yJoYk1/wMcpzG7lculO3vZezoP+OeoOn+3l6Xa795oH7CRcPZxFP4gOt5miYNbA+
fcCGOWcLVXdZXHeLenXcjraZj6IDC8MvYLlPNWEsBgBPdF/NalVci/MODg4D2ule
rjhQxbpdqdtZ7OCm0zo7pDcIYpUqSeJXiBCAQ0deMMKwhABIrydepJl+wYyDmM5q
E+4mDlLXngo8IDqg8g4aRPj4Z/EEOzOwMguOCD2KQhMVivNNjxB2Vi4NnpNoujzq
UrA+QzBnk8gjXumkVxE/LOIhzBrZtdpWxm+KAXjnpXNYAFOvDE/f1HAXxwTd7D6e
42Px0alVv/UQtdDDXOlN3KyYsg1vrYxZc8H4oGuwup2GmsE8VER/14s0S/svns/N
wi+eyaCzBhSWXPyITlGZDlBurJQCJjqlPzFAsnNauxWtuB15+Gu2fFPb3Td4KIyX
uQNL2pzjyd1kEYmlJ9U3dphkhcCa3JoZEEXXGVUi499X2On9fikQbR6L+OZWBGUL
41gqBZWusyr3PxM9hoi0+leX0RLqTIPVZ38WmToPnPB6zu11hrHv+wO7mfSdc0bD
/5xyjl1+XYU2Q1Hb9WO+j7zWM9a1nnkLNjdY5E4l9A/Ig0IUSu+j7YUrXr9PTrxg
0NRbGEzBhdEBcW/QbODm1y3IUPC4CvZwrxKyAeIpPPjUzimt+m5oIxThJSHWPeAZ
45myXGxLM1qBCP80Kp51hqcQp/3RxVZ/LASYY1863xswnuJqTeCDjnMj2lm3IjPF
4m2NW3ztthnJwE7BZrzCWvhO95bnbQmB1+byv6+BLxL6Hb5nqcb8apPLHS9uKpEs
W96k0i+clIZNktMdu2c/EwfyiNf1UyA0L4OjpNxUAGsnKvR23DeouUZZ343DBCuS
TueRpaEezxPEfG6Cjlxve/0qGv+3Pd0+gEgxTpyjwJ6B1Zf22wptbNRaT/C4Iiro
NOBIDhOO3nsKSm40yIenHBeah7CmCJBWjbGFlbgfQND61mdFMTS5rZlGeJCP6Yuo
Sm9hnkSB/wdKGEoxIBXaLnc5ZEmYKCuRdiiKmHx9XjFFDvwmldPl6bR4ySND+PxZ
FH56YxLtKK8T50Di2AXgj8yTNw/RhX2zRkUQbgCJ2oaUuXHtYUSDk9Aha6CqZprH
0US5W+4EKQgGEOylMYr3BVm/yBlAMtyvRjyaZeP30AlOH32l7WSQ7Aj/U+v6DYmn
hxByWMR+NXQKjbaallhIY3RVBHLDGMnFdj//a9m6ldTWP2nk0IzGJ7p0vT5giPtT
zVBxx+vKdvcGcb66IbpTf5+myN+s89+TNIkugOTMP9RzGllBeYtNP27+ozst7dGh
GLnZf3is0tC4+IuCRKkHpWMw5P3CIfRrOiNfhuOD1L3us0OMGjO2niY9aMJpOWWj
CPvw2Q2DlhBQreHHqcYeVIg7iYiElMQ9flzfkUjWNuPat/DqbXk1OsT5Fc6/Fejk
k9m20JrkxWp3X6ddATJYyTQ2GQ9oVn3Gb+25HLbnd+QnT0gU8GKSjW997zs+iRfE
0ktnWMX8yjLMEmB0PERkQGknIiqVtuJruKsuePO8zZZlVuSJKrDwy31ap/Q3F/qq
ZEa/XaMdHp7DdjWN1DMJiQ/nN6PHFDdWsjBoydf1W3MQeasGYmttxP5nqwr9KwTp
tCqsozalJGEaWBLwDqEgX6CVDsJIdVuJSwzdpkxtVyqQm1Q65R3hWB32Ox32Kc1C
OdpDQcF1hf6OP98wODB1grhWQLbLgrvcc8fubF/W0U3htt4nbm7MocJ2qQbQDRUQ
QgQ+khgzKWPhmbwce2jmkE/Ye7yZ6bBB9qJhjx+Zs+I1bxq3yIgkF4ekwVMrzqBa
x+N4MfU2FWvCoQFuGjc7iBa2gHP28E4jaqtaIAfIAHB4TFguaMIaA1RCdB1qH+S1
DXngJNurS5Rk4JVyKqRkZS6jJ+ZLmrEu5covlU/5KkycfJ9mlgUqfBSSoZZHDmEB
7jExQNj+SIEFID+dHwJvdJLloIOvMDG14G0cOaN9Mwmsg+xc9AHcL34UxcW0pqd4
f4Ke70jvt/BY+0CJybYf5GY7Z1yaJIj+1qn63ByM3Q3dUs/S9eFaj4xJf5NBzbZV
QLu3UvG9eKC+wGg+L7QruQgyih+a1gXegqZ+mANK2LDbT4j5uQL3ikvf7Tr7Lb7Y
o+bVVvzXnVOTz1cyQi+Z+rfWkEeXXH6apesjGjx0qL6Yw0FdDcZdUvXrM4OY/6xL
5zKVz+MY4tnM2b+4xPeMVwxiLZhA+T9ImyY64HAI2Pssn15geUxS8btHSU5U/Mdm
J/Lx7xX4WJJKdTHYj8FwDC8NtGaTBM6gCCrXnUA5DlOpkgP49tlKnPzUk1cX9CYQ
FybO1zh3zZ6Nv31+LTs+h5dx5gHOKbMEa8GOM4c6IYDkXSD2c7oOjsAg64pTzN09
RoIS5QDnVpVi34elYmXu0MYsEWJZ4So/Tu1Tx4FRrB5/5W6MDhkC/QY8ui2nLKwe
n5PRY9OLy/cLw8p6RfcLkT5RcCv05+mcy2RaNg1Q9Ic8lTSjoWjXFIRbeYJ7wrwn
BzU5km3p8BnfXoCmUhTYVjxpxrc8D9Eg//CfTS0lOOCju5IgTeHjhX0GaVKZaXB6
6kyyPM6pLUkrdK2CSIJUPqyJeUajWyGNr3qd2CQHb5zR3qoJVFwEUettzOarjklJ
tZ+5g8kpkUeEpRO4RkyXfi0E7Jt3z+b43F4VJC/o67XgBeFd7pk5Bo5VfPbyxfSE
vtjmFBqBDtlVkoBhdVUCWIo5QKl9jrijPFyuT5U0zk/e+W2vj4WlBYE2+EG+GFy2
f1C6ZUko9cOUtI5+Px9/nMigXOJdfCm3vyw6xpAHOJlVYYY9gwsF2puoDUFt/3en
MCHNhdz5YvqzpwJras24vFHhL2NsSbe4xM3k3blRlQPKu/qdcbfYBm38fKISTJEE
SC3OjhtImd5JJvRjly9RluLHddA5f+VV4s3jhNGcsGE7Sf2lI5O6jMI2Jf6g3Tue
wFmRkTrwvWQeSxtCExCN+NgAWB13u6xbuKOJw0MAJNtujg2tRVrV2CRFW4HWoAA7
XiyxcEPTgLi2opjir8jhRvqQBQa9ykvF1jYVex5D93cnyJZxMEkHxLMqetJnsWZV
HImPRaMQG+mDG3qfKxfUMjf+0xZrqhoeI87oBQ9v0hCO1jVttaaSvWMuxKLDSdIB
+LyfixemDWntk5XGA08hzFH4HKpavT2fv4zFAUmcYlHD6YaRpnURZns79+xIPVfP
DOLALsVY6J/8vRMfvG7REu0wrmRej3vd7lFAFeAcSFuTiRB6KukU2DL/IQphn18/
NDJTR3DT5YQ5mbxiZU158I8ITl4GgNdovkc2I3wvMDfxovSKNHZHlnW/ZcUSI3eN
t/qSFRarhmCQ3RUVnAENObTyie8hhFmflVlTg62zN+9yZt3O5MCENLvM6Ffqr2tf
bKPS17171PolMYueq7NKQ2OMs/VVLHCctgrl60V2jVXA8sq42ik+jvE7yJcFSL8z
jRpa9C7Admf7xYjIAo+2dDbnbIkJklYQm8wxI82Yp55EUrCUn1o45ZEz63ZzP0xo
3KCN+D5EYlhZhlogcnx3CYfw6si9nA592tn98Hx7GNglQpq7YizJXvBdN6wqYlmO
XWET3zCamI4bQDZ9enn9UnADJ9fZ8jojjhhL4zCgsy1KX7itVN+N8ri44ogZOSKG
XOFzthWqpZpQK7Z5eTleK3HTYsUHYu9OU3+S8bfxuElzTTgBpI75pXO5M9wroVQ+
57RCYAdqSn8AODp5Q7NMd4re9kUb+AmOqJDZ1+6/uQvyNBk4hlH41W/pGic4OniG
br9/ew8vA1XMXqD0DGjcz6PvGTI4FD1vgLLPVH9q73pvgBd3wh3t+PhuPxJFT7vJ
3yBnCK9ITKJotHN6LZu1U9YqO3RxURt7z2eVfw/yFjDxNzKza9HwhjoKhu3uCPUn
FYbvw2b2Lu6xGoTwD8WbM7ItcSi0M9GHapUljr3jWn5cLELrUVMGL3VoRzp+ZEe4
cfLyQeuRRS9SudHsbg4BpczA0Oa8Hnlb6XB3Z9Ii3vgbfoxLSh5V7/jPtLghjmGI
dH3lbF1fN3PcHHGJWotiZm6+LjMn/sxcOsEPwcezDGHjNQcog/YnQ6jZenQMPb13
2QMrT5bncFoO6EivE4pf0phsLgQQmwJFK+VpiK1LijTOXDqiEz5RQtfELXvSmf4K
C0PRKV1L2TvgqONC3X7UsUimEExvjDqlU9+seWwE2Ltq2oKdA1J5NX22MCzE7yoL
KOt6Hgs2fpT9UCxjopnu+YD19IXU2pKFse+xmbU67PV2sPgoPPCb8mBnWLI/eAoj
KXfndMroFnpNdx0nfwMGzNqbBOQuHEANzLw1N3nFWemG50S0cQax7khYEHksjZ06
tGRNtnpBxOMgu1azOqKf18+lFJ0uyFLpJ3rohLLinGbs6woD7bXS90XDdpT4Drd4
OVtjSD0cIclWRPxNcCuYYATOsJ7tJQZitaiCuBfsUsasKQKBlGLrP4UwA1I/omj8
Yr8IvMiA55hfv6Xvq7oEmNDIGhvNsBn5/BUSo/rGTHNrzaDfiDK1l7a0Ox7ukNtx
CqH14r+Z/imEW2mJjFfpINCQes2765yxamwhaKrpv3BbCT1mfza2N6uV8+5WXZeg
OaX0bfJtdOGpOeI2v1m/WLLtnD/EWCFYyzMzD/p4qivrq2WuR0TEO6gqvs1o2yGF
fyJAQWEBAY5eQneiRs264srL/4p4Ydt6pp3rP3BOpyQRFtnmftdsjb1X7SDx9ACC
BjO0USwtkrMyLV5PM9BaYsh5Hr04nD+//3xf43x/bTS14xyHZr3bnRf9pRl3eKyk
t5Gu1q3grGrPEFkSYr5Po8ZamPKv1OXGN3inzBOER9bjNYEky3P2OdUOC8KyRpRk
3NNm12lEuvhNY7ZuCDv88hhSjJxoCI+oIsi2/wkVHPWdeXby3xHt+IUT2b03xDxO
cmecQtMzImpmROhObiii+kECejU2gk0aw4tjFSiSEXp0YhghY8S7tvBfvSzzvWdo
4oBgjlhv0gdgwR6QEPDbrzqeTk0452wo6wCJDB0obNsjQ+suT3ixVsLcVsDOtMPn
L5tUZSqnlN0cS/R25AxLR72bgh2DWaVXTajTb0WkWS7LmM2RxpDx8zC1DX2e1sxy
Se2mv7UWNihUuz5MFVDVRUdGgB41qpUV1ay5wPyo0dMABiHEAfLPYzRGO2vga14B
dkBq3aRZ9vaqWXqfXOfUZGX4qmDZf2GOnK8MUWccziGslK7gDXSB2n+Twm2MLdDL
uXrAUbVLaJYQ9hB84T6j+sH6PKR8GaPmtewRkF8JLUxoP4elv4Y41mEhkLH4+AcD
vR/vCKq8y7GgDhVu92biWVfsW5d9gJSVXmChP3xxq8NHjXnGRdmowOkIhwGZXib4
erSRwglfY6RCkxCCDQzZdFIjJv+UC5Zhyss9qEIjrGCQoRtq7a5FNAfB70SCRBKw
aM0KDJhUkBEZrtMF8rCoMUkLE07XuRa7urRXjpR8/nzx2k+VX1IqjdCs0QlT/oj/
t0VzvszMzHzfyd2xJq3fI2Uj3K6+k5+j0uoFftVSgrI7tUasOJuwYd6Z+E1gWt7k
nOA7vE87ThjgYczqBzmEiRPaX5lCbafj14egnzXj/GXxFOyTsTurF62qXXBYr9Fb
gRLv/Gk6PFmXYt2Kvv2T8w8j/+fXND4wzqAsBKgEbouvDjgVwvb8MzSNODUvY66M
VHe7kXNHrMX9t/C580I07UbcIJKYEUDS62Jn8OByRqXoRbns7x31fggUhdxM0/PM
VnfrDVcTRQXP4lMtHqh6kbv/pji4J1d1U0y167C0BU0H/J5mE/3+iENsXlZbQsRH
4qRJVl4b7nAhAdejJWPqxLhRsoU2VXbh0IXTHeWks5Py1pKHmURMyxUnJQNV4Z7i
9p2UyFnWV3Kicetzvv+CYBrC39l4lOth5M5qjeLEjw6jJFEvLJ3LkOBlnTRBPQCz
VGZX2Rq+3F3/9XzeNST3FZ1KiEGNpkkC3Qmmn9P/pkzgTOIwKssKizScLklKL1i8
QhTTOTaYiSnB6jH1blyMX3JlGOBOep641BAQTiS3jcFgh0kW+9RI9vPpTuK2ophx
2SoUhHBAi2lPY+A/BPrAW/jCx8EgWTSbkBNvKGXIqjF1hQUcKjTP9qG71bG0J5Yn
vXrQSksp87/2MTNBQ6nGF+9/8AkgdACPEeQjRUrTYp5fmYXHjJxjqe8cDKKupGUB
Hu3+MUG8UBao8yr6Jw+GAkg0ciAU1s9T7MZ8hoE84Hforler7yvu85Ce+vsNY/2r
grxkI2Z8aX+Ubs/rDT7Z+coCVxlFEq7pYksSfP8rlxWtZ2/qN33r6RZ1LLSBgjV2
QEPm5cm4NO7N0MaLx4kkItcRNP5GFTHj0YdC0sdrzKM2gfGp+XRZq4IJncAr12Hv
K5EyKRiuBjCAd4INt6OmrpZARiqPT8wUdI+p0mUQgg7oDidAQb3vUEl+xgN/8dF0
TNrCiwOUMuzyNySKbW11+7X+rnyu25cHUlS+bbk4jdtta3NyTtgECzqNnxb2Wtq6
cfFM7SKiiaPLw00F2G06uhTWpTx/j7lrXU1r/o0tueYEmBR1r33T4qcANgKBJnzp
vhcIY2BtKc32mMnhiOPF3WHRYJTyf5og99NwV2/TbgCTIS9Rk/HSo68tmpqoacrU
s5UjoM1bN0IbRGqw8bgQt0iWrAJMoKV22qCInRMkdoH+G2a50ZMS7NHhQBqoL6so
6jqMDQQUTr7+m29lFIwT8IVNVZpp5RQX6yMiBPJWu9GhlBqPiUYXDRyA2f4wm7zJ
ikXoLnfiUyrpW6a9dBrn+NYTs/NIj2QenJUW6BMcpiuAC/n0aBi0APavEyxhiWqT
UHy1cl8Srq3nAfJqUfn2jJnWtKIXV/xFj4BOwuumPbxE/Xhr1JH9lXmFCRAZE0LX
0O5Qh9De7XYO2mPcpOya+yVYSh64lgPRhtIk4Y9OUeTXr2yc0jHAVuef8p/5DUD6
rhvs/62VqikRHpe3Quptc/riMVXkAqk7e1CRCb+sjVGdXAR/3m44AfhGmT+X1yhR
lv1Rt6lorzYpbS7/TTFTFL32UQB8ko5OAVpVGtOCennmENcMyFrycXVqi6usrBpM
6IIKZt/vlPfyj8Y7KKpkVuWKilfQ66fXqdS0DidtOrLEGVhO/CZhTw7qPuIx88dk
kOmCw2+5mUqC/Pnai0Bi5zXJqW48asVPHfUsaiDOYa25KopFospYnSo3iwLiSfkp
RSX5k69K+pkYulhzXyDBzqzRUWPgSqwdhqy2/XER1e31SmxMVpwr8NlASkxK2uNY
Uy2jFoSvDrve+TCt3jGV7N3wFlTPwFrzmzV8c8/NKpNJmw5tYG9/KI1T3RBLnANv
cirk6h4lvaqHOGSPt/eWPCF5bXTARDjta7HzTH+Zr5+rB519eg7v/Iht2HlgjCoX
VFrYAtpy5roV3AiEQHg7Z9QyYouGxPtLZ6vUsS7ZW2i0pSsGRIgF365mrEwa4jTq
UGpcEErGHHOJwayQJEiZjrPDy1u+7EIrxWJspYaIjimJrr6H86txt84YwaTcC5RM
Qih2zQb4sq9yARThwWWmZrIrRYTvmbqysx/qnotXBj7wDKiSKofA0o9W/p/12Mfc
mvxS1v8NT2yzXDuYb4NiyZlTnIkmIVUJnOz0RhpzOD8k6L6w5gRVjncVjN8iWg0X
mx2+ndaXPQvuqN693kgEwFel0fKnLbSglv5YJ3ppzONbyBb7kgp3JlIdMWAT7mer
RbbMfbvHNlUVZ4D1cLvG9VSiNuwhhxeXqUH9ZkuD9SMoljj04XPOtUu+QDPjgybh
G5QWSenwDWktvIxrBeD/x+/MixFcPLcBm/nZ68who/JEaYSO9Kn6yAId0ne/5Azs
sBjfHtHW944om/TIuDalsl+H1TiKJ4Tf9VBXwUF7FfVNRW60FvxJnhpS8ELD5bwC
++GH/djke5EDNHDowbQHiwzGxqpG3dWGxaZMsm6kCSKwQOaGIp/o9hNXzPz3NtD2
1R6ovdHmvTz1Jaq0pV2Iy08fZt/Uobd5UIYigM1sWDrXeq3HwrmjFlhJ8HR0Z0yM
omzRNhUi7FNPA5UX9SM9kzJYR7qwc0mS2LGy9IjGqOCUmp4oihD4jLyWZ8XBxkX+
bD9N1PcUdWITntJGvkQzCctxYd3QvYgB87PiXDo0RBhtze0muEiE73INhEzWoNAC
0K+1g1YKX+6sYUtASfFtovfRYy1MJc/UEtnYAwRKjnFR501CYuL+2yfF2B8DUAR3
UWwhR1l2UyrXTWkpAo+lBwH+3JOJK8kgPrBzrdB4ct6Dw/79lkEcegB8MtHM5rWh
DBB+v9V/fmG1oYsschEo++TkMFdGNs0uRn6y7/QMfmxUioXZrgNdjFHzc2UJhclB
iNaCvlYJO/z/LNG9RtoDmL2nLpe05OzlUAHLzb+9bD4uVZjJXs9FqNm/MzD9iwY7
HmvRKwPSt4ZH8JnTy2f+4S7wLsuMFWfhnhEFk9L9PjXcwcJaoBXpuIo23hFAh7gn
oS3PgQivEEKURTwLeMlwgsYjd1V6+SY7BI9L2KZH8fCiLNyuRIejMReZ31fGmWS4
FF6L0GCngH7HXlNSmsHwzAdSee8itSCKBZjXA4RcTJxz8IeflUFhdrSRVutzv5nJ
cx9/ZaCxy45tfqIRPtBtZ4b3bt248KqiIafbwFTKfWPhz3YVGLeMyMtvpPR0Clt9
m6xfy8GqHlaOrMexk35Pg8WnxFdukS49WlGyRHgHdHp7g4rDKfgPuBV8UhJzU2DZ
nUOZi8rpxib1JLQ+1x+BumUYj4Yi/JTLfhDpGm/OGUQ4QZR1w9qna6tT7+/mW9+9
DjrUx7dLNZIR40Umfej9gVxodufWOc4gaNLoPESJ9ZGq9/XYnjWiDrBhz6ITXGXg
/deHeS0OQPS9tnH37h0SeC5js/1jOyM82dBaprakEEITrUX48bSktsdld6gV4mkL
aWFIANSrM7o4VEqGd11ng+jUMUKbd93A9VhO0kJ+r/0hYA3qgkO1bmXM1d784Gpj
jZgmjK9x0UKzbgkYy/q0/m+6ihS2eLxPRn0d6Zp+VF4soMbYMjSiirvDtvodc4ti
iE0E9riKIGMZJ1q6IU6mFllNg3sC1LrPSceuusj8wIkMGqVs7GuWf6JRyH3q2sCs
CpP4AbCxZ+pKXrXmlAbLPr5KtSe47ZuThHJVG6gB/Ozro3Ak8Lw7/4N2zbVwKxA9
M3OD5Foiji+WezSmyRN1wtJkbrKu2+jT6j8KUMz8iIHiOSNSKz2BAipDuYpQvmct
goYSMtLsz1XevF1HPdsIc/NpZ56vLnO6mrxwdglKzXM06pOkl6x4dQNGIxloBqbk
fWCq0AZPsWPdPUvSRV9Xa/YF7w7vlDVLEMguJg6ZJW/WOR6KlVjPkiQipQiEQMUh
gRJAeOiZfxU6O/5s18tH/ka6YNK0xzfhkgr4v5pgFp/2QkrG0WC1G9zfhNxEGwP4
RUg/BD062eYmmzb5nWedNLSlcWvuf6sAfuXtNQXR/6M3n948F1d2ceKEe68sm9GZ
GIS35WP89wEqDDo4zoM3tw9HWdoaVOs2h0Lw0BJaKdGQ9bKsoEXlABdy921gfzXz
deXP+3FwP/advJSRBwmbYvlFPP4wnKO3U1YFtmslCuYlpehg7cXVillRvy2lO9lF
cNLaCWTKarmE8Icgf76e6K+K+ZOJ/bf+C+TJ/Evqy89TDbg+QsBrlsX7C/oSSwga
EwIcTzMSIT0qA9YA8uWBvigZNoAOhyIvDRZ6FdyMhuKISlpI6v6ymvA85xIiy5x0
G6rm9fRyqer68iA/yb3RLW6+nd2Yb5tYS/oW1Z8n0PPzM3pxC1v3xqxOSByuKSHT
ScmAIqO32mzSBK9kf6ihQaGwt6ANa5jR+2SkOZAQMLdGozup9bxGtjli+Z9xVpQy
ONs8T/HluKf0fPxeNZXCmxYAWDs4SYXI968saQW0Mbf8PUmq2f0c3K1Rajv/gUim
cf1d850U+JW32v/vDbW9mwGfGm2GUjc7Eu0Y3dTGwR2f6g8Iee7N+ShQi+zJ+Zco
mjow5UJAMcy1weM9zM23L3YNMrYyVsR5lsx9913TfcdsHaudorQcau7XQPHQULcj
DMGiyKXXv1wMZxvZBGyHc4R4PYB487ktsqnAbaL6nF1lwsxPmt+vC2ryLVCs1tdD
bBLW76cx1BUroR+MSoUI3x9Wbb6f+0pi5VFQ1TIpOYS9i1BbpM66s/FNrLxizBx6
lk5B8dUB1xiyBKRBh+TLcpaNVU1mKqiHdceNlBwi+qcRBeLXtf/gYEjsJunDS7F0
aT1HYTWH9XjsYmMFLLTVjXnl+9IwjWrcR4FkHAaPgoKVrBXKdjmngihfHw2IkRCl
DHKiWntjnFYAYbTOwVKoveVElH/jIN9oCWXDUVdSZgptZJCRMROunFLMXDgPG/yg
CN/YiCyd4HbvkbMC6LR41VIxArywj+w2fUrh546VKwU5+4AcoeEvbOdyk7Xa+UeM
8zLqV2SFbliYdotIhVBb9PF8a6IkdxBACuDU25lPSwr+T662H6ZWYAOin6JQzxnJ
GL7Q/aazRmfEUS3jJj/3gT4kpjUpM4NFF968t1mr/PBfm0SIyxPXtJMJgaQvVdJV
jLi40dEyi0Y8e8mPyFtlRQbpjbt9NbLFp2wKtTNmwm5OgE0p0PaP9OsvMr92vBuh
pKms3xNYp2mzk0kg4ZKDZbt+9JtGEDiY2FXeIWKVJVrdvpO/sSYfLPoOCQBGNLPx
iCRWgEtZfeIECBIre5Wo/k1oTy8Gg6M3yCU4Mf6ag4y3CfyehKwH66HoalA7Cuzh
l7wANkeBYM4JfjvqSo8muIMpknLGj9be/0V0exCMt065hqGBT+maM4k/+/GJ1isC
GdpvMJ/M982B3KYk4T6VriSPN1M4X7Vjm8OG9b/XAqVDv0ycoCjkmDXc/kiB2q9h
mGkRW1fDiXuyE8AluYelPKltSsB0yiRf5MtOn6c+fhYKX4HYyrSkKFv2xJO0kumh
haNsx3Yzl1u87AwOA1wX2pPJC16gZaAniNuwfr40nVGziuPokGEh4PPqgUUnCn2l
pAdrBe9iVCffp8nqPaPHMRVjk56+EFlqs+gZQNz0jdnVvBLi7Ml8u+lKEgOAVjdN
ir8nMg7Xl0Z+IAOGWZyWG0QeKWYZ5uF37BpcvJvxazf81tfKqHQez19skDVP8l0p
T3cao1XI8tryOJhs4pvJHGjTV1KWJI0sBlMDzjg5Y4I6pNGy1SfEDBPsjm/T1nSa
8MgSiAaTHHZrOShjVefVQZSZCw2MwfgOHXizBfu09KAq1osnByUWc9071T3gmaLj
J/EaCWX0rxD5v4rJhX00PF2A0IckOHGu5RfMpVhf0mNQezHdutkb+0/g/V78Dp5s
bAK91+noq7AS+aCVpqMRcRZnxEbTauUKxMXa5lg7NyY7JbYT8fnNlbxbi+W3OFQT
uYqD26Y90GiVxrXW8/685PuuiavYy8eDOSt6EDaduZmjhpfGNDM0bg7Ba0m/2W4g
vaVe0b5rRhPyLziY51R7+J53P1neSC+NVlH1Td/FvC9SFH2P6LfjnDglbg0Ye9RF
XRdnBxijCAee2dP6jmUAfBoCDgfLrjUWJ7XPyqx/ywa0/ztrqShfYU6iAhleFS7c
wvLpJ3EMu6w6D4Xh60W4ytnV8DoinR5ejTdfhs8S8uuBQHkhMXkIWcoHW7jKrlUP
DozdyQEVbTHABJtpWCU9DdlinJ4FMZc7YkX6IrKPu6k3H8FgYnRNH/byhG0xK20v
qXZhAiOitZeHQsuAfZg0X0TNsj1JOD3Pg/0FK7k9hZDMuFX/0VFBMzxbaEe/7bAy
VTKqxLKIewvyjiRHbHhW+awVUsfD42cli4UqCL2EJ8iHfDvHfkEmPaNi27HSwpoe
azKLzkvSIAtb5JdDiASO/nhRXQ1uFXmqDN49nQ+9Q3woA7cs9I4CKpT7F6jAiy0A
J2aA6iLQsy/WSmBx70LuLFLVHLd5axOko1BwtIX7wsmbF0XYf2ByJjTU36fAwj6N
1LNJBCEZVVi1lEWKsPlb4b0VTSXeH8nOeLS5v1TBjjlsDKkzEwCc4dtWLj2QJ7uA
hOADZR+FMD6ZI6HHQ5lM56du26lJQl73jsenBmyShlWlvTTOB9v309iBxS236qsI
S6JYFMYSAT/IsZ87wVsug/hbK/SwSuz+54O/OMbM0RYqSMvWcijUCWgbIZ7QlUvi
0ZnfVzk1dFy38+KSZzzdB1aY82NfSH5XUIY1lkPdqmSoZZwCURbI3tVtowpKIU9u
4EJpuXd6fCYc8Py8b3AvT6nsNHAum4yZAN2zWCxoMgrTI/3bxLgqWRmtvZvjoqKc
3s/1ln39gaPi9/rcDUB5U7o4OvklDKD6foAcFaEwcdKTv328a/4+j1sNk+iEizUx
XIbzaF6+aS6eAGPwl+UNjkpYpuwxjg9OPdYkaqC5ekJOhoFwHquYBlztyq/kyVgP
rcJEbzUWcniXqUzfscoYzgW7bjSgN7mvkN2vI8AFRxSe4+HcCbCqsv/gnPO1YlZK
6tXfYuMatx1e+WT9Qn97pdcPMexKciDD75TC4POBBxqvTEaIfeUgnR69OaSAoxAp
7SnK3O5Gc/YwES5P4sXkEGFmmGwXWgn7GK/JLhp1ogwoskXdD+LkD0++6XH31tNv
M0EOBmoEbmBlvvB7S5OdzqGjTAKOidxmkQEQ0MlOgFbf0u/BVy5l4YU7MflBH0e3
q/Rxq5Ny2cDDteRHwveNuqMrlltEmubwiZWhUSFiQTqxARMq7T5PqEShSYFRC2p6
2/Al1V/Ny/ME5FyHcCg06mRV2bq5lYHu/XHthpVqXmDi2ox9JSW/8Thqs1DjZgIE
SEIQtMp1lwubbAEFthCr4ljQASlVtgFiSW5XlWxQ6np/fyGD+Stz1wEsaoZVj+MS
7Ibr/mCgXRivlPlLOg1wY88jAKyqPg/rIP8NZvtQ+KaOtl5946etCJPyIl1D6H3V
f1iFk+ol/oRMc5seoOtlpaT2NR776UH9nJ9RF/PTcMJVhAMzKdudlQVHnCK8JjrB
YmTvjEMUfcTbvDleRUZLOwnVtIHcdQ7lbJ5q/qt5O1LoN1zTsdRLZDCksQdhFnDw
384gOSIKrdbKbUxhaB/nNLO8lzDGoFi7IF/HHZVN6M6aiyhhEeL0EuCZnYXBbN0w
9X5fWXCJM7pEqfR6DSx2YR4mfejmsBmAsh0roJ5Gte5ztsOUUSEQUDPQieZJ2G01
0J8Ofc/mc40C5DMiD2MUf5lUea2LhlclYW3XD/IJ+fhja+K7UD/XsXulyMM1XYY3
7k4gyXmIibj0zjr14QX2/QVVR72ExVEZ771bmEJHdZ9+T9IgQjPQB6ClF/FCz7Br
ymPfrClmnV0Yd2bYCKYnl9OlG1MMtOaxeeUWLIOmNi0NtbtQvAEaKVJCM6A7fD6G
yrWxlFTZOeG8V6JY+hAsqOeWxZOrpMtv3Qxe0BOXGkpHJ1Q10rIDeYxoM6g+Ep0Y
weOYTj+YJqfPRENW3VmGl64A2/gRrhUidb+P0jBRkgqJ7qM8r1OUtm6F9rDYS0Ae
W3lLueJcQdY2ejdsv/6fKIzjjFEnIgPaptE7xk3LyZ5WNfxY9NFCd/Zty6D6tkJk
+lHcAgDuWPJFLrrGrvlkRDvbSWqSh8jZqnIJy23Ye/guYEUz9eRI2LkG+Q4kPRe7
iUIVtk01vJqvpUQTyAv9d/hS0DMInHS4Nk+PHrr+X1X+68+v6rx2gj+LAaZpFMwG
TBGDAuwcW9JOngYVXhDihV99ywS1fAqGEGW6g1A9rreO3w58FKONSrYEuDRuzVpz
POX1MsoOrS75583/2ywpE0I3G7bprUyMjKuwnFHkArjSstdrrjAqzA4eS3WP1fAE
ib4BHqMiUraAB5kRNX3n9OhvA8lxwfhj89iK4mpkTw3TnUTyphN2BkFoPhuvvLQF
qsb3Z0N1s2byDq1iW1FbQoCIEcGMdnKLh9SNxUP8Ka9olzRGgR21qFxKi6kNxBRe
7ZASphpEoFjx2+AHbC2JEFWRE/ip6Mb+ZH9B9uZqBDH+rWaqINb6SvtOlU69cxAv
twURRE0Vzr+D7R31WEpt8i2qOV80n9ajS+MEF0MDsuqEi0IcfaV27/QoRuvxCAQG
clH7hIoVfYU90xCrTR5on8a9LJxhV1Z1gIioqSdiyroZWaLis4ZePP2ESpqRSNL1
EKWhnCydTBljG5eEr1iGaVV1x7FHDz4KpwklVNrM3uw5paJe4R2GrMUKjDwRLci5
zaEJ/XazLbKrWv7+IwE7r8O0wGI7AGvx/1NjWMi0ba/msgv8yJv/mPx6g5b3UWwj
NJGf8kTooObJQExW31zpwGVFas/IAYUQTmvni9hab+oGfrdUJAwltqz0MDkG8qUT
iK8qERn/SKaj1TubSp4/SzIE2XP18zczutUFZTzkjSMyncnWE1goy6n7l7cNmJDY
dVT/B2OAF5ClBsgKX1KoC1eoqjwGvvBWgodK/TYCZmiDSBMAjtvvLNuPbBGHxB7/
lQ/qBWRdZfNTRtawVnUhT5QuuWZ/MkknK05DlVz2ng9hv2ZJdgMuwyd2sCjtzxRu
i7q3B7JhCituM0XARIOXOSV7NbltzYFdqGVvh+7+++RnnzYR9/qpvS4wJ6gN3xKb
jf1K4Qs0QykrGUoras3aZU6k/rL1n+4nJ/C2zT1e+ot96x80NjdCHnvJIc9jRru7
JWhg1fz/a5B9KSIA6rcGm/MgQzYmDiK/7RdO30KWQUTuw2NzBpGkp4++pmf4dVCy
4665kgj+mTj7Egq77r1J/UGIeTDfM3llem80JWHl9+I2IjSH198W66KyDIUSgguL
EuHkiiW+D9NV8oF9Y1knvSMzYi3CVXzSMEXWtmVnkamlDc2pDdBZRaxm/keXAhhq
havoiYEqbibtYhMzkD2v6qkc2iIiJl23YhcNNK0oibcuEoSPLo8pGJ5FieWP+1Ks
nCaaV5E2GF2G9PhaAVyBjU7wE3kVJaENM+5tcg7tLEYQ0swefZSQtBXxmyFuOZV2
fffASPAlHVC+ZMxwv1OIQVOdsSyilB5mZUgkdgIXwdK4ixZV/QQ22Kt3fZp6pPbu
qn+x/swEfbKSki5xD1Tl5Xl4g8OKXQKYVzFSIabBJuTiK+IO17RiPblRn88+e3qO
RUp8GV2FU+q94s+aICLgnCX+Zzz3GTM/lBE0SAxixjDTKLT8UU8ID+/LbcgCWfUF
CmBINJpe5I95Zb0r2QFbwDHC8bgoYTlla9dZsHKzlxeNWrrsY0FGFlXPlCyJqhmz
eNgXEvbRjaN5IQRiXzvtPnvHsFRSHFlSOieOQg0BUsKHw0H5FKho7P60Tiib8VtK
Yj19AuA+h1mJjPt8wT3MtzXGuiU+2jwhN3FqJ77VNKwDgaqQlwDSFTjYxIqbvapx
1J5drZmHcLJ9j7sNjz8SuY3obL0Cs0EXa3YynMkpXBcEuLcJsaf59fL/Q5IRWiPZ
zqIUZyQk68QSJyLA2+9H7ASiaCe+NHYqNILBAoFVECzp8NozlOFkLSpV06DrLCce
IknwDOuHY+x+q7bhZBjSqNafA/8lPtghkoCvhyuVcm93gPKXKpK+0PnF+Yqtm0xn
AeqhOjN5jWGT3IXoRCJpIq2caMyqdR78EdmHuZopc9b1OIBQWlfY2bQwL23/vktt
QlxnN+tA/vy+Zmd6V1YrGQRj8lo+FwzTjs6nS7k9sWj2tLleHhpQ/pikgZVi9vNh
c9nbBLcAp1H2WNbBzkLzuuUkIhGaHxaMY6Cwr38gLeEXwoN9gKG2+VRoaidWban2
NEXyzKRG4FiX0b8b/rlC6mCPZeZboq01jJ8l8iX5P23/yjl/u5gojY9f2lEiWKs/
AjQQsL0qGwqsBq4lKkzsJsXiulnKLMPGf2QtHZNHq6Nne1BsLdaQuWUGPkM6MbRA
enmeUFhk/ql/9Y6rFF3EMJ9juhf3ssaoH1Z4mUZReJa4T3aITeA2eBZSd5235mef
F2+o9OuOlgdfXcd1txNU0sBzG7iiv582rwwsZmDuGGJiSuy5exORYcHGW21Rwt6R
4ECQXyrPNKKWt0+u9edihgU6cECgLgtnIfr/zq5FpkHFd6PTKrCKIgXYWe3X1/nF
qOZj3CT/x8oLUlQlv/eU8y6RMOARN84o4TYA1mghwP0xtYf3oy+7z5Bjik2231hL
3nbwUg0jYAy9NraV/AarOKxPqOeyzbTcjljgBdvl5jHyHoKizHTNcvw/OOumGg9Y
f9XKMqlkI/78OJKSaAH8dulzbxrE+P9VERs6L/4kMF1nBrWYQMy/R4DeQ9czq1b9
Jxw4F9tjFATpL6YCVkwtDKr261hw+4jzdOKm2NsGdU7YSweOOEknoJUxW7R80rRY
91kzOBpVxI5K91ksj2vUG3lPgb/YJFHAus16/Mqss0agxv6qjSIbcg6TccO5r8cT
tYsVYkHjPib67tpD1jD2uh784ec64yyPbYoWk2vlvWBp4H+3oqhWTlAbnKi0CV3c
pQfjfEnxvwjrwf5pOQxtkrn7CINh1w2GikSRN/ZOwnmBW+ahPtc55LdgW5en8slr
G7TUGaT/xn77S+B+USe9DmAYsZn6Pj1H/7WoO/MNKz94RQUlhPCSModIrW+6zv9J
Htwzj60sryXuUFqsUPhtpEn2vmcXIEuFNFA8nPGTEeAqXlbX/NnIJ+0d+97m/YkP
20ilDBsqIiOJxzNxIxfHVFfIs1Rluyh2+asbCNynSrjgV9MlTJlQSj2efDO5d+WW
C08MKE6vbYZXQeldTSnHW+LvltPyCTBiqtuTbtfnHMsKN7VgqkSonNhVB6JQCoV6
ZYGrob/0mjyAG4Vhe/ErTfXfCpqEg20kOnTSR3jM//RYLOEifBKq9PkhN4d7RQ48
aSBEbWxjBvY2IHd9q17XUtVmVbcd7rxkzC3fiKvJ7pSDihnoJHQUOgc/IK5ev94V
4pw04YAjxEu8ltrkwrU6d3Cvd5Lc22+Tl/iA9liTkyhG6pi8FolrQnxf7aSSWL9H
QulyHoXeo2DFIc6vRneGXAqKrASlg4xGL0lXP/kJmGfh7NwjGelyjeDpJf3hz0Aa
OD9ZISgMxIc0GalQaq7BJn+ZP6Yf6q/jdvqta0iN5Wq/pvcJCmDvvukqax9ImsMt
6S6gQXS9SUpZHQn8cev3O5z945mMrZIf+Y9XCc1dv/yZ9Ma5Qx9Yyxi0WNdPjwL+
IbtY/2CdpstkjFY4UTuUJaAPSQSbXKLNjV0NRAd/dg2aoeCJjSedP2Tod+wCY0qj
sPlKSucAkF5jC+vudjEKfyPGwfpgEsEF3ztZe5rUR93IsnLViIviCASnjAr2I3bG
UHokbaY29BqDojKwFuk7nhuq/WOdtEXZPjHFJb7ehxsa6+Z//r5oLMAXHzBK0NYq
nOwItMjgPVtc7ONp5HDnXtPh8IOwE5UOUThA7YSYotalbF/GPylqBenwwvaYNYAZ
k6umaWpkkMJzZtt23OHW8Xln7Sx1760AMTFriAoxWnet9h+jRfxu/UvgYKHPolKx
sb/3tSXfTS1dUgEOlm/CXf0XOxOKVhBQOCyLoIBSY/Z3U4WIdGTvaj4w+anPRmh/
8WRwDKD0apuLHNtN6valKIl/2Nw/EXdnu1sFUA0P2ipRa8LSpP9J6jU7xMdfGsgt
DOMe0d3bewHtQ9oQX3LHgEVUkGNpQWoYkKZHZqY5TSOOarCVbPk7agzt+WbzjCDc
YbKVIu+1EM2NptLOqhTcs1NpXptOFFpgIoK+W32YeAvlp3QWo/Xcx+uZV+5PxkG0
6iFb3EoBvP1tqMORCCTP95Mia3cPPloUgD3mHJAuc6T4EBeln/5tOPiqU7YqRqsx
KtbEBL8ymPOn9W4w6QUXjFebP4ElklWSnSWkb/0zIoBkZBbNB5b8jM7NoXhdp7vG
A1K+t5/SRlniNdNQGmq0CUoCQsHGVj1tzGaxk26yrLUmBlZXDQ+Jy0NTFl2Sesgi
EWsRK9RWf5rYj3NLNCRAaoIm7IFdkRWmp3RrPwv5sqNDsrb69nfGMmWk6XgWPNOh
/Iq+xlVPJGonaj2Fh20zgRD0Om3kHRLVa2wQepOavGaiZ8xjFSEfIjssI1zsjz2f
Ya91PUxQkkGi2oaUGNryscbGiEMbdAqe0YU8fsvwJc2gBuk1ylMQrNd57M73Wbsw
m588Fwe/rDBmba4woew0cOdseW6XKFv2W75+ndxgkXXjc9NbIc6ZY1zmlmJXA8DJ
5+4A/V0O4i22DuEZDNbK9oZiK7t5HRl8Q16loLxNj32n16m4KUTpp9dhtTC4yEfX
uQKqyLRHVUG4XiRsE4OlS5JRMF9cBMm5S4VRk675byFpVVgXxbnr4bQIiiQyPHED
0EhZw/VN5zqTt0HSiGKqMZ765vjytZEp1zVfKs2n8pvXC7YrjiRSkzgqeuAjduFC
8jNSmfbmZmUVYtx5m0K2tOv8MH8DtQvHQGDnGVFLFjKT9L10qs6gGnQQW3cUWamc
Wz2arr6mJGDM4R6w1n7BUmo2dU+AgQXVCH8yClVMB7II8gIg9tC0IdFxh8Jgzw0h
15Z2xyajjEwDV3PkmA7/y8QsMgFm0/0yHzDwfsd0yCLBgjqAAGSOqEQuS2M1710i
UacCGqd1/DzthMPtZR9BNp9oMw4Gf9upm+/H29gnSt20wX+JnjjyEqX/GKiqVZRL
tsK3E8fgeQIC+CylyZZwPAK3L/WFJKTNcRXz+ihYUXeJmD4/TDv5+PdhPWrE0IIH
NsIwf3UqgFJLmZJNPmNsT9wMkK2/HuyvrAXhUt/N+tAt8Ob68QcqKaB8R9T/0B5L
k02JTsr45M776fndDM2TdGUz2ljZybNpgKK3gG113j3oH41oDI7hxSDBon/giFTl
OYOCcl2HZWsSgMi6Ti39MjcaUAyhMWagacwNiuPAPkIFaq62D7OXPkyLTIWKzzD4
KoRIQxay7TO/1Vh0dIkIBmFYUjmVeR9EvOyNtRvDJUyFJMJo4gYMB6AkKP5IyxQk
ZR+F7dejIPWMmCCSsx6+CcSDGBlecoqdLGbU7/8mYmnc2eJZlH7E7CCv934ybusn
2ovFzXyzlcAnLF87BRhuBjopD7ZTAUop3MoliaozLBim6DDdMZRUowMtYnDGZsrn
H+dU44y6zW/mPZYUVx3TmEYDD4JjCgTaw2rKK+pZB6E0ABWT+/VjAniJE5V4bwKF
MYDpPr9YMB5BAZ5Ok3mRVZZszxCeIlymmTBiG/B3PSg3fljVX7BrleEBktTI2hx5
muRz9jPPhd4kV1zR8GrcDoa0k5aq/9NuxzMhut+n7oc4L36LdOcGymA5B0v50rdI
fNY/DA3hPzBYPGaHyrN0UKKhr0PenBez9ilAb52RFgFs8SESEBNmNkkNYiSecOVG
zGHMtJE7YwNydALIXASD+FZMEzeMWp7FXQIQnMCQhxg+R4YJQOAzwxC57RHrPkZb
esuXI43S1fcL1CG27UThew5yGe/sk5UKLUNyPZdItn8Fs9IMnWmHpM1fcovAMuof
T96m8CDfmHRx25w/z6oP7rwkA/uhUNFsvx3d//PNNIANUUSPk9Xge6mClW2ZYI+K
q1vkKYhDOxhud01deOQ/TUKtPTy9bqFZnooeoUWG7McRCYBYX5vugu4Y7JyEfpKA
nNLXGEg2Aa3EydZbZCQTYY90kgaUWN+cCAupmJfMu7csEEBwzGSvIiAStkA1QilF
HplgA4/9+TXPhdyv21CJgqbWnNc5E0dS1GIWe5GkQz1uI0R1MJYpBk5kGq8T1Z9u
y5tNZPmKFM3cEIKaIOe240dF15Gjpm6tR39XFKioiIbM1ucg2+EQnULsERHT0zhG
X/Tnn2FVjqFv2fnyV7f+AroNrC7M8rqcBaJgjFWr6hLUDtT1AU+hLIqGQPWRyDjo
cYWO3rYWqw3qwicxTkfHEUht/v5p/rOpi3HSlNhJk/BE2iNnvyNW+FQQNV0VaQrT
Y3DLgH1HagNYN92D++GyPyzKaeIdGWC4q8ai3TykvAlpIc6zlU4dmmWkTUaCf/sG
ANqRvubvnF1EbT6N+IfOhYMqWUIkJQeYkJ+3dkNH/4i+172nNUiYl0nFtjgWAbAe
xxyv1qIkmvKYY/X5JTVi8hpPeWKIjbb89Y/1k1RL09LyugTl1vx0XbZgy9M4HLjE
9of/mS5A6W9tFMWyK4K2SGuiAXWT5vPKcydc0JL1CbvMGc5mHRYcyxfe8fW8xHyh
9JmJxIDFaIFTyzF7t5Ks0hlLKWKOKgFRiSBXMk3HHnc7ezXpvznXp3y8ebRgyFeB
mV2WnPS/wDfsVMHyNHsVEXdh8f5V0nADRNvB1EsLuqmK5ZBMcFz8Pgpy4j1JFR/z
ClpF/bJ6unIM/2MkuUBTaX4cB1GNa4giJgncPqPA483jwiqcLrx3m7nkIjeeL+6P
svQv+7+w499gRTeglEZxRcOHua6HlbAacLR4iWIqLtI0hSUXMe5wp6HEQpVEPHrE
IL4Dkzf3li4edTWScDCTqVOSwUvMORkebNXu1tQZadOBsrviUrpIc7TFH6XiTN5V
xwOjJqPPreSTkGwt9V7zvqlRzH/qEaiKwQtvECALTyaaQxlsdOgvS3KQjCrfH7Fr
1cBmHotlSNJ5HZZl/Mg2HA6IThdfltCj0ZVToTA5WzDeYpYFnr+eAS9JfCuVNI30
Xa9avc1Sai4i4PHlXdZCS3HuCuOL0JU5yFaEH0tS97Dh+d8PFhNH8lPM7dlbApsH
KSOrHg3e9jzgWfl8FEYK89Svx5By4F49bpXSwmAvZg4IBY6PjxS1SRhLjZ4YiESJ
UcIsBcm5XVXtuYbWadIPDhSbXTSJmYsZPOn2JG+MAvBzSt8gLFBqnXtk200h2gX+
M352y7ny2kQDj9afHWwrxp8kYcRTWxDWNQqv3rFW/FQd/Jsiu994nqLJq7U00xcQ
UUioDKzFkMq9dL/NJ8Y9zK30sbE/6Dkmz/v7BMqdWlx9IEJqQx+v7Dj2j78XlkNX
t+TUM/Mw7NuMRZe3g/PSiJmHcmEj+xkapU7vR5IR0+4RKBfQ07UxlyWwfvE6MJZM
mEjW0+DzIKl5QIzJnJfkfNJybILZoeDAT7BrQuAKvrqz9p348JrKqdg8vrIe43Pq
03Nus7V3/pXfz3U0iEK5g37T1SPkFa7eqGMpRE5ZelPV8l1v6cKS36NxIlGTXwbS
AmXv9Fgwswf81JdeIdQqECktIjhNBR/8IHgaoZb1mEkvXa3jR9EyLlS2zJABlvv5
JGSZSBcKDBaTr5fn4xY9BvtkH4TuswljnQyhKbEK431LI/9/2W+qfyzDNUtDsErZ
8ptWPY6iYw2680SzemNPozJxwK3SBm2sM9Qd9P9TOF4FG0VJJimWU9lKcJXKSklB
3evtEEHgKei83SAYyxFwMs+K+4HCrf1i3vsmqP7Gna3gLnGRGlFlWeGwu02ervAc
+ccNhbDLq+mulIynzQU4lbIfoo+Np+nZxXfx6cIyH+LtirgS7svvvv8XYUXRxuWo
RxpB7yw43KuQzWymBYlQAclxQhe8B1F+O2oAkWia6dCpX9nFPdlBcBKTaRP78Sge
5qvSSTe5BPD2nvAfTXX1z1ttZ386f+mwjaMn12TeyoA6S0lyvYDqyjpmvohsXoXR
suuS2Hxo1GOZqS9chshJQPpAc96DBjhSITWciFEA6kFqKWZJmD7CJmW0xLREPwxX
rEqbIBHkX3uXFYvpL4axt+ZZgZtkdnKkONFTUE4uxvHbthA/bDdCFJjyrkQuehH0
4O8WGoRzg3+xgZGf7CQSoeXlPqVDe5va2PhifaG58LlQU+HYVdd0x/DSKE022mNz
20e6xM9Rl70HZVDMnUE844XK1jJBR+sYWE13dDiG8/aqLsY5iVz5wn66ZsSzO3MH
ZXBlVNZCOKZzuVsiMvKUujUkxwHFTmJKCsTxwO5ThUOsmAVtX26kt14b/NPaDPr1
bxE0okOYuVYFEe+H/YGihhvMa1wJyZZ+Az0ICyeSQWHmvrjIlMuMVhq9Rc5/EtPD
upBZORnUW8Q0aHDcpqeJTTy2LipN/tDnYbUOT3xfJB+ecMpBfWDGO+UYsYaZGgT/
GH9R9blS7nD3s1bXXnSDrZbfmqLcejKHWa416EWAfH6WeSP6P2wZ+JG5DocsXINa
golYfDJWmo+3KcPS68pHZfi6i0zFQ5lggrW08WJmeo3u9MFFJcqEP2SYsEoBTAqd
cvsK2fD+q5b28BqH7hph14vu4jjDioKZzmuzdHPTzLJ2eW54kilwox3O/Rx2SanD
D6fL6UrB96883Lj7B/5Z5TKHGdLu/qvYwx9kYZOUmnQzJ04rpOnKtDpkR3Y+m7Z+
PiH4iBJeipDmAeaHPG4MdSJUTtWPwIQBq247xpIo26c3GQRurmbpWc0feXZlVHeP
RjiIWI2H0RVFre94F+FkCOuI+reUbIhQtWasZ8GrOy+/NT1O/eUhtEfdlj2qJees
RUOJm9G0VWUW+w8EWJVQgpEuRNKZLM5+h6LNG5+xuAkK8cIUrfpsiQWDU6Ewgw3b
4YfI6a730GQJa30dKfxqeVdXh+maNSZ5p+Fi6MA9Su9Tt55haGxEr1J40CcEsGUW
uYKekk/1uDcaEeSwsrYlVRQ8Y3rxNiNMUfqeHXbRUnEQnVXMKSzS+JGBZoZ+0pyq
YI/amrJJvaN5dbuDOHzno/mpbp+6PornnjM6dGXUzYB+qEpsk6qLJDVGezO5ay6v
r4F18uMo85rh2zfOhUKESRgIqmx0KnF+RDIvnF0HIWCj8WC6UwzasWj8Dt4oq4o4
B1bNtLmUReELPKFujlPkLxTSGbEsMAjxpGwSfz0SlGLynjEmIr3/RIKjyCmxvxon
NupmlC1/ZY42Trq5rtpsUcNRs+vSGUctRpZjGi/IYS+I6oVAuuV+kweeFVTbIskw
PZMwIYcBjLhBKk8xoEKmObR/hlL0Uxc7LZcX7G5uRhh3JeZs9xcNerT87ROmcU0o
Tl326U4VQsGVtOWmIVwbDUzm6ttw6Qa8Tbiyiw2UHoFWn6on5Gy/gyGJaWB/4V6E
xzVKJraT9++F6gkyHzcmCsEBT9I4rhZ/uLkraJxEhyiph8RfJLrnbQkxAtSAVSKQ
j3EHuaoR5Lx4Vn5CSwExLilTR7iioGQQWD2x1sImz3a7miUx2CJtYZB8S6SsqQo/
7BJXZ8vE1RzESs9CnZgBwnSfI+n2tcoSw6/gxMJNAHpeyCFST1ZtsiW3HxE70PXm
dvJhzdHM5VkzexwyOfLlyFXK8eyfJMAl1IhbOzslHUh+9sDeBoNBOYzKRRBzloVI
6QmDmTzSGEDJldMkDmkY90W6rEk9bij7rVfU8VsJCNM4XaR4oLbj30Djm2tbqYL5
N8G5TK+b4AdxmsmlTmJW+rXDE0SXuIX0cq9KAG/6NhoMsUDZTPfyJ7NXl9um3YKX
kdt00O+qonCoI46ByZT6h/QLw7TBlKowBRaDnrk1swTGpZKJvY1vjTOGQWG2g6nk
+tWZuH6oJHw6sTZvTYU2RbkTtRnVwQSKLmsyZt7iR4qKLzVL7in0EFpLFpKkTM91
XV/q35pEsGWdcIhDYq8mG0HqHbQGXz3KMbcKqUdNpUBtv42pI/d7Zjh3aFKv6fxY
XPNqxP4fyTpS2m3eAueWi+0SFjYp6dEcVjC1KyYgIVNhOFAktRX0VNBG+xPV12W6
D9IeMeJOFJrH1AYzxGfvjnpO/1d0SJP58rAM4VK/1IxsyGky8LsgEbfsoMGH4iQl
bquGY6G0Fc+0l1ycN778Krf7L1QgMAeKOtY6gA6tbZdYpYLd32fgLnEO+/DeaE7Z
ZLH0ekSo/g4I+5SN/02YPq1jngQokpmw7EuQ2wNDKoDIPN2f7icolUGw9nXcntIG
+9N5eO1oka1M7I+fx9rEp0gD1kVaorbPfHOLeSTMiCICx4mHBW9abspCx7Sz7qIJ
RGBbhpxtsdtTxmnLRQ6HNaPhVDhWgi2DoS7eyUUD8R41ElwTtXjaGgVIk0CLeFbk
PIyHBfPrvAe+SJIW8/CX6l9KPIs+9lY97rWdehfqhvQapEUoCdOxXCH0FAuSzEUH
mlCzZ0P+4ys9Ewry8JdcE1QlG3UIvPzD6hDsJtMKEEe8Jn3lG09X82MOylSHsv0B
cwKQFJJwj7XpnIaCyxfq17bM2uvwQXaQ5hhlpMAuxk4qfIHHn66LQ8z55NT42AYe
RqHpJEdpyJJ/kHP50Y+yNaPnVYhMhzWzaFLcKd0y2/sIcmozc6fG25oy0YLpx7E6
7wykTDpEYMc0J/5nr3HDcgsylfwUryp2lQvCVDq8DngVshutfp170uynv9P+pqpG
lQx2uAHPFh4jDnRiC5GxAWuU3BqJ5Jedzy54zJOp2DsywBKrKFUCWxROYnvbelmF
7yfhtfX2ohY3e2VGr/1SJtD7aUgR9LYe4gxZW83r2V8leuNy3AVSJ+4pUjUBsEr1
dLkoqUYS8M2jZARtKXPPz1Gwq63PNeRjBevVXRlPsfA5S/QdpV2D5CbgXipuCo7a
Tv+Y+vDHGbDkl/KGNQSzJ+w6HSE2KQUltbDUQR+hqD0OQutg85x+8bDp4h6D/R2s
UHO3RFz0PK2P3WbiVy/knYAHqpC3FbBKYpXcgprAxGZhDlZMF7/ASDHZBJfCNwPD
SST47hzTcogeXZgp+cS+/u/fNrn0NJ5jB+kKQWD0xxf1W7aztz/ntGfBmlUquPrU
gPLvr/9YGhOZryBKjnqpAeov/9h3JxZvv/3tDJbtQ69I7bq4kjrGiIFYJRz/1rMA
3+1kv/7PUGwN2tFA0R+d3CT5i1/kVO8c//5AUhc4dCHcyvUBP3Qpis1Pa0db1pPs
DLQKRPwSzkDaqEHd0Hsm7+efLKEq2Ggv4vispH7P2ZXenRthp6/7OR20pCTTsaBr
nOhtyUJxKyKW1PsK/ARceVCpMZjERhlUAAlvHs/SEJf/VnWIHipGYH3h9QdezPnr
cq/lSbAk7KumegtJu3fIJLpsbGO9YFJ0nPUxEjk0yjlyQLpViL10B2UXB/+uCAtl
jh62JRtm+kJw12/SvjROCH/G0V+T153gOnC20laEEjxlFnoMoPAAVAMYj+cXBvLl
ssZhA/vRDklMpbWRqFxxyb3BdDJ6CUUtakBdEQWtXWT06YTnt7AUxPKdcYqQCGG4
JRMOYk2eylTPdihwRg92wkIAvPx5HofoqUjAfpZWXb7RlNE+T6StYV+qpngZS9HV
ggSEO4rSr2tuFBrPNbKv5JeNqS5UOzCPHKuvC8YFSo2fr8ur0N1Jmvl73fveKCD8
n0LO1V5mJj/06pvj/5UAPhIDILYbidg5aV1ftywhpuf+HpByybLF+JCgNfWiI+t2
CHSAwVFd3+78NRM7DhJBOPv33sKqCltnjQZELch+bwvd/POTQvH7CujdB5T9eACQ
1WNpPX6LVLOtjdQrzHadaXxopU5HszJbmexKPVpUCZt9VfyQsY1+kMoODwmrqtL1
HXORZkL+zZ+CIVMp5+1GLzgieE6G3Tw4DhPFOeeCkBPbuuwjBpUCHV0prYVUwrb4
1NLjRS6+EbOqrgvqS2OCO7dc0I6GgF6kFGRKJ2ChiE/HoE2kaGhPp1eF8VhU7I/D
vdBhIok81vZt2EimppqmSFwfijZF/BmrfJLh5tfiOVwdAX+cA58zR92kYQg8q4/C
CPRMQn37Y5Shyb1NMpQId/4+Rc5iTu6wvON5gUT8BKWM4xPy0FUA2ZvWIJPiZHzP
baZbKyUwnG2Knfc3YFbS2faMfyo0JPxg0jSOKapIsmev9a38mMfgQrzytGjt2yOu
/kli+q50qAWp16fSEOBpi+rG26pU9hEhoa7jrR9p23dhHwdIlevOF8jJNuEQr9fQ
DT7kRsqcrz+5sKUl/fD9wSxmQRedraKMFI8S5Ev9ATysSvgT2Nn4mGvG5uVFGXN1
8siOZ1CBNCcbFRECJvo9zf/tMBWAc8ZRPy6MiaBqvxhOumlxlxz4l9OzLKdKvarr
M223FvrHzO3uEJXO7JTZ4P9pC3q0jEZUY/WPPVrxrW6jGTplSBbCYHvzEm59ESEY
AMN2lsiT1ZRrc+n8tC6qIo/Ug0bvGiL89s3UccYoNRFiOuSFeP3FlFXi1rYmLXif
kV+TUtkBA4EEpVnlEUynDDlbqxupZrHtgBwzL+r3aymDpbpW3UKSB1KM4m3Ukca1
zcUlAhkeWYbALgqn39LVEAynkUiuuen3br1ldzaw1X3Kd4UsoMs+IK+DAfJoEjgm
XrVtowc8JMcNwMnb2RNnoheV2/A0GcFftdoZ2JoQbSwmtykChP4TuwyXnXxQGjS0
wj/t9XMQXGqGBOE5vhsBupNGRczVSnOglgPb+w1urkbXrCir765sumoS//nZvXeq
HCtD0jn2JaiD2aWlVKjHRvzhapBnRbFcI5vr66zO/nmAvY6AYmE1e8ZTBk03wnza
X8Zk2LhGTHbxnbtG9Lj7nG1yryF5gzxIBGfu/+d5Zny6RjCLL9Fm+taGtddR68qc
HouGLAxLxKSNV1+V/xMLr7kRTX0SoL8/Z38Mtw/m3fcwFKcnWoaGoyo5MFAGwXCZ
Z77cFkCyrotvyxi41zl1B2Lbzvym2Cf2jFGmmLFk3cCyeErxWcStHAqI9+zGvMjo
0ZQ81Bc6q/V2eL2UaZoEZY/jU0nsDbTQvN4IYS1CQIesqPzZh3Tz9VazphmPavcW
NYOsHlti7zfC1fndgK2RNU65fbCIisLgF46vpY9rev/Wmr55ViW5JSmOzgfZW8ZW
CoI2MLruU8qFBQZzsqOu3lRX7buPCekJcBMfuE9bMo/XhimFPwluHBVZeL5ysJmU
5WATSnrotOdOahqMyBJssr4cfHyAT1MTM9TcXlee65E+sVAayNq6/3Xm/PCJC5dm
DACOqRZV37KPpASokedLb6yoP8tTVUR1tYSqaR4f15lMal1IrS8lg3I4SzVakvG/
5+4UEC89GF4KeHU+Le0kCy9kAlKjQAy8U8SIGkEUv8ljBwjxwgKi/LMiECyKHTwL
12a6AeztlLq8H7kVhmUr7Cnt8h8zUp9L/eMmCOdWISo7JncqiYud40DtUgAjKUEc
CLc4SIPqzQtqkZ5viNNoyCDqE3fc+rB2AbEWdiTKF5qrcCqiT/5nFX/6G2FIZQ14
RHvl0E/yRTsEK3/L/rjFuGVnkLCX1t+VzCmFeVHi56l4gJxKHk8vqUF1LJrfjslb
AzlRClAhPV8rhW/8r0ePwBEbC7NHMyn3zp2UqAWeJofpXJeQ2NjWEDw6aoWAVROA
Bq62mRP1idSHkxKMyNNM2cOhen9T2+4Jb85WKJu3QUo1LouZ+sBzMa35ksliuMHf
aWjd9e44Xef/0EERDA/WllOBGygEQNYF+NFzUcRHYxY91gG6DNoaAKWmNv1wF3Aa
hRQunxbhZ+eVSym4JvknozNbD6DbXy/clZ9awqUwE8QoyiFOpcj8zrT6b/gg0suY
KkKErQMV+SoEsUGq2lgLnciQ5829LSUQVIvra1KhHCD2vbnvkphAQp9C/Ol480SI
JRf3dAJvJlj38fwb+GiPIB2cExZKtl5+IwYFncdLFXzIfrpsUaLiZlMZRKaeihdV
BXwsO87Im8inrgRS1pX3ZIQCLPwr81nPnRr82jQvorqvmOKcWGRtDefTw0ute1/l
ZP6yKOxUJrXptvPfLGWZKkCx5qAf/IXoY7MvqFuEYf3glMEIpmQruKIHLeyit0nU
ESYSm65aFrvCQHkWw+XqE9FUadXKjA7hwVUpZRb/Rc7c7q3w/hbPUXz/1ROoSn7H
vgWU2vblCPptQmoQK+7vUEY/M4L/IPnurPu3pDcPgzLvfa6gYjgf9/Ajcj2hO73T
7+Zn4/KhelOHUk9zNwW5/8weuM1pv+90bes3yDXgEQJCrK1ZXwrmBUiROR6hMWB0
Zzywe1bkUKYduzcyhMyhyU4cN0iJK7IjnsSdeT27WG0k6s4bhK5a9wIu7JsMJpAi
jdru0j8R1dtx0R5P4BQj/AAv8bCzSKx9lCLcFINj30+dshZjP08/W4qHu0+4KY2a
9h+mskUo5nfdINn4Pg4ZTBS52nLtPwxwGEiwJWzoM/YMF6pKWnxwVZpF0IZTNgq9
6yRi7n+5vBH+7u0nzwlIH+dt/gGDTmMGX7AokkWviCmaPF/NV700bEf5/cY5MkmJ
oSsQdhsQYs3yByeADA/JgUipMLDaNkovh6B/jfBuTvI//IfNTRZZ33MQRdiS7lPN
rFUiC4zT6obIZSh8M4QXkTJtHhverB6lI5ryiQbN39slRh6cEI/FyWUMMJWZm4iF
RQIoukXC7xEysRyL+LUJx5lpN31WMnWreGwDgpxjf2S2qRR5M1nRp5Zy+JIB3Nzk
hD84fBUWrlToqxPOjzWv1AZ+sHxIjlMJ5gwMei9xG56lzieLB7+GFCBpgHzCepYA
ZQGXn2EbZUPpTusCvRR370PkwHXfImNsaWxsMApTy/ibEnOXmvuzyi4aU2KhVITB
U6gc/4+2U1gP+auMEMODnOntvJp23f+N1GFKTg+/U5ROxXKDH02mtxh8fIkEcL+B
F7ff7tr4t7BJ7K5QkId1kYvMPDVCwbxWr3T9e+Y0j5V+Pm3VRQp4gMa1Y57+42ko
T+tKkYoeOXKH2bG2O2S5gV2AKoI7DJy/hI1J2j31lFmeMjd0t4PPeHMr7hLfJnv0
NlSuLufHs158PHsExd8oVJ1rl6ZzgEpVZlAOPAtEuolMnDW5J6gQlg8ff/e9zJA4
uSF4p6W/en8RewYxYwgd+jHIyvRqoG6qQCzv7uqlb1JJbIWM7wYUz+2GCm28Dtrl
BVDVe8hj30uATazsktYaNoU1xK4Tv6fW5jJErbYnu00/FzSZ3/emsGy5KTuwwsu8
wu28gX9ibq75bFUk4FpkTuULHyVuQB4Ont5DGti05cejD1dnaD9ki8FvRNkbvKFo
eu5AJF4go+vVOJ+aeOqSVRgofgkAJw7/Z4p0ObEfx0gYAoD1cVkP4vX1UoTNJ4t8
3SACbXNsArRmklJkcbM2hDvD1YFLpo1aQbXPyhL6UR/Kh9aR9ujhBvtmHqsfMbuf
Tc9yNCVxq++mwQXSToSgUAyH0jIO4fCgXvDlJdDBKwUw131xn0PBfN84+bd9PeQG
9SebPKfgHk2bPl+kIFWdwhdsJHJ9FdP2vXtFeUGZgHSq1bcVZleXp8NjPrPGVaI6
3n3pC43suMfPBhmftzR1/IY4/Q20NPC+1OvvIsyEa404lDBq+d1Y652V9oU4aw6X
D3fca3yxHFhf7bUcocKaWMss/NXWFAFLczuEeCgF5a0DZ33PWyZmaxUc17qqQ8iX
mSBgbs9QIEkV9n49kP2zjKbVyh3v+3I+1g85mWU+4z1t1PkMobjOfhVTF0Q16aLC
PuDkJkIwFPpyGOgmnjKHFWAtyHOZ3EAvOOWsWHWVRoHFGn4tkCzkkT4r8T2MOgGO
PLyAOIn1yo54Uuvdf480+CINJZfJed0GrXRAaXICGohQCC8U/1eaoPKlx5oiUy1F
2Y3dq5vMTBni5R7OmxOCk0eP7JS0sVw/ng1DFGJGdie+1Yt450IA5WFvxzcWG5zF
TWsM4qehI9lwdciIZsad87SHObQYkAzT5sPU7U0L0lPIXXSW2hfV6MweYchw1apD
7z5pGD1bwxEsokQMCYHaUc+zfJ8widDkqFs3ZLKxYtyaj77vfPbYuvl6BKNT9bqD
LAFqmPkzRoh3ZgjAna+ADQZvmsNeEA+nElayv1NistCtgt5qnIgPKAnSK+cpaoZo
TAEAxl48ycWTrG4mFpFnsfIO7ZiK2AsROO2tUhFoYErRrtBlm0Zy76WeCKMAmw05
0vBHySXYpuDf3DeILRP1tI5YJ2QVje5ueud2wfz3eNEm/AZoFjyKjIDznTF3K4gQ
PICTpJJ4L6RUGRYU4URxRHJe1XlElPqik78NSVfPiS4U9a6MfJUvY1T4EoIZHBMw
pA9z42pIksVVrSemruOPQ4cojD2HrRzRvhRQhYLHrTquhQLc8AdbkpXYwxHOQwZl
uDPlav/fL3goLorHldWHlbHSAc7t6YXYodd/EWvFj3Ill0AuGF5pI+plxP/OGjWs
2NwZ8qvtmBihIyzk4nEIJ+NlC0JbPJPeisiuf++Y0OMvqKDJsUXZEbAOOP8tAbdY
tJ21oCWWZ/lxvFntXGHCL58HyJLDx3+x+l1HFMbit7+xB89ZL98LfHVGwFIqYe7L
6Vj7CbjF+k4WynBBYFBMSrL9HvbGi7Qhla2NmdbTUhrxfQt3ouY7pQjMg432BUD4
GWr26K0vXdS5soOiFxflA4TzdBGoRVYl+cvPoa6Fsm67eDvArgCTlHA6pUn2VfN2
ub0aU0BG0IddGoQgIzE2oTHTSyux1/IkqnDmzuG+f4hxOm9NLRG8UNngjkz8atgN
M/ARp1jVcAMnROG8lPJRvV7528IX7wWm51+cmhDECOYsaixR3Uj5bk3PuUSW09yL
FkRAyyItahU1STtyzk0K7pf9ZRNKLFm7CRnxSCN/URo0cpuUt6ymbZkBx0CY1id+
B45V5+zDvwZ2PfDpJMm0lKej64RnueYDI1mqw4jH9E1M7aaT2aT74XmMlSixi9xP
sPa5K64j5KNYDNvd6uUoD/lME5yCq1xGoq0JbzTXUny5o+yonK5RL6LNK0FpqzGk
Orxp2+eXdTGRjsNtkj1L8HbQPInvp87AidUO/desGAgGHD+qUzWgFVjZ8pkh8zjH
34dhQs7l/HmD8UNWgZPjwWbkBPrAOsb/l9VBgq11yCCiqcxqtAG9X1wb3DEzNwQ5
YQqjYeZYpbYcMioYMjVTWXxxTOxdZsYAV/famY576bOnYY+HMrN8eDzrWDRFFVnM
enj1/OluTOEOyIpmQFzNgRamM+aewFKU/PEYSIJN2dwINhAmqV1ZS2fSxra4oFZC
IlmAH+eUV04h1fbRRnNJIgxF6lNsy2PrNxDr5qtz/VRyIskM0PZSGyp3apXouGkF
pFtdQCe3s+tZm0N5oU/KiXm6uv2o69FvNrrJaq6QudOVlYp+by+e1+MVq6x6AtV5
zqEChpdmjK42Ur//tQK5HtAtJJ3W/oriMqTIGotIlrTs6+3pa2FwdE0RPVgkrNDX
3+MsRCrpz4+uDC7GMvwnON2ALEwAK8PBoKWg61BLCwMJvAJex+W3pD28Qf9eKglX
+CKKGEIeoTeijeetuKrUzUFuNOsK4VHQwpXFtGwyuHbcRaEA96mTEdZ5nkcL1HuN
jIed0LGl6NQOzZ2J+A4GqHdtQlLu2rLSS7fF1mjXVE5fPbyie75mC0ocsYDhYQMB
uoB9il5ZlwlHHYZYAuGVbbuGOOgO6PxQe9e0G+7x7OlxiJDvfYpHrsvYNSV52O42
rJ4hd/KrVWo3WRxBA6OImBT7l6sft/f68siifafv6IpSlv/UxEq3OPtYUZyTXgxv
6KX0FYH2kWhizVQgEtOBFns5CnrjT3ev1HY8TToHgLeqIIQPHdyIDp2aFPtvG34r
YQ+S1UJrEOLPQutlhFZFUV5dfepgF2facdUxwV8PWi4TLtNYpPCTEpzfkhxVCnrD
Qw2jHhZsKeNWU1OqCsGpXU47EeBySqVjehJ/xkHZRH/Vk0hMcwSS9NMhPc1Ig5+1
b9FSDzkfEGWP/f+hpbejNrbkPLtFwqaAgXksnaRMS1Gcy1WwsPyUZNyE17dxPYOG
QNellG8y+BZb0l3uW5+ZFzsXWWCenruWlRY/I7BwUCD+ohmNU7fuzOWIc9RHH5Lf
HUEOF7EOeeYRp2EQOV9zU1/MRQVCgQwiH7O8RSHJMjqBJPpUV9cU2fOZvPF0rk9e
G1xA2b/qLz37Zu1a1SIcCv7zdtn2OXHgsjz9g3YRObXHpFGZo4UBy0oPf3NVSUZO
3EhsmBWQhQSbcCTtO2kZuWjfk1j8AEYZqgWK9rlQf4avbzGVZ7sGh4N/lZ1g84a1
ZzWw3ZpAl3Cry3vYN0LpYeOvkbAbH+jOBLZdM5lYtEroJFMMIw+Ap/SZZMlxheju
+thhJNRYyiEOrfzaNTzTfdd3TJYpTt3KfpZJOdm2g9L6L/qrryqX7K/JZ/z/yBCz
hzyUWcA4Bqnt5qjlz80b9j7GITH8iFmRNspLNRyW3RzwOTeU+2icrpbB5tHIaKt2
VhwMdrWeE7s8szKHyf6dSEU8ZuYPY2CSsrx2ybKQFiGpkt4nbpJp5q6OLF4I3a/M
EgJN2+zgRsJrK01btMBQlJmRykxBNaefxhtNMDkzfbUgBGz12VOB78a0/UnYUHFp
34EAiFdeS0xV89P2zC2izmSwhRkPjfWe8hD4Zz9bExzPAqj7cEyQ79fVO2CsZzoz
6W/84xv6pNDsznCD57Ik9+6tfa+jt8fCv4kHZvJf/bC4PjrxaaTWs7+94Tu9pNao
BMZPqXJW3FCft8Vfte8pgzFMG7HVs6BGiSa4vL9p7G71U0MfYl8jFtR6c6ZNuwmG
YfwJddtFe924ymoH39R77FhUyr6df5IGuOJ3m+d2ADmCHknTctNobKysBFCxeoA7
240EYtc3uasvcpjluN151eORx1Xqrem4/aEZNLV/FjB9QCMFBmcF8nOChwRynzhK
LC1bks5c57BCKodxQogR7mP5R0fx7+4Z1qempwZxdkzUWfNWAPN8NYduY4Fr9PvE
npm3lylj1joFAvM4jw2ESIR886Crr4X/pwynAS6KOlM=
`pragma protect end_protected
