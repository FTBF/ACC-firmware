// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 03:56:19 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
d3som29cclRjaCj6XsNX3T0FQN9ejh1DoEF+lCsbiv2nJ9ef8xrY3VAcmQz5uYPd
2cOIG4nhDARCnSj4CG6FD3FjP2TPfXxkLCZ1b48gxced6ii1kywaRta0s088mcQ7
7j3njRD59t6BSJ0vFJD6SjyYR10VF7atxOIjRQfssjE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28160)
OIuT0WNdLdis6OVIefEBwEjXGW7ZFsx5ymQy+a4KMZqE8Teb3WoIF8uQYN19TnJh
5lv9cNUWvmZKv6GdA3x0f9cMfVttTL2zwLhRd8lsw5xI25OYssE/oJzPK2j35yfo
We4eoT7JspuGIdk4R9Oi3VsccblA8GGKHHpoupAg4df+N0qvQhsc2yfdmtk4XO6x
bzysTZocIFn7nWI8dj3cOan/diYwa0bTTIZEgxgEf1KdoiSYTqP3WbKArb695Yon
apVuRKYIPCo395fuafYlMT0by2WYPfyoXO8oUECbX5vJTopAkROmDZCa+0njSWZ6
9564EkoB75gJSeS9E5WWB1hkXvOheFBUtsqOndOHnJogJNpas9Igx8PDHO8kDRQ0
J3E1dlLWKJ0XYShzShzgysZ41sgqCzdWFEiXCaje2KBcITG15prdloXZkeX8q5By
aXGMJmQ8U7co+jrDozsoJ4cKCwO9GL3nJpJCxfUTC0nrJrjFi5Y2bUFoqIYVDiFQ
huteZZszKZoWCkE4nK9Bun+GtuVJP24Q2E2v9ESetWgK0Cm/x9n5rdK8q60AHKhJ
Ztu9yvrG+kl56obZvGn0Wja9P52pXnpPje9StIul/sVNom7YbcJ5FF/ualZlskoq
7JLO7X2BbkoRkxsxUcLxQj7cC7A+1CFFvpAzKfvAaleYrJDWkBE4lIe5K/cdJLx0
hiY5fifs+vh2Mqy1ZopCvq2VtOe8VlL+FuhHZpkzFbAugs2zp5Ez3hSQ8mkrQGze
r+tivmIbPrm5h2WiDCLIEwDM+qWK8QatoeQCsS8/vgWftlICpbBicOqOaTxilbUh
vXOU4p2eKtTe8PgPIv6OQWavzMdztMVXBZhFynrGY1JOXIWD7Wrv3Sit9TwUS7sH
n+zLm8rY0lQbln9nYUa+CdQJrdG6oxOBlz7H2OD1UdR5CCaWkL4nU2zFN3FWUni/
zivmMLKR/YPEO2IvRhb6SwzRuY77R9sLzwq0JxwhNmnrfa8dowDAxvVNqbxIcHFC
M7lpR/j9HWcYdLnvFVFnVNF5NPNCC7g9enOTHmk6X4zjBEBrfftZ49YKOYQfJm5a
IOP0j1gTwZMsCMDrfqw7fV4UyL0wyob666Sg/vTP8MoPxEQeaskfiap6OekNodpU
PBjZaY3uhcywWctJKif1bmiIkyALVXYutA/Ssrqk1hrkB1v5XwoqYOPsZNNFwaiA
QmvEfbrNa6KX7Tx/mPR2a0Knujg2gc+8i7ZorbT/UIigRRa0jYGEraDgicwQ0vzw
w2zdum+B7lcJz5tF9Y/ushKvSLXSIWaJWx2fwpZwmbWCeoj7DBDN76ylx7PSpLRZ
u9zDO7LZalZA8UDVK+1SYojgk5MoX9dvwgLiE14f+J2gu9Ff/hzJBYkdniZ/wMWy
Hslt8/dqyuKj/CKtAGYwN9bBzjyNeD7MXC9KXNf2BRwXmWtV5uGUTKmErxGBjIoz
OSdm5WFSrjL9QZjRlmVSnjeHUq/gqMenknF8ouBTUThgVFtxcCeH3iP8AmM2BwhH
HhkmuMqdgwhWBrT1gXVWusiP91oznB/B2JLwxmavDo8FbHw+t1dITtQdyvnk3CUv
KzKEE2jm8o9svrhGOhOYwUP1ciX8+9VawY9b6UFNEFXofJ56/1Vil3Rq4quQxn8L
NE0falGZZLcDqgQo3L+C7zggjQRUkmE8Y6kaMATQ8kEsvaTkgRwdnhHQnxHcp7fi
jDKSlVdO2rDii1dubVf7jOtzaOX1/wbVSgOeeg4d2Hcn4K+0Pn3+Cs5JhiakKS8J
NvyjRPmxuly6As2FF7ay1442wY/qWSnDSdddaGW9ZXNzHsAs0fZjO8rYU3ssW9sz
dXo6/3GtKkwbGlGN3ECKCu8rPMgFwljRFUp5W47SfdPrwH4hf4liXjkhwC8Etjn0
rZHntLLhNbM2XPnfJwsl9RL3thtRYjijNpesAa+EKvd28BHKvFGNPycDsrnBY3KK
oPowJ91SEV/n0gP2rCGJEbx//fuKNQjlqRg3s+RjXP9+FOvxTnIBwSqF3uRCmywD
e7gQj7uY5WpCxyYk5pqDDV81dqwknal6xwM5RWgV3EalTD/BuMHjNQfWmhML7l5w
OL9NecuVb6HK6JpGXDlw6X6QD5j18subXdX9mh0CQ0KmqvjcC4lWfqDYZHJwimwM
EA9+aiXM5f0AoOdKKHR+feQRvmHXqbBadnmayD2EPdUh5v8oR8CW2mSmkhhDh+vR
JEEVZ5K7BybBbOh8Sur78iJ+Kl+NGEE3OH3ximd+NH8kDn0gqiqqwHftqtZs1MJ8
L8X1COCy8i824wxgyqIVB6yRBoyt05jAedjH1/YCXUZoJ5ickT05iWxVAczLlnzK
93+Ui7605z1BqmJi1bHCbYxLL08bvHTWYIg8pATxD/8WO8gMmiwrtDOkrI7CXaeZ
KHvqWOAS4O1wfCM6J9vLRFx1SS37ICfDvRAhCsfobojkAKw6AbHsSHFmk8u1Tr9S
JHbNbAhVVPbGySjdRgU4iv5zGfwJD8+Fqmp2uN9fnguNdrNcZFzs3AbhtisP5cyw
xhQaQNdj8yrSMNG9eosElQnR4YuB+SR85NoZ8tm45BO14i2yRHrYsw7jZAmlqXng
fhJUlQvYdtHPetxc3rYiMI5xSEslGKOyN6v4Sezl4/08EpsaAW/EL+S9h8IpeMxm
w9Xaq1kWxwGLyIHU8LofwPf86hA7b9s+u/Z16CX1I0Kro2QDhGZvbswmyoEroSO/
QoTF/ojqqAn5LbeFRaG0md3rbFyTauCfC9IfvuOUu32LBe1klHN+p1UCSJSzhZS+
PDNYR7Yj45ZNUjKPbZtKq5wYibPN9irdN4R+ashZg1sKK8YMqgqRgMj82gmb8JDW
sFCYwaGXaohR09F5jvnCVLjjrM7O0V8/I0/jLcNFsfVQePakbfV5xCgtFHFwJkpe
o5arBYLo4IUaPMvYTrxUahTiRYMDjn4z5Pp6eePS7TNvTPfueBei0i21tbQd49nr
cxfFe6VU/066dWookFiB5NofxoUzULkoMwppck00yaBpXRD+ubQhWoX7R74a+BOa
6O4HsPmWSxoZmOWsZ5czlQebz7MYLd7/Zc2Nc7ttJ5WJcmSdEBbflcQViwPH7mRA
z3WZAnYTNBsS+ocXdjDw6uxJB+krdWdQlZdodyebdrqF6UDCiLDzyItp4EPw4Cii
ubf9/PmZuoXiV/BFab3gDUvm/INy0SnJn/DSQufm6WcSB8vgyR+/5epT+OYJymYR
8RTtIM31ZrGyIjD9uG7VkM6o1Oo5oAF+9gPZziIqc30+98QOrHM62DjdHRApWyJh
BWp8OwNoLN2xKhEXHExf+YXf1T6+/3bBlgSb539QmTa8dKkzXlabjUJr9pt0lNPZ
QzbDHBzR+QhXb6uJbbAXlKgDuNFpgvF39Uw7f/vR4c3Ge3ZkcTyS9MrKzmksfYem
S/xmGDVlpcQr3mP3ds6v0v6N+C4TjjpHSxkjC6yi8ajXIYqsrlQqs4EtH6jxxrSW
8w5UdDpRhrDTXiWMJIumB1vraNhnVyVLeSMxnTHfXZDpg+RznQn1xW/qtjLf2uQM
Igy7EQy7nDqVq8f5Ft+QH8ydc9cHwDz2gSA0eAhO50oDxzRvx4CkNMSLOySw6ltq
Mec+3s3TRIAmhmYXx6szjEAinpWKwnouUnnrsWkkT+H1aNx/qh0k5SNPHvFeUolt
meY25j5tTD7XGcPMn27C4vjgfSu4LAtuE6ZcZjfWybOLAKLakkzBxNeSfX0pE45o
PMozJTfOZuUW85pexh+1/Ic+ygBMe6FVBZu1hdKsGUNI0JVkB+5PUAdfW+OZ3gms
s0k8TXnoXsib7YxEYPT0+Jmh3N7APgqwIsUlc1baYd4DZ+HFPrOjIaglhcAMaBSJ
QtflmqjTerh2afoW0wjM24KXNkiqmp19gwcdJd6a6vgqa8oshb/7/OI+s0x0E97r
S0w5r9w6mKsNokIFZnA1ghlZ1xxoYeH4ACyEMbRq45Ql3mnwZ/+KvMPS1ajBBgKo
Y2/ZziYqTd7S6iYP6TrjMFW0xhhMMQb3SroQGFYcKcTAG0OO6f9ngOCdjf+AACyJ
oqNDjtLppUhstU0ETZu2ZuC4bl2t27ZasAybvLPI2FVVAUo+3lNErS44fk3F0NWg
ieR7RhaspyAjdPmpX8CE+KeoEnYMvBI7m2A/NNRruUDesW784OVQbWA+hwe2NC7U
t2VhyGo/jo3ffGC5qu2owfw7QUCSRBti9mcZsay3sP0dIRo2br7RG4JTU53Otcsv
qNvrbAtMuESRygZl820slsREq8WlOt3H1ehqDFn3XA8spRFDLh9IJ3Ue/j/xHdVI
o0OaIYENHuG+eRAnPduJqGi4ZyUuhgbrdCkOugTJ09qzqJrsLoGHIVsrDHSKYn1X
dLC6HoM4r2Bq+wIBvujqMMm8Jb2NheZsDg31pmrjloVwDiRmRfe+A7PE8e/q5a1a
yJy3BJtuiddMB2yHYYp9b4qCcoWx/eKMTC4j/VNz7va/ulA8phJBdxewrD+prjCJ
QXWxFQnL+WGMbrCbSYZLhZL5FdzCfAcDlSPwdAfuprYTQy0TxQYdU6NrzWx9VlBn
cS2SkgCh0hZ44Ec0bw4d07eiBasE8z+5m1Hl5k6j/DEtakfW73ajL4IxcPQNn/fv
eqkhN6z5/qH7r/I0mw6TugL7kAoittCK8E7vmhFwXc6FWK0LBTJuc7RQ+4meaRvA
yaENuRMNPtTkGHb2bPYDQ3+aTLd2j2sMLHtiPB+aPl7WN8fUiaQ7kFCr+bGDC1rv
i9xrCWb7iFt3l9aoo8c3uVBdL+JwWPYm1KLlvbL/Gy3WxV85BHF74EYtLn1pgK4D
yquSdiipq6dtO2+kFLZUrTirXN/P6jXaTYfuXP+YVGBLGIwqMHD1ECdT6HTMdqMy
2JfTVymgS6UpIyI4b6GN/sso7lwt8L2bqqq9deD6poOvVvpp4CGZXhHoP354Zjzw
PK8CbaNOGw9lTNyoWba1aLsIrvtKQUBTo1EqNvNvkYaslg5pn7DzWf8x2R3ZO12b
n2hr2DgsR4DvsPZ4FNE9VWCEPzS/klvOo7eQpAI7U++HxBf2meT7N2k6ox7SC94U
kJ9K2wKeNRw1TECew0xTNDRG3V8Kv7r8PVpwj3aLU0nkY+dPjA+UIiJa9rRazSL4
ZVKsIuJPoVQXexipwqiC88p9v6PVjoPN1mKAYo1kEvWODpHxwj9vsqmIfCUjETcZ
sU7E4KAwV6M2fvtynugFpwerMeOSgS1GPyigRUj126gXGaeymenqrr6UGBTWHwtM
sV9WHWDXIcF+s15HDw7vx40+iAWO0Qc6HIeYKDDrifNwUH9jVtuzmjWfLocMCbXG
hvF8LTjRo7lrInA1Y50EhFD+pnqmokcrxjVMyzccfx/y822+6OZmxktrOmqsT8Y5
i0bHQHSWOszgH1RhpWZmi6sybbVOzgII/F2i56Rb3fTmm1wvlcSUB7L8FfB2XH4N
I9DUpW4YhPnCiSy9wJX2sX/Ozii5XETIFkXr55aTcMgW54I4wTypDgiFEF/XLsrF
ZDB2oZh6cEICRdHizun3U294xEAkmVLPF9AMO1qgBb17w1LIubcra3dL3k2qIpsy
0WL9TVbZcj+fHh71sjEybz1e0ui/TmkPXRVMKLSQUvD/6a+bqO6DQJ33TcsAri1d
mAGHqyNzPu3mP2Dr4naHZ78AMk7p36YKjoQKXrq+PB+N12Q/2fuXytuN+cUx4X3+
I2T5ohBk1BL2ZPBYoJk/leohvsQihRKgiS3r2xtr5CEWARv5NZ1rC/EWnsQw355O
OHjvtpaBqTFUELYOHmuLWxmyOxeqZ4T33t/JcJzRhM7H9XH6NWschnoffS/+HfiV
609TItT6KU/rXijngA3rNHehAjzvEudAcIgL+I6RVnje9FgTzJHvb9K1BQmCqWAW
Ta4Zs1Y0tK3R4U5nYNdmdGd146Q7APJJ856hAJHDfS39i59bBpF5OTR6+arHiy69
wZT+cteZQCFlok1opMIKpl+cK1SYRF5klb3IiSXFfmuzuAsqb5/ldnjenCLOh1Zl
YCYZ/Zhd4E0Nwb6AI4tedQILd+XZhQZ1prQEQATGmRZ3VLq1QaBLGO43MUaw0Jm/
CbKlofApnbT2B3nvJ+z2tFrIqRN7Ju/v7MKLv9eccI5/HcOerj6uLluRsV2SCnv5
/ProXcM55y2A7WbAjP9sBMKBTtnjt/jwnsQ8TJxWEBtiTZcCmk8Nh+A4/6DSN7bu
IYFO5iSB5sklM5QwTS3bDqbdyDM1b59+87RSMsCBZc+gDlqFJqW7py+ORr/1vf8B
tey1KQRZxMvpiWq64VDHSFOQEfEKYxQYnBY2D07iAnyg6Ls5FFTxsqeU83ekES3E
suuU0qIm4xPrRftG2+xLjkb0c0rvgckmPB8r2dExeht0VnfzawHi4XsB1bpr5yDW
Q6taph4NukAlyMFQf3/FYF4QTtDhq+WKhqtOpbnwBy8x2p7SzacTv7WwgWVjLzb5
81Wjk18Eij3nSzjURozuLKHJ9LrBtjvbQ2abh9oZvs/XwJ9lE6e3psz2NReT2M4x
ad4IM9Jw7clgmubV2n7UtSj+hUdkYiLnjVXdEJdKms9HZJuZx28LZf3AZgqF2qJn
HTPvBwkXTxE6DF2aQpqM/YL4L4SCJKyn73O4Z0T+uNZIIXyuiX+AcU4jn8xdEitG
DgTGQTAlUZx/FW2ZsWT0PlkFnDNJERhKtm1VnQpNZ7blA+CH9fWgIL20QTzXZ0re
8NoNgQ7dR1x6r3ljjDV6eZa5R04FtwNYfbcedys0ZmDKinCGPL/WSVhOV0zP8We1
cRS8Q/VYE1P2kXSxr11VJ7vQgGcV1sEyE1edA7WGXnciM6Igdp/szWd+sUFOMgke
4xsmyd9I0DBciJunaU89VxxWxyMIGvgh7xePhIY1oTogHRv4pWE/RJ14DC1T3kwj
I75eSHDo/cgRXEOh7O2kSol1tLL8sDGtdTZ4p0THSJC3SN4n2ZozMPXj3jZLd1Ng
6SqNSffdcwUL+eqXwjhYLvLlEBfQNkvFUJs8Wv9+xCasWd9ZR3KfH2RT8sMKNYWs
INzt7nZN6Br7nfeeqr/jc6nxbPHX8kh+KcP95KJC8AlP992R1GnH0sWARypFMZVH
N5AI2tkiSzggi4i2CaAAvnEX5aFtol3cROXNhp5oCBiL1WefeT1q0Q485BlalBc2
+iWmMj6v44aE6vp1Akkz3WGfp/KJfP1tNdkHxllfjiRexZAH4wH3n1Xln4WV+jAX
vkFm5z382ujcFg0vsl30IGgbZtodRIg1b6plLiKbJCMsxYaiV782P/bTYrFc8M5r
EGtYFat9cP6Rg3vkdcBqO8vxve6cWdcbkm/tFx2gFiYRTc1W2lWVWqqb2IEb/JRc
lMp9L/tW4HVmuUJZt1nsVm8ghsMN4hi3u8oK1U/FZv042L7Pl7cnDYCd7xb4+PuT
zmpDF0Qq9EuSFzewIXnePSVC6lRP4TxUGZy5dwWHjngczZzim/E+A72ILox4f4f8
HmkbL6Wu8SPpmHTtDTd/6lZDxRqW3Drt3gUxjOAAPz7xMWfw2miAk1x/c7oltYYU
8HsOLrjHpxt1hNKo/ujuTVTiNmXbYOk4g6CVnbEUTPbp5JrSLma1aVPgYzg/GtnI
I5TaXNJP0afFIEITKFYI/jloUOO971/lzhVTryml7ecE0WPwbGadKOfaH8az69nn
oOVl6wo1gJDL2jZbe3e+xR+aiS/ad3kl3euk/lywmMcOB96hA+vUfqhRcfpSI/uB
TEXX/dUcva4TdnwhYfHt67y3/7AFToTiWdp4Tv2V9cMkdUkTQVCsz2vwc1LVb5w9
PK+24GF/nSoRUeEUXDIjnY4+0O84hbkHQmTBt4dOxYfo1VDfCtpxZnG2if7f9/zu
cL/KIjlMMn486m43pDMnfrOZQQQCuJZZs8561OnifrhgLUTT/J9ugCG6TQbHY8Cd
mWJwMKhj1YmpYw98RSxtANBtZoTZqcJqKHntI/NQikHKqdu0QjKPkC392C51k0Do
FWc4utLkHwI2FcmsDres9ahVSTjQI56k9JU56cKbpGZaefHNi27rz59zW5KDyjVz
+GZZ3CvUVf1f55T+4RRtypZ3QOQ+JYitdANjA/rdp5FJeg2Us+tNIcCU0aAJXWNR
PtINYMGrrmYTGp4a3BXogbbrBYvcz5DwA49i4o0iwP+IMDIkX9Q0AitIcy/lScxs
l29MwWFyPyYAM4IX/NLb5ZsBRx6MgMvWqYpQvHMVQi9o818aDCzkS/zIEi88p3yo
YCx/BkV1UbUvt3buYj3CIbzPMye8fbcdjgIWTXM9wsiZ85C5ND6dvQGrTLHJSLTg
HPVfCqG3/NR1k/65glloGQdiAEJwebPhVGDLaCnZmy4LafcdcGDOzZM23I4Gnk3M
bwvLaBAXfONVfd6rDCgK6MsqPh9xf6vM58BxXQ01bc/ns9Vrg0hna4PB5Ch2o8tc
Z/Pavq4YJ4jSj25uJacY7q/4EzItjyc8lDOO22mKvsFdA/fK0BLYIiF0hw4f2Th/
XdmS0c/72gdvPy8ctOHb/nwE2CtVR0tAWSppDRCnvEb3U1Pwc3h27MPtcTEhwBNB
UOnWczqUVky4wj1XYkmthvN1DhaAlY/YagB/2ATdGDtdZbAf6ixOAQkKSfQALgvn
Ubmafd7y/4mT2vZKCN51ctdErUIvo8g334iK0Vsgx3r0oPPUftS0sCLQtd8wdCe9
xLlQIcEqej6KSf1FZU3M9vZQhfy+h+o9cbvkWosyIO8v5f85q8DWA58xfAszc0mY
v0ipObv20YyHgPnjP9pUiyRI5kBc5/I1lXY8M1vo8r2opYyJCasapW33EG+/0+kE
djxx4cOn3dyeDsKqLP5m25v68X8DXtBb2lOWWuwqkkCeM5s/0JjbFW921JsR4/Oq
Tl14SaIX2xGBhXCZnWE8r72V5pb+XoDoggT1X9XVMbL5Cyy4+nYIqOM47wXjcN7y
7gTUSBg+hGxq5FRY65Bnnc6orwY6TNeoh9c1MATWkzdzjLqZD517ikgrm8ZujOef
LoFlBJPWs31PO/ZbEVr9jMCimH/Fj3sEoShq2zr64aKDCai7Y7ThIvyXbmjyM/9E
r3k77YYxInHC97kNYij+bU5DXneszNlIxkV9pWf7ayad6+5/hM/WEw9UHOvobZnP
jCjPMgCc5gyJ8O+qwXuZheLeuf7Fi2XdNz74wtapWlktQl7xp4spwy27g+26olsj
i5WMGWXHLbTYQxcPe3Uhvux1y2slfCneGXNNlMJ/zbBhOjhIbTshutyG4IP0g3Ab
BAFocIcjocVLYU0x2u7Jagq6jdDUVXprJLQSyA2K0J3ODYlr0WbokO4BxKTHngg3
tHFFsm07G2jkX368BjuUh8mfdYH9fYY7zHWZpBQfs/9o70BRZz3Y6j52fh58GDpk
Sbayxsv3TP0cVqYwhXWX9z1loN25ujHPwKPpYWVgJ/k9WQwctk5e60SiSqq0hFLC
PUiI2Hsft879Dcm5Eib9jznIIorzJ6EjsgjF3whplMuCicL27b4z4pbbpldaqKxu
UYhntaKkhxprst40Am6wnHCx8Bqgyx07BMhLD+pVLcUuyPLFfTD76DM9rNnB2tRQ
xKiK7wK0a5eKfu5AseA+umBChFAmxPMGf1IjS/DyLuzgjbIhredqIQZBKPZe2S2Q
F2PJ2J5sfIvKXNHTfCBB9AA4p82CTJV06Mx3J6ZLpQ5Pxa6lG3b41uHLln8qprhu
cArZMru/2/VIuh1+PE9M/Uv+qaaQxbYjx8OM0yeW+j1uGBHG9/EP6e0ynftHZwhm
Txv+vfodJ091QSYl2tgQ7lpE36YX/lh3nNuNb6DZWZlNBUYrwZ3MJvLZyp0PBx09
Re37XTPX0KVcP7fWGZvISEaoOYBWpl2GuhbamlDT/BaoEm9B0KRDHxGI7RjTggFp
Jf2tYbvQNRO9el3tnTzwGcqCzI9WnIBae5LIQNuAYXsfnGvW5Cp0OWlN3lRSkemN
RbzDRwaE3kfNeqDqAMtzA3qihrtnr756/Str4+zS7LhZnhfkrNk1ZzcYOmjWUyFo
e/yizlRuj6s/EJ7fttL8piMyARQCyaIuOMIvGF5VormW4axLWh05GxrJYi88D2KQ
qG2IKh2d1aB6vL8uH1PG1POgkg+iqHnxoviGZtpfSTuTaJSMzyMtx5eA9FUcRS7A
B3/C+mJM4GJUlUTvVoblarRquYHbjyzDxLmDqLQnzfAezGHu5CSjfo7lpNprISzc
XYsJKqqno+NUX+jpP0TqvL02U1cBiR1efzmfsXG9ZA7M16McSq0xDxc7hJiTOJee
AzE4XUCEjaOZsm1UY5v1tMseIEEHBbb3NpNm2+V45bfI3bD11cmcbwtDsj/8ONIP
+GLK+5ygMlCeIG7w3a+RtqChVNwh3CmSgwUOXHITHCjAgiJjV0z7QaHVE9M8PvT+
GNDUAPeSJEoIHe5Tep+BC/sFzuU585S1AhgkQ7t4T1qrPCShPH2tWpKoQbS7vAfR
Qw2GTsqWf8eLqL5R4TXa/7ft271mTulY+bZeZR05tpza8BABQ0cSO4L3xZyYKcog
4r9UDVzxExEP1Mw4B4opma9yKAbC6LBV6v3LahqMT7wkINovebwdHuzGX+zuz3K5
2oMPqQJUHC4qbdx3XP9UbYYqpiK/KthYdZiyL5pn65OeuQ32HeE85tnh9BNjiOxJ
t7sUaGbf2mZXWyOc8pKVfhAdfDbXp22XTVo+G8gOj7vYw1nQ++73Do0zXiWGivzc
0cPZ4ONUZpsp+DUldiJRZJrNprdIu1b9N5aZh9E2b9rNXlMfUIr8j2I7IeMvn1yN
tGY66OoSnRmCgt0GY3guv8u04scJrlddKqVH+QwHbWbEk+Tweep5FfxJCvk6dNmc
6q6MIgQCvyX/x5m/kdA67VI5Rzzam1253PBmqr/8qIneqX8DR73h7NzoN+WK2Ixh
z0qA9+iy9p0/C2F4FUr4jyqORxTp8QgG0Gm8dM87gJdVtZ2/Vw9MmfvcasNbZR/0
cs9lQeGgMQhdYbZG6eIUYBywFLJggUqfeesreHka2XzirQmlEeI4mg33v3FhVl0+
ZzOCtbAtaZIS/1XjzERmKA2uNqxYy3ChdPD+pTnVCvkqGeXCMFLfUBxZESoFTg1I
sF7ukvNRQ7K+W28YM7kZ6XKFaphZ0iZGN77sNHdtbGNBPvonzHVrCxcwgtCjo++Y
KcEsfO7r++G2mwE9Nw+cGKIZJfHknJQG/bHTDKqii624HPn0xSgJQWm2W+ScEn6u
lqRA8URUf8n2OHHm+wqr0Ge04ALfk3PQT232IiSk7MkeFJ4oEKQ2QVFhtIdG654y
kQgzq3Necj8tKbU0oFNOSm4JnYYJOUDXydl2kZa58zbSdQ2h1mHiay6zjONAH9iY
tEFw2dDmzh9OZvyWqELmOPPeBot92a08vXVDlZmDboxd1Q9eFASD+Aa1lmAtpDHW
UqNeAiGldPaxG4beuqkiSNog+39GRJsn9QNIrdazaWdrzoFMTRIl6yQdL/ZTHiJH
jrfUOE9zABk85qCOZgFugBjIS5+OyE8RRRhCs6jL94UD7PhxrUof+2sDqpq5avbo
dJAUubk4FEoJRrpW2TyPY8dWIHqCPAhxJfHO6Lt/vWWmdzJoktBmwzpRchAZOjTQ
XQyt8yywtOyXcLnhx7kj6KwUZkliAHrohu0dQRNmpqCBB9PIIr+Voc5bfDz279/i
m19p1iz6J1OqvImZlFJoKQitryiWiIh5NXfywaPwKi2o7QYRyS0lCe2JMpgdVnFr
dNEv210glt340BPvAFiW0EWA2VOA0PV5ZUFTE+23NlDt17PmKZT9eIeAlIlh2zfq
AbFGoujOkZ2EGHDij2KRUM8W8mXD4+fov+5+7jS5N/0aDvonwnR4oeoeS9iRuFnH
C4pC6Tmq6kfSVVPV81ieYXotym6mNORHMM1UvBb4t5hUetZf5gGPgHYH522bQ2cS
S/xfGDorUZ/3w/Wn+CA3GxZ7fuIGuNlrp/i1Z3Ik/HzHdq+HOdd8byRNNmDvUWKb
t6wuUtb0ZLGEVeAu3JvYcRE9aQMJ+37wbaHsFHL9b/LI2B0nH8OSAjXA/snvC5uG
LmH+2YO/2UxzrBofCjzidOgKho+BuAMZiENUfDzOqiW3tOk9dfigpHoS3PfZvtLe
dlx9cvQS7Gu6PMcz6GBquLariCxcroiXzOA1bNNekJVZwEcpFSQj5FxnyK9dVmMu
edkpUe0B7B4GjJdF9gAVAnFIf4bBl14OY2vhEfEo6JOSFd7zcl5kNNXuWRwusxXx
dMAJ0cCag8+/0wdVEEnxkwaZ5nitHpmXfi+B0MePTzi4D/l+CPDD8YZ9NxH+WVqD
5sK+NfF//Yub5rV7j0uyLUys960YBr1G8fU9sFOS7ACrRI2SryFZGURa+5Z9cBoK
/bEie+wnclZKvfjuxfXRyMEkCy6yc0yTlea8tq05llU6ItlHgUDvKDRVz80FXnen
n6nrpAQiOv396FmfCC67gD11OMNtapxnPHVHAIIae3jcar5JCQP6HdgxCdpD26A9
LlxmfHNcyu6Sxa/XhkUe0JPofug18O7VsWXmdf2/8MzcaaxMY5RBUADyqTBMr2np
lylfnEHpfQvkT7B/c+Y3uIclyQ/OaIPdhxEdAciKzDNSgeXsT3kAZzXWqS4wJv+I
6CRBIG5CWEQm/oux25e5TWZBcaqxQLK5GnEbdjHdvb9HMRTDUdEJivVjLu0Weaeh
h6hW11ADlRcJpwItUIGUODq9F3biiS3nGxz6NyrkJUH8mtU8plULpuEcIGnbKEPe
MZHy++aYpnsqC7BWYHTRaIyTEsz011rw5M3+pQD6j6OLwE5sxpKHxCkwXyjrQUb2
V6l5x3/KGDQOMv2i75+heThXgJMk/CrT1Ib4KylM2rQCI2+aICVoyArTntn/kaQA
KMiZwW9/zL2QLa8eHGpxhPdgFN6PzDF85fi1H4r/QRxtSaaSBG4+nx5HTwLP0zdV
+KhdN5b0JWcM7BfaMArnkhCQEB7hRt3zcZnM1EHpi2/jjG14wOKt0FSF+ll0MUZ0
1Al6RgRyv35VOEn1kd4mSbY4DbBWeNmpMhq8jyZVITbGZjSAZwF/oY4xPal8J7p1
O7UN/i6XW9k0fsv9spi/UYPtvM6k23lEESN94mOZ8bah7NEXzcevVOBy2y01fGK5
6UaoVT9QSyaTdRMW2n2MImcAKtyTEMgY1ol/ELJMRwgyo68Jd31cdZ8USjGi8Hic
k+0YZXGAhId93nQMCuyDvAi39Ayr+wd70eZjqDfwgb/hBCm97Zjqc5hzVvkRBL4X
aN7bDjR4eYqBO9g1MDUjWsW0EHMpfYcECH+DX6b0uoLL3XdcRzJfCGVdsHayeGfo
JKnYrrKU+4NQDWc2dCONAhhAyuley1GYGvB6IC844V5mO5+eDIAagVNYunnW6G1S
8zHVnDiLXE8Lb42SgXY9cYm4J3IBHaT1wklBvjGkZrxh+Or5NanjyqKO76r/jp3J
ATUcYODtyu9A9NSEkxzNyVRP5GZ679PXahoAXDF1SQowiiJ6w4aerBGHif30Tfv1
IQMHigxKNxiqacwmv+yjG2OI7YqgIv43wB5iO9Wkb1I8xfp2FSVgJngtl6ebAn8Z
ul8/D4VVgwv9qVas9fzlrUBEvdznYp3T9JZSik8sLM2t0DwFVEoiw4h6jNo8Zlvs
wFaTnYgNt1DHGLcFwjQ1CEGlazCUimV0gCGJ2+Rz72zD3FwqT8cBKN0UkgmHdLNn
sj/+GggWGclDyKPn8/N6zDQbc+FSO3qOtDDb26ObTJs4W5vYhdwVShX/Td4aybvr
2V0kNK6UpSiaydKJsHsmOs1Z371XecVqwhTZnjTnhCtQFrFzOi0IUZ/zXVigfomk
KF5yL30TmuuZYqpLvmmOrWq1ys1KL4gpK/Ka2OG9FNa993hMtBBboto9UEfIs0nh
FhXemB6DnpArPq5e6IGsz4/Gbj+wVA/kRyFoAjLgVv5yEkOMs2Q79U0IZF9+iXov
n7/REUewsQCNUSE3o9Al+JoSNAlHxHGzNfja56Y7gmXBH/cpz7YyqKuItG8NjaSE
Mz4qpn7g9JDHU7sxVUQEVbdxYnwn0k5yLXvN5gLiI4G6KoIMm8rTi1tt/GH+m4vB
e8BhDGx0gqf14eAilvYyx7UqSN2PkLGZ4EYeVg+8NvrYYxTwuatgQ+eNnJQJAGm/
Fa6w2Q3QIavmyFEGkwvqJuy1DopDYl0mFSMGbQIQbBq0frEF3Z6XXKlbn34it+i/
XGZtW6Uya1cni3Qd0YG59iaKZ1bvMMdiXL9bSkSY0M96wOOpRmYAYhCNd2RVs0+/
6Z/JoJhE5cey4fqNzSNtnX8SyOdogDIF4EAosyBLRYr7wI+sLclMSM4CkQsNu2Sl
MS5Ah/NI9RmyjSiFFvC123ophGbgDwlxBTCvBwqAjvhqcTWm80WxIELqqd6SRczA
aMagidJT3kecHHrIAhhu1yohp5DimpV2VvIOeoZUf6kB/Zm1pgqUXZ8PfKRQKc4A
XDlDXBluJv4usE3u6xjNUQ3GqbBSlWpDpSJHU7JHRxdGhGeXMj0UPo9sHwW/5ivN
DGjsKJGKYYBJ5zw72SDMOrfrSSgwHtNxjO2vOsmyPaoEs2cZfeP+B9tjRbbntvC4
bB9oIga1nYCIwo4p+NAgK1UomhHyGsPKiAkkTEL2pmIP/r3Ag5P1ZjUvhhkotaBc
wBB3KwywWbqqDCr4MXRjQbPIbx7ks3TFL4Dd88Ih7FsKQ0daWQuDMjd5/bikZLOT
m/2BJskWYvHh2UktAn2ZzTFEs6qoUTE7skd/GNcI29NmCYZEIZ+9zFWQsM33aolX
/7hyxkVu4I5hx7gh9r/jKQ4URawXcR+vhZtAcOMhe/tVJA84f8qaInR38lIQ3d6Z
xOHnPPzTFAyxtLu+szZf7IsQcsMtytPvpBS0x5xYXLhT3QVhb1HfiHWm8/rSAVba
mDvRd3QXjHUeKelHEx8MYCTxEuFgHbGQolL8USOyCP1Tm6TbpRNIhf6oI4YnPbeR
ae9uDRPdItA2kNG7VTCyADzCYBntz8ccm83XqVOm6Yv4YEFmpRaxp+lLPLTA8gyJ
RpcWXRxkWENhoHKGhPDLXGxderChiGxMcvixab0oUUu4ds02EtlKeS4jCF6loLMM
p26o/zxgkTH+HcAxG429lspESVyz1LuIDv7d+vGP8JH+Fhk+vaTrpvrcaqgt0M1b
BYrO4p+sECyASZCDQQKOYuphM0qNzHoVMS3+giu8yGS9y+NiuMVfLWK6KpVlejFv
GfHlwBDUBCXVvHwJVrCjZqBhEINjUYQGx+yhhcKjEBD2WfLmTJG8DhRLzBR0ygTZ
ZGpYz/pe+s9MC3dvlW7kGDaYnUgI2vvx3K1bLpHiN+LNs2sHhQboS+28z6204CSU
h1aCNlEFO9r/vm3l+1EhLSTvjH1taSwgvEM4fGk14h6ns13lyyx3TFuGzAKsMZ+2
U2eMxJemNonW1d6jFSmJN9OI6BVH+p+mSWk+ohtAwrVFKjL+n4cam69vd5jP105C
3s/a+wn64LOK9GZsIwiyquOgtbxu9XlE2u5yp2M3w5nZbwzP0aK6MbvK2Cbf59pi
jc+JI05V6/FlEGg27NC/Dks+5wMzM5o7XAkTZsGf8DaZV96i7NgkeEBeFSkr4TIC
ROvqtTxNxWYhx2RxwEuy0gCfbBYXbzZL3PGxI6CzrYOzCITRxZQgVy/ODaSqHQCs
8iUtsmOe7s+Nx0YM3Yg66lC5VRlAUgKzlve7OTwD1lSSbhDVD/I4cza0gEYMCW1L
JHYDMiudLKxGP+Je4RFZXkYcmgJzGLVv3Qr21fs6p/59/frokVHYUg09A9j9k8ts
zfSEa2xls5KWxdkWE1XSjvYU7u7Oqrb1zEmpvZUZLW84mWZ8kusUqlSYp4mFeVMm
67gZyM7x86gV9rfQEd+IqI25dpaHPntJJ+aqKwLazb1UUO6+UJ54C3HzLXREQ4mP
6l9yDjjNUFvGepQkk2T2K5M7zHp1CvRGocL4478zEHYAhLNa18/Lk5FKJdslB2S8
9qPihAdqF9kjS3TNwIN83iz6iBQtON6PszOfI4ZRNErAKfmKRhsI0yKtwUw/5qiO
9KQ/5coiCrKGR9w/eCrHgj6mzLnjyW4xFGdFY/fGyvLXupSC2tjEj7gF2bQqtS2Y
vfJHB5x2Qvbk+/x23vmg5yfbjxk92CMNpJFrjzh6sU5eZ7DGNG6C1pb8vrC7IJfW
qKNqWMJpEFdUn15e7xYgLIVp0ZWpB6SRsiRbhBN+Ahkxw/CYpAXD2Ff21hYZ2yP5
6rWZlLBIsxXXBdN0uey1nAxZCnFzgJTu7jaHWHfhWwf0biRWvRgO1psH7EJhtTnQ
fEiwimJnC2pB1pKXoDzbXIt5mYNoC8ne/+aT71y6B5lJToAP56vBA1LxZ9yjMuij
IS3P07189FJB59XFId2ErOxYMZP6KryJR3uHvp/XKaX3D1Fw2XI6fCCf2kTc14y7
gC0bMn/+3C314nPraO8E2UQ9sLqBPANZaeV3jHIX1ZioajTMGNY3CeXBKVQ9NikK
CEoatWO04sUG8YcOH3VGztOhdEZtuQmQXZasC+h7Q3Pw0UYbEnxxvEUN+Hz/jbf3
CQUanttZa7NA6ozmmj7oSvQq7aMSS4bJsUOjmJUpZ7QPw4LJiW0YD/UDFOFf4f7E
OrWYfI5la+lJFftHVhKE9cU6JIZEQ2nMzBBQPf19e+hOyXNLjgznclBPQY8AGeRX
qyi9wOakq/2eU4kDSN1QOuLqW7MB0jrRKA1tlGlY5h/GNqJevYB5usdsuz4kXWLx
6/XxhqfHPlEkFp1a+3OMLTGAlUugJQFFKE8eeqBrhqghHBI5/3aGyPbJ1nRye8XX
iCZhgsAM/knAzxk9QwB2IcetBkiRFkXtLEfmZFPQ6Bb8P6exBPI3WN0LVts5wUiT
EWx2Zs60v1gV73Do+5xSgF4F5DplMDjeYaOhuiTQ17dUSGIZnWJB8Bn71DYx7f0/
mEvGNvTkCOA01oqhFg6Wc2CJP0dBuCtcIF+g78pNsIZ8Js/jC0BRhMGulcciP594
tb5Kv5SBT5iDm8FSpwS0ONCvpWKJ1AaGTu5MgCr5rW0V+ggM79mWhAJm3LFnfanE
hSmI7Ht/hYSFACbXddiYmfZZxsSVGMiamgCMYAJY9ZsFg7PTEKVfuX2xhtFTFaQQ
gE5Rcs6+C126SwoOhl7KgrehMpfOw1TFMw+toefoNgwz/KcCA9xZQ3nDGUogVp61
euPwqpGdZZ08+h5VZQWkzKSQGIP6oXXN10siXdq3nmAuPd5VrBHjuOSHLKizhYhC
lYVpv6nRbQMZFTfohtDi/KNKyXKjBh0M/p0I5gyqcf6pMj7BR+8UV2cjdOlc/sNW
LDT6n+9vyfJrPVdG20gI2G/igk6ykGB0FOIWGiVDbwrQDrSdzVeFZf6Wg2FLQDlM
Jz8ltZBlMShy1QlasMvRBc/+9KByoQNqN6h6Y8ZLXUH3qQtEI+67EKbHjimw69RR
B5TebinNOXqOxlzGFRD/dJygQjxQKFH3/2mUopuM8vcocH/eWvOdfSx6Hor9fE4k
wUIkclrAFei9Dllyv6qVi1BmhrwxsamfySYnl47AUBZCxlmrdyhlfk1iDgiAAFnm
4NdeUlzsV/GVfjrMw1/H2b5O3rJxQ2TwZPWIQ1j+5lEOqN7c1WaCh0NiGCTZ/OxK
LyjqrO0440DdRlIrIajGY5Umec2swOyyE/hMagQXhhLmUJSykjplW11LfdIPxsHd
F0Vgjpy+uRgF0VFoiJtQxvVQf619Nfmkz5K4zUpDnUG/rp+wNrMqlAMo7f825eM3
scOTuRmJhd22lDlHGH+3dVDvrLPTU+5fwFN1GAyQE0ldA/iZrMzPqr8GcTuj18SV
D6eLIEaoUba09AeuvZQXEa+mIZd1Xh08orZNbnVf7gwof8aviCgQqoDZIaYVBbaI
rKLTBe2MQ3V/HzF6gTbojMdm1drf19nEDUE8vN8Hn/X6Th4KGXVCA96oZdJjUiD+
lbd+7tV7lo47GAn9f0/X5TwqlwqVvJh6ocai486bf6loLw7hzEfC0H5UgAvUmoEO
hQfzG1eS8i2GI9GwLn4aaqLbgq4PDb8v7C4gnZPFnMkxNl2sAiUDn9RKM1utXfPW
ygrtgQ2dtsjBCfT73P6NBiM3QcCRWjjmz0j32alIDfyT++ATJMcYhfnvUEW6gqwx
X6mY1Bg3XR0FmfTf5oZR/vgv1/4Hpk2joRwiXprfKHaNJcG+/5fyZZ3CjQ/WyZrA
CaRHKEztyZRdsKngCsDB0zWe2K4XjDiaGZyANmIWBacITx5HWYMcGgepQaOkNu7q
ZtW4+18YYmROPPEWnQp+nv30tEH0Yx7cOjlIessFOhOGCc9EwscBPhzjf+9vREFu
bRKpVpAOj7Zy7U+Iwo3oAJ8c0pTrgsSsqxLKB68QvOAdLhfl7BueUZ8AAI0TB5c6
iGeCanbzEcLlDVxhYFpNGzcpMmO1gECDcqPulREK3Lj8wo0E+cAk7+wujUddqUwF
U0Tso07sE2273VR+tShPcHs5dA3iH4mizjj2lU6mj8jdSLaTorXp7/AEplJbePoh
INgJluVWeE6jKmYp8JGL/MlN9uddt+o1wGnrPo7VXkVrqRb75oVXZIHiRN0jn7WX
dRP4AoioU63cvrm/2NouLSOoyqIuittdNpvCZh8BPQ63p8LjVFR2y1hSx8/zb5xd
Bdg/w9S+E+sm16JeyBY7liUj4v/8wWGlvu0SRzjOge0JS8TJEvYJv1mRaRcNbvMP
in9k/5UW7kXJrKH4JMEwKPBGjOkm2/Ae2HhAoNiegdeZeaq4r6XxlovKVDN0TZg2
Lf5mrurudEa/1Bc0K3Bj4FG6rBQIw34qHUlqYL+AL2Q9XDB0VqLM/UO65fN7XYrg
5PNtsnwLr9TBoodIdjgOKIPe4ZQXwnJfmeO3oW7/hNshDwGpo6QqWLJa7zhDm3e9
UL25glgl/kMF5yzWmuuEmvBNcoAmNan5+hYG1sdv+E8/LqJ7yt46IrBU65INICFZ
TaTBLm8NufiKKqK1URVa2y98UAh3zOn8H0X3PYhapstSobEpOkcwU7UWGS4SywQf
Nx3hH++rjM32giz7OS/Hw1XzIV9gU2oAMzw8eDCGNL1ko1MKKXecVMh1r/wEXCrZ
T3+/RbgcMwyE0lT+yWFeHnsRZHBoFy9fEvwSaHJlZ0/ZR48RKnzFWDHtfZSJAyZA
rZy8CmAa/vJy4I4vRYo5TS4YaszY0qpA8YCYNcNhApORKev/9/kdL9ngOWGF+DXw
L2jynZLgS3nDpSh5mSAc5ddrtgegL/SaMhsWgFEpqKrA0itcoXsTxlE1RrEnljHR
/EcjHJEbthW3u6Mxe2yxA2hWG3rlV7mQLdtB+v83my7bhBaZhnWdps/1pi23PiUp
QIHwQEMkfqTy0WHe+0hEYEkyCExKu6iKs59OqGE/JiGvPF+AtRgiqVVWyRNZvloc
BOBtyY8vVj+p4L+3tB9N9SLE8X5j7os5cZIKb1+lQ+lHj+v3SgEL7DAKQ53p0Zjc
HnVds8u5xom1Ew/RIGOSYDxzawpEqAU/1x+hOtKgfO2FCLaUbcO7iXPh01IeOEYC
Pv5kxnKwSdNMxBay7CIWJ7YKeuSLw8qZHjuc3nPuVaMEUTw2hxWol7NL6C60xzoE
h74Cmr0P5KVViTLgTwbWze4tnCSaF3XjxAd3j5N/wJ7XwYXHR6vCwbLlEgbRFWEm
pZmQ+y6FTCdtXlswM0fY5/Gjl8+5XEE/Jy4Sqg/JSSy1UKZgp10wTph7D8bHnwPM
of8LO4MHKCkEPmy9GLkdOKUq4r5hnkMyhlmaPQVwuVjBe5lTjxJY/XKrlniJMC07
/2yGw8W4gThYSlBlEUWwpNofcWUUG/X5D9e+CablrNedUM1v9zXS+cI0IRVZjJVq
hidSczTOG5PqVUH5UTqMBy02oAKq7HZkz32eArWMApvdnqrw/RSYmW6IBlJK/T5d
j2nx0gmIa6bdTQKCdBa+LUZkV2b5qeOUg6zqBUqZ19ScY6hyqp7DcShUOFiszENM
vUG7UHNIo75uHlxsGi+ws4G15SpXWh7InHgnWkiIxLL40nRBPP1FeYnpudSVJ6qV
FYBaJeOv9V+nBPUSHViuMgj/lkDbY4Z77xm+UspbkS030FA5lO/rQtltiMIoCB9l
mkLBAmQ4E5wvogyre03dbNGzLatGpBcIAltChlu/tdjdJp4gLc4+nhagBlmlRkXX
1rF7B1cwiEQmWDsC/Hz4bVnEqDlpghQ4r1s4p1HgJQaTPbcKMVnQp8l3B8/knftG
3w5R1Pl3EJdBm/wzt8Ul0bHoYiW7+k90cx3xX3SF2asEulLv1MpDpro0OXJ7u+vG
zh03nhqMuDuEZtE+4RXkl2McZRkbVRLnQSJjF1fccTqOVoMlC5miX5GduJw1zzV2
cq/BkhBdvdV51b4Aqj+NXTrnlfTVxAZtPu9Yjb7ObN1z8jT4rQ4PcPVBF3GPGRBo
I8d+NWXO1SAF1BaBdraazWTR70g7RZ5d16eliVCU2dPBJcE8BmqA7n51frQgl8Dj
R3P/SFTCFusnmM/XVWmSdWYwQN9e03m4hBELksm9XKg+Zw8Iv+nAG2j111BG9uWJ
mSf/yCN1mPPP+7dX2aIWaWrDC6mogXAoPa0ZuyI5zEXKiA3VB6XGfWGzStXt1Z2Z
vNwU8e+ErHY+Mo2Wa0T7wFjGbT2rt6NrLq8gx/YZ/wLn2SKwG8aN7q8tHBYM8k6j
dnvOzK7+PnyCvrXA42LAktqJAXWvOodWb91XlKs/T7JI8u2KoN08lOD2xL1bDQo8
oh0IOpcfazp3HW3jlkbvf9oeNd7XWlGqyHqm4loorrUBas15SoHgsuJtlCBPuRj7
R9IypSmIAR4CdFuGf30qHFeDyehw4Eqha99duAICuCnjgA5gQ7mobLxJf58Bvlp+
6cl7OJyMPdxbNz+hDcDwRft8MVsGvNxW5viwzbrdAczdn7IccxgniGo0NVi2o2+y
Jk7Ntb2R74vgnthjBxH+N57Ys+wRxyNd1WIy0hdKjq2SmgZ+BX+5Ew9Kv2Z5u/49
fS/nzT24yApSMWRFa/9IwTuDdbM812OQ5UvqLdTOCIotHjoRAmgXAYFKF+914hZc
COfCrlxVWwS4FYvwbHAV4fFqsrsKScWb3rN3eB/mj4vfNFeju2sHvGIlIwfUfNpl
3vb4ya6aQ5JXdhKUL9AfIxL2fI4b3ida2c1XaXk4C+6/Y+JQEo/hpfHE1EMjWSCG
rZKFXjfOwLfU9EBMBR7ag7ZXZaptgHKjwlo3ZP93SLRmOxLMgFnGUs6bzyGoVHQE
aD09KOHe9tu6hK3hr64mz5btY43tINUFFLNn0JQLpPEkgud251kTy1F5od1BIiEr
kixWR7Nlck7mYn6EV1r6UTesW/pnxQ83GXEojKQv3aqJoe2SpxsP9aNk1XLHLixs
yvBa1qnKYm/ZnyI9Ucdyq3iHBE3ZaTRpUhQ3bVkkifZbR0OsYb8ZXeIfEuyfm/Lu
peDFZ4Oe288zC+vxJUZ2l5Zf5gqsz3rDG3T3RMFuyGwxGwszC6X0sFzofqKWLacS
Jy8fzLBbypRzGpy4nOoat/UCD/qJgvAnFWOUUUMoL6g7kwtDAb77uqUhCX0WLKPr
MrZ6cPYUe4qB6rjgEFjo8sROf5VNzS+IadFnrPBV74z9D4FmawWO1jgEHeMbgPks
k4LpigwNCCW0JAdjAeom1dv2YkkwCRe6pEKO3M4Ii5ePGb0iT9KQRp918DHzJhTT
8KrCM7pF5i8i39oyVJTIJXoEz3AKJ+vOogr/Z95FHCDPhRTW6b8WTtaHj2clME0y
i8ML5ZeiTNUx3eBe6kUtG153HyOTudMRrsxOWD2JbyLsp5EpRTwBZmlopu4OCk13
OXCsggY9K8UV7WTEIdgzZVxvIXtHmOKs44CCuZNHtV4FCVr3SD1vdoO5sEZTrfgW
lAYXxt/d7ObD3mXOFDpJq7wDR+dIIY6hXl5hD/sCQi0Em50BsFppOFz684aB/QD6
vJHf8QwFodBwd61vkoC6Z0FYnzO5zNarhxgXaLFO5cI93MbTjrsByd7qQhNTGiAf
Gq436bQrwd6cm9Cx8LFqgxWbOwlrKds4gOGK/KRv0QZzNa3swm6Ms6GiEzSq0L1o
fU0wWhF1U0nfXygCcpZEuLUnLKs2ttaDuCtFaniAf5lMnZOHjMta+Uqs/umjLxmp
WHqwUIsQK9lfFuYp5fQFVG6J97a9ldYXjHYZxpcdeVCjIeoR0rJsZxk7aOQVHgQ1
jRnthImF1Pb9dgE3cl67gzerxPdc3Yyy5C9xCeHoGP8I/fdpuTFq3PKdcQZ0nB3a
KRUvq4PdiF+Y5jC+9xXNsjCeYIuyg0uPigFbuDleKjqe83fmKTYOB1TjNHvt8Nsb
gflZVL2iXhu0B3e33FF2JFEYFWhSWD/zfGA4gMYCI53sszF+iwWdEdqgaAlmshN6
0kBtmYHrZjeWlSn3i5N6blpsQSjwpW+s39AgnfiMRPfgSGBXbpD+ehSJhAfuPcx3
I8rKdz8dnDY+BfqEfXfcvegEArWHeBJOQo7K4dNUrt5TNidrf3nUv6/cWwyD1iy7
Y1DDYcRnc1VHE5JtvyfDMrZvNGiIb29oX4G0x2kvEHuyzvacS6MV2TbNtl+LEA/R
zesrPlEhUm10H+vfA7r1AttiGDD9TsFJxAGiCFYKdf3UdLYnHWx5Uzcm6uUIWcG3
8N2/wUaGHKVIIX5XTtnaB9Gb8clE0Mr50d5+XbsaIO/8NwvVtQVUGAmIMMinRNyA
jCHWjuI36YbKYKgqOyLCqiSp26EXfaGXCp6idNSegnooW5YdcWhwk//Fj4N49p4X
dlRRiWTLSAGh1MQLksXRrS7HKoQz1OFEttJ6Vk7EZmkRM1DLzG/RMU0UdU8MdUS5
k5O8AHOOQ3ggD6Ad4HAIiZD4bhF33/TCyFnJ9cA8p0Wa5OuS6ShnQhtxxFhNDaII
OpMxhhUAioJiRkzqHggV2HvUUWpRXI4bgqVqrJbL2gOflQcCLIHwMhzTmeiadTrC
6XOgNOwTLJwVZ/Stv+UqCnMQMyg6ugvgAs9reOp1I/vzENUhJhWKrKgGZ/DrrSx5
YjLtvqlYaQA4B8SWWSC6e0AhfW6itgAtF1azZ41OF1N1rSHWOcTxwUZPQjsleCiy
MJqOEQ2Ywj8adkxuZOxUAhtB6LYCBJ6+wLu0lP55PdNXtvt8hZSmZLE+MOyUuID6
KFtPXDUue6MauDR/gAO5YxFVKwQUoN/HuZ1nArApyxXEUQB8L+AeGLMfCaoEvR1I
e1SkxB86/BVpH1aT47XApBF3Tql/6msm62g9WA3gj+ddoRztqMOwP/YZV9BAmdQp
hrO6Jb4TGR7e/YEzeY9P+MBgp9ir89FwcivGioy06zJ6MQ3V8mHPQK0HBdP3VdUM
yhlbSvSt6OrinRKhFGX6x0Xqf0/7lHw4RqHGdF9XHTTw/JzbMVNl+fCR20t0f1e4
dTH94ueHdXa6jkNuwY3KKrN6Hz9IqzcPesLARt7E3omhEjRs3FH/324RbByrbvwo
u3CB58CxZJL8cJcSq5R4T0t2zQyGa8VjANalntnB0zHyu2GxtZKpDgi3LtWYmEeR
LNsPDv5ssbzTgh2OdauoseN5TF7rJ0plRgSpQ7AJ9zi6jwB94I3p1gf44Xk856st
HslihAj4QFkFmoA3zzdIRS9TLKBKNLGfap9GyMaWBjC3penXiBQpsamnDd0/Sz3n
lCvyoCKPbRNcXYPNXbHgh9cwkrNhFZ0LcEEdHWUAhNVtLdiatiCk0WN8p/1jz5uS
fzZHf9suLgFrOfqQlr9cBCd64fDGv9A7h6OqUW7ClV35nmHf/CWcj3awhmSTn4vP
P2KkMeXjlEv3658CU9lH4BCPphUnwYcpWf7nZT5f5xkgdqFR6yKSVMb20cvIYi/s
B/YALyjJ7QG2GWAaEIv8BdblSNGOyPGj894Huj9cbfR4ez4BxXXU00FACoo39RvM
lXXqiGKMrSHUnP38ZqjOpEgUYeu0gZME1s7L64nLPVygv52Wa+TlDw4UXqIrR0kc
M/Um4R2YDevFuVrDpPVt5RTjDum5NkbdYFdMWQYT+XRDPEMt3WXRMpgKCE3cOHkt
apQ8SxGRL018NaF0vJVPk3SZWhijkZnce6EjCZ7GxPR4mESrO1xQpsi+TZFWXg1v
+9FDeOJx4qf+1KOmKS8+rLgyEGnc+8GBetQNxK/6nxI9IG2yG5uDFuUBzGwPx/wI
RKyX1iM6LeR7FYnvenuzsVN3TkGIRwWzEaq/SL6wQz04GFtV6sZmfwmrY1T8KlS7
cjr2vYK1MIMP1Z1/CR7BOGqVpA/gedk9B03CyAXl45UvCArKaoS+ZyYDWDOjwY7z
nC5MCgQeM+hIVGunp2klup8ggEYNgf5837D07c+GGqwGpL9bppwPmZsg4jcA7t2l
QSeY98+lSOt/KgZona3o67IM8x/+g64DLNIxWD5JkgHf5yvYuReT3v8o1JGbCcwD
UrOF83sN3zwdfC1oUtDANsqwWqZHchzXDtuk793e8RvHKJEaNJaZDDLhgSz65Lrn
/13LtrxITTIwcDIknX8iaFeYhukSQ+FTiddpe19hTNRPXOfI1eboFPxK2fuZMknk
l1f3lv1COP/kjrAuvpdoXKqVgfYcVsbDMNrEDH5t0luSoYt3LyJmcajAyLvZe1b6
unUGM/jVxLi4PD+go7ZSnLOB9S8QuWmI5r/c7FFyZeR/ifbzxMS149kRGEDA6XYz
pjL3rR4wVU5eZDnrK0H5THMsqahlA/CBoFd1cxdMAM8fSZN54hfi1HRQ4PoDxQ+Q
VBjSd2Q0zE3OB7iqn/SpcHKUf6elHpF4jIdtYxZX1esYrBvdLkkegY6YkbHuMSjm
f0ysFg9Fg4k7FsEOqQX5wV+5kfBH/VYYtPqCJIZdklbbmiXn2qO9y8ZUQ5stn3pH
3tMqQ1AFz6kDJDYrTq8c2NFYSbevNxFXd5KJacL+ayQ80mrNDr6o45SJpMEz6sQ6
/1pZCeeocoCnzHlqjRObDuI9AaVsLqWqVF8G/q/ZUmrsQ+VkMQs9TtD12Jg1f41Q
NMIAUPel3lgmlN1TOSDMbnBFpeLyysgWX2YQcggp1130+yFxW6GR6I6e1Qs32ODn
9cIGiEllWcIOoUAJPl+5Hu9RNRpSzrbhYz4cOHYwrOpbJmN8HW1LQ9qNvvYKMv+G
/Bs0+Ry35AwQT5/kep1Jgo0lsBoznbljvDsLM3GAw6cGw+tr/4MOxbMGRAOkaZBg
+CQPap9ItNYewXdAv5Qd2jIgfXbgZL228IxU/s73l1TzY1pUYGq0I567pYOiD4xc
xRKswursJ5uzFx2jjuGrlrmX5rP/RvJa7DBVWdCBJ215Gxz2y1V9hf5m5yRQp05O
rfy+r8MBFev7RY5e0khz5otW6YtW8gHRnrAgXKHUODg8R/7aPUYE9aav8R9UWj7b
x857Bsta90Q03mBxOBBO+OrfkBzjp+2tCNwBvgpa9zGI7YmTadW1Ecssu7KzgNmN
+0pkptekhaZKUQGKM4RZehpVU/9EPPQ2JB3RlxoBWGsiNm7lIs9i/EpK3FJsFLJz
XghqrP9s9jMpUg3k5VTb7bNDs3SfPX34UZ0CG+evZcOkvaIhdG2nzHbD3MkACFUf
IUHV838IL8R9+UA3+Bt67UTrfbNU7CRiHBboc7GLUYeNi1G/0XpWIx8VjeHWHS/b
IRsKXIIKKhdN6OGmu6UItibkiogELAkwq2MLkREnuHfCKVn8Rwb4xCIfZ8Y/reGi
nbQ/wx1LvoiAMPPOu8tWjTb+43LAO5nt51DK2Y9bImZ0CCz4YHKAYBxIgJHD/qsn
ncHozVCoXb5oNNik0KDx4CIKAnIvoszPA+PYILRAqIPj2sytYtNFx85NCog0lHK7
SA2RWlE5IoGXQQd8x6+4MF08P+m9YZ/HkEzST3QiAXwzdFPPm46aGHeJjUtk3gRf
0oGxTiIOWfyMtn0KVthHdtEkSaiOvN/3R+15eWae/aIbZHd3SKT1mE6VYRfqZWlj
UzzoGsVTSmeGnZSr83uvcP15N5XKAX3q2QR6RttbuIXMVvl8ec0LOoWeSjpFwAUE
lgsAH5b5MST2VFYXHV8V3zwc4wGGh0O4dBdTv7MIvigLZz7tBxFiaddgxFq/S87q
oRlqWjV0fiV5IzzPMIgoP6b5cOsD0D/navOHBW3Nur8crD2nXhIH1DSJhUQLPSzm
MgJ9InyaD6IH0FS5gBqD3j02Sr3t9D4g4oRMizZpmKifOL/2Oma5+Vg7TCkKEN/h
FmFE3Me7ZK7BHY+HR3sq+mqIn0s8ZM00h5umkaQDAvL2Y7ajgP++LIrTFvQRmEsw
q27jALQMWX2vema2SnyLTwC5jjzv++u4efgJQdzRSZGB2yaaOCH4dLQyZq/fZNNS
2N7npwnb+m8VUUTKUIt7UL3CKkn9/D75fAMy4UncbatliKcD92U4VAW21O/GIsJn
df5knLoipUWw2ULj5FrH79l7/kfQYz6cSMrQwh8H7kazRyKUM2yW4PJJJsuF+eMJ
dREls1zAtBnEaALgMA8NzAoWCx6y3mChk5msNc/fd+AME0ge3mZbIGbF5tCCxAM1
vJisyno1Uj7GOCNRs2MAMk9qwvl2CejFCO9u7VA6tonpFnsrN07NtfH/ZJJUFlBE
bnA54Hh2Vt9mPO4GObIQSPuyE1mXab8f6/22SKGy471dSU6du6dVxd2QxM9kFDUv
Yi0hAnrnjjXLDol1ftpo50CJCLTzp/ktlNO47ywaCz+k9dssTPuNZxAvsRBj5pZV
78qt6NqfhL9uox2hkD7x4QYduJj5ofPOrlql16aiWn8j7tUI4dTptOzGX4Y7iaLe
VwpybcaTwg62qNTHa2+b7My/LPMe6Xd0lmcpFXFmkmzIyE+ZMZ7B7SwGE7jzUv2y
5uQD4DSGE2sbI5uDahdDheL8lQgWyHaJvWTsMcTpVf2Ay4KbLkLvq9diVNecHQm6
k1UmG+trBbOpjfe3dSARVuyJK4JT0W5ohlbJgqKuH0R5hyecEoSJF/UoqjX9THt7
Jfbv3C0ODGIEl7Rw+8zVumMj8xegJFm3PzwzBQq/7QTRE1emnow7kgokz58D4zTJ
j4kp+KhHdDyAdsqyLLH6sAGz7moGVLIlFstvrd/mF5dwHCu1Hi9JM3AsQRo+7XVF
pqf4MobZB2PayOTl0fZkeaCdc4tbnQJrvdv2rnDsdnTCG1TjsvYFfKQSpc6E8GTo
/lL63+nSU0lJWmDWfvqyVNIzm8L0dsgNZplNY72ia1+FqCSvYxCrSm1ES0er+qLl
mV9WvBETACI01Xa/2ldxrUj4Y1zFFe6Mdpy9sh2wApyXY09qJr2GvG7p+bEkaYFE
GF8DXzfdyvY6eU4IXqUwtqWf6t6/PXh3fHpR9tl+AnCyXpJmqOUVAhx1YHxHWiIm
jzLb+xdVwmyQn5RRl/G6HjbHT5/0uQ5Xoi2x/hcpqst8EBUz7qdch2SZsu5+35CV
PEUU/q/l3SAqK/i7kdUGFbgIKIjZUxDknxhB/JTEI8WdQVZsdz2eTIru1N6nRAVi
ex+O8QGUA3aIB1YdEulSBfTx7Q23oL1rNzDeVZX0eCikYnXmImNfBuCdsyI3mI6c
BD2QHifaawplEyv8REKZdkibYYHDu062u87iujI93Rjk6RhfO2/oF305kuQTnHx0
qnPVxP4SHtdW4fEF0Ga31YZ6ie7TwCgxPINITzZQfhN/URJKdwp0r4swaawTNSop
7zmW+RqezdC6EPu1s/f3lo68ZgKQ/tIK7VrnGkBiCbL/wY1Rt9I3dPDoLVWVfM73
27/F6o5OkWwHOO1G4ao4kOvjTuy4MwqOHzWZUgBA9wii2v0kChVA+wITmhULFDVD
x+P3o1/kfXI6L8KWd6xUjWWPVv+fStp1VwPnFWVmO28wWdAqZRKEp2Rey50i9/Wh
/q1Tu77ZNBkb1pEIWZZcgpDvLYZE2Mr+nJAUW9qcnMjxeRwkt2Swk17qCnLGv/hf
vgB8xrPJQcyPpKbJ0noI/tWPVh8Xi+47NYdGdEZsTLeJPyWZGDyIHsDDPVcdSo2R
BKVh+koB5CgcI0e9pdWmIs+X0KV4ZLCABGy+c7iMI1r76Gx75Rheij5C/8/qXQE5
lATjOS9oBY+1YtWMw/MS3kD9u8PmhB6wDsKOs8OB52WmclOz4gH3zUa/wBaIFxWj
9tdP1SolSsmbc7RA5Au4PPjKAkoO52S/xu096IdNNtZCtd9PbM6XD2c4Jxpmmssm
U+5U/ffRm8J7oYdluDU56B+GDw6GJTQZJiDzWZtkt8Nni90fIskrNTBFFoVyqk3P
zr8Ney8ThJVTwlvM4mkizrPpL7Du6wU5k1RIwWoxDCikEWw3vaJk+53NPoODqe5E
INrM7eAu9p8b8wpnmMkAHxKrLI2MzGZ4ha+bQXjgb1QKhM4oRUmwJG7IKRlHrgil
eDbh9D7Q/g70rTjzPOsEqomHQFQ/iFyc3ObrELLKq8xK9HrKOiilyMDSx3+2CFKC
QJSrvpqhKeCdGd4EEj/teQsNKJMyFi/5601RG6E447dpXpDUcwgpoHNuRKkwuD5n
amHXCy246uMq7jBw3amexzyh5B+YpnaCdbgVDY6yFbzs7C3CZrtvUiQV3ZcavkdF
ht1L8Ln/nrUix+k02MKtHTLUz5FjdNqYhMVyeOxluBxPFb8jcFI60KY625AA9oPs
kHT2bJU1lyse4aHRUx5g8NgztseNbCtrR4nus2yLZ9z+oKfeQNyHTeF0UMOXtCld
neCjbzl8Ki6XvEvz+H6jWOjb6j6gnX1T1kRfojHveu4gbWeqActUyGQkuvUCHSo4
/gnkFMxYnzsmndZR4PgXP+qeUrYYXzzAn2bAU1VCeFwzTF7HWTkEu5nCYpMioG0H
NeyhWA497Z4IGUuItd9gC3mEFgc4gqjW8nH2BOLcrI7IeYP6EEVORsPRxzzUXLCi
yVnF3YozZU1ytDUdGztK9Dbj914pyFCWOttKcdRlOxQB8oGC3iNVZ9KigtjcifiT
wzs+AT+M3IT506ivM8p1BA9LpaAaO/w9JewRTTUjBxMmBV4i4qsmKkK8HmtPH7nT
oeqyvENLDIloQZx4seG7Qjooyr8WgCsg46gBHmE7aZwYFfWB4CM8iM9NobHD0Yc+
tVlOhbwLUCOjE9RUhT85yTpRsimivqXRXPpOV5gjercNZ98/AlQzRQ3dKaL2IhJ/
AUM1n2lur0+7QmqYVWO9g1gQLxr3wsDDZdvTQPL2vjRXqVX6Qbu+D5w/u1gaXgVM
M+T3Dnm4V+konCrKLjscJytM1ZsVGBSdwOVA5P2AYMwwgGohn9N2SfjjsmVd6/IW
lGGOBmQFRuyku91BLxpgL5ypwr/vor1LhWhA77LKx3E1bGOZJdlcygpqYjQ3mFXL
3Wp0fFKtkkpvx0WOX+eGEnIggJvJOganUTx6nnbGrQy6KrkzXVygUTvAPpMhcioy
89sXnFBm5jbRuBKmt7EEShZPlWrZ2YoXTl429TMQTHSQ86+GFzgPMMvcWL+E/7UI
HlsSd1igUQGpUZSe29AhzUr/xmV2iTeAmsf761ldC5L6oqMtdTe9JlfO39KCeHJi
DgwpD1YComSgqy5YBSga3Dwa+5TU0o3ZP+Jr8KBNV+ng0An/nSBlXvFJCPGNEARr
IN7kb8Qg+5ILMmnxsWfFaErbJV4YFVT5FSSxESOhYWOh++KnPKrueZDQclFZKE2z
hUAd06Tu32Dj1p2qAlGzpbgrQYeFpq32HOJekTxmENTjk/Hd5kPUo25kcppYKuQj
SxWV4dmfkY/brSIa+n0Y6wp9isFLXvKjn5mtgD9xnb5Ejr9MRt9g6Sq2FQ3Phfl5
HmUqgfkJaFFCEHYcfWpyZ6IsGeOeTJeb/cxk6uYkxuRMu63AZYZCApLti2yilGg5
wSzYIQaTY4TLSG8xKZd8AMq4CfFFL64f4OVGJkQOYcRO36AoBP5xruFxEbY2tVKL
PozK+Yz5NL8Q9r/8LAbum369tq1/tnk/eArTyEHxUwNbX3EBBii8pWhYy9btmcfz
7UB2tKfZSmUMGPVTbvt7uUy/vNAddKKH+AgKoIwaD/5fbHu2nqx0Qf1DLVxh69oO
Jmkjpk6Ja5ul75JFKXsx4ajxpB8lfWe0+DWlfs5Xd3hzprD8td4tp6Yq2JKGR4hA
3zR2X/3Ia5iv7zC7Coe+2moDhjG2wZbAqBOmPSw3w9MjXF/FJcQ1TI35xvyaVOq+
+kzGivrBpkgDK2BZgj7wAdq1wwhG/OHnGzEQIPAwEiTWSPzWtR00piWNcJxE5drF
W/a5v5s+lAHXfx3KrZMFuFmlbKr3yQH8Vq4wNMrv7zYHtZw34xnjrBUitMJGtrVs
0EvIMykDQna5Udi9kKEZji/D6aKHftW16jnSKkHUoYxWvxCdhsu5jL66wUA01joT
FD3rJ/O/HdLHUSNkAyBJr+2rUKx7rr+lotbuMsPSUSOLVn7eKukYwOe19DgUPalW
5ebc9xl35DaWTYjHuC6iGCPTSC6nFec3nVxTxsYLaLd9HKuSUTP4pSadxPwKxkFK
aDrhuDuvgkiqm14U2DUvcSdeeFPBMptaPZegW2GvwMSxnQQLSseJpC3oG/3fnTbW
5NlDiS0RP4h14AbJLtcRxKAwCTgOFEhR0eCD5kkVFclOg43l8ODiQdPjIwLNq/RN
LPPPstnmUCukl4zlSj4T2cp3nZ3rU+zYxMwpkWFGPOwehHuhznQDsltaRc0gkvbi
gAfct0YbXzV782tpFT5bKhafkCbkr7W0JyHemc9jua7G07ZgysmVJnGF515xgXUg
c7Gki8oVZsXVzCNMhA8qMuMUjgH3svnjoPCcwoIO5BzmYadIPlKR13rBsFkKM4jK
X5s1eUqN+X8M+DftTJaKHKvT6tKRRo3arGoVeiNFmIvnn9J5boLxZxtjDxt7k4VS
TvHQ57hBHtd8byAITmTAxYL+SzApPJCDZjLVu0iVd6WNlmveaDX6T6D1c3qsHxlO
3McDBlluETC3BpLpHxn0YD4zC/Fg6rQgznaQC9Jjq8immeoTp842Q7bPqxI3lm5R
nIuHUFgGQpQvCLokwg4cnzeFSm953C0QvCz/JnCKU+ojTBTtVwiclKD/acU3nB47
3FiUMDkxIbYyjiBc47AMPo5OpgmToOwyaUUhXTfpeSpFAUm1jsdmAH1I6kSDykaK
bAFBqSC6j1b3grL9uXHtYsEWZgX7o/6OGjv0wH5ltsbWa0ZAFqzQ/jkUNVOLuQzc
hgbF1HqBZNGkh7WHHbVCcodAnqATMpj1mVlU4EnPKevPVzQ1dNKJQudb3rwtefTm
Oh/2sNN408vfTZ4c2JdxAg1tEJQ/GmY1UT9ok1MiDoOgmCeB4zPHr+/OHhx8B7fa
SWjJjxvgk+/NqlEn+rwuthjv4hSD7BBlNUWqtLTLc5uyUdRcoEUwWHGf1UYdUsEG
tt77HVow6aBdoV08AcIcO23bUDhxR5eq7tLCHPzfs11yuxfoT98DD5uCMBTo865T
E7PfFs5T3YQVTFwzxK+S6ctyQ6e/y9Ai3wswAHBl1j7TUyD+qz38k1LSUPu7/Jla
39YGw0RQnnZebgLM5Tmc/Q8xrmp//rkUI4RmtRG3lKEVIONvWjtSVjCjAbHZqZV0
12uEMekbI35lP0tPpTvGx9de+TKohBftyDKCdX4s0Kw+UqTsuwpUOWdrnlyAebAC
KPuC95W4jdjGg54EeV5C25NlgERuLoNzO0eXZhsieZhisInZJZ56+dAbCAo53izQ
wtccNwA+KAqQBirsrUYgW/kS7411RI3rsGzIrublIiZUFjJkZkllttykiog4nn5C
78oPo/qAZoEhwqjbtLb9o1nvMQmXQZ0hqRs7C/wyoLjmli7TbwVCoh5chUK3sq/Z
VYBmk29zhS2wUUmv+mz8jvxNC2X7qvqgtHyFN17DTwA6YzcExTk6V3q5SSbGBvZy
hkNiCpBqTDuVa0v6ed0aS65df6aZdR6xX+hJIIXuksXTTt6nc2zKkj1BrnmYZE0q
17FuHoP4Tf0L17Rk/6UPG4Dp3wFVE91Ry/OXFap3aYea5Z4xbOAQwG+oXFQzdGhv
FlUKu6bwDvzu7qWlSO7gSqjJOSvdozliwD/JDJsSPoyVnqtKKSZ1bf7WI0i47nqx
AL4mOXyrBx+ZDVC+7uvwMKu3d8+vsYqYJIY66j/pucRKmeL3DeD2zXxkRmrnX3Sj
aDZy4a+k9TUDeVrhesqC4F/TxF3rG+4UpXk4Vkw416EFmMoyxp5NQp7ma/VdSvvx
hzTx2pVmu1h9zOVxPbxSGM99tKb8j5OFPytiHR0GPKoZ5Hepiz4TvdKSznpaIJax
65oI/GwRoWJ/hZZPYh4mX8bqbcah9SVcD/aXh2oRnFw4yBhcxZpFXrtSI2J5qt+v
hXn6Qzt8VRykh1HwD9khGAO/K7+vU5a68ark+s7YQTpoxqxXqMY+Gs47pDAx8oqK
aUg3UpS1YLS0gl8xcvqO4OwP5GbKHZgnJEABCKKn/uQJYmrU/PdCD7eHa6lm+z8Q
+d7pHpmXa96rEeBhUJ7Yjh2KMZUqQsm7tf1Ws4GqWXEIconrUTXekVa8TCeP25aQ
BZdqGDDX66b2FSl9U0kLoFA3HWcYdxDl3k2YiwUaAunWiVV4dSCN4SjQjlRRki2P
1LMRQQ4ruWxr5e5ow0H+kbe1QQQwvQkxfewesb4+lew8p45fEAbXJfRFG5SXGGpi
Qn8tV3BL8A6aEp9kgae8f3JSpnLlrE9KN9fWsh3PSB1nxCQ9A0o9Jrmbg7bk0tG8
qepPfMMF4n99vLw1imTHdOTNOQqP3Z7ETrzVd3kUt9zdltOUx4mmj2nYzo7v7mYa
c2I9e/y+TZW2+87U1fe8DqCchfSj5cPnQryuR1R/Ajr9HnM+lL7bfv7rFdGn8Gex
gV/ooGfoBgQKpWP3OB/zC2khv6UTFS+xIjzj2gh8Yyco+Wsloz8dfD6mGcxtKuxc
r7Alze1gthbRDioNoWmFjDfcyRpL6PZ18NzqrWMiJ8zUUjVgxpctvEST1Km+16+k
jL7ryqBk6Npe478Q9kZMGuJeYtCJaCXwlHh7XWZSa+z+lMepCCOm47eq0JNlEFuQ
ZxQTzM0Hv3j3vsgQYoT2gHX1wqYbtXiA7A2qK+UK1kmbUJUggB5eLqAuu6tEzyzv
3YrQ56fwfxWZnr9SunDXzeZUS9beUwWu5Yg3JNxsU/PKLNXeoIZxe4NqHRnsjf/3
Y4dZktGTYwPSkBmpTtbeP5FhaqskV18WYc962HTlCyz7SOgsaG39vpZ9KrRUZ3bj
wEegzBE8hzuQzzYyRobdCQ7p+2TJAydwslhDiXueUC/35LCi1jk447l3ss0h6Gcf
mhmfC2HUOhDzt/fOLkz7GpKhpQuHresWSVHyCUabSSkp2RlUz0Pbgyu6SLuiEqLS
SQsgrSEZkLXZ/lySU6M/yZAEBYzpKT8qOaGHPVzTKLjD9BmXRGc1W9W775JR5ClU
t/WYJ38BA/38R2ZejGTGBzxYw+hqO3SoAIzOUSs0kkKGKyth5Aau+P6U+6kcZL+9
G1wEMqO63mWTH8btgRJq5sEKK2Ow/ZRpbn1Zbh9QeTwqh2IISg9CsEWaRqn/Ayym
ls2AQZ2kiyJv79ZNbXoUgMRAFxn/urs6kQuLPjFcr6LdjXsR/XMMdMDe+WyajO/b
c3rI6G9lcfmMY/k9Y98nuC1mrkIAQNNp5HtQN2b5HIrEne7KlTWTMiIWtnyM09zS
OXYeyAUhHHcZZiVgVSGdbEcElRUz8zU6f3UCNzd66D0OB6i8+ofrD0u4goMO3Cqo
dg5tB9W8ZYOwidypgPOK59fJpGI4TAUtg32ISPsf/JT6g6b7JbGhRn+FRs9w/su5
eE9iVo1EImjxXJUPNLmk+8RwdEmICFu+NP+qw5MwWWjFCsf6XJPgMCLi0bXaj06X
rk1lCu06h9B+TgUG80wwWj/nYX28mhLOvg5+b0gej/y1iOdvFTwGG4kT9O9P4awi
2hIqMhjIte3beS7Z4rfQ1sswv92RLDdDbJoLVoXgy9GmX2J/uYswd8em0eny8Qog
gxptIpwESLaUWkScDqDOPL1zlIE2OU0XdQjYovxewNMHAKw1S6Fdvva4Ud0gWH5t
1mdGLNBYWz0C5R9Hf8k/zXvj226VwFhzc4Lkh/fOPW6pAqdUwtvpHkusMrmcfygP
awEyMxcibVlzHZr82YroE/fXI/cCgAVO5Yjz9Tano32vgRYX2W8SxcQLYZGNTVAC
choApxNKySkusIcW5OJiSmTWM4ucHiI3AYXU/L3dVi8UFpqLu3W15hfrml/iqIof
xwxgzgyGvqC524tVK5hAuLrKXx7yvpUjamcMTuHS5lhgHBPrqkpLHNh5n0tFm6Rp
1pmAUS916iA0tS6HIFTVLAJkUZ5h2K1X6OgZ/H6rRCb4wZeb401tKJsrrenbX+Wu
fr1QAK0SGf9/ZrMm9J/43N/OQDnbYyEB4kqWPUE5EYfGSABXSdZP5nBxktAMgYDr
3+sNw8ZxMDQC17S04KOg90Ta+loAxP0WQr9GM14f/KjWHboui0T22Mu6dpaWaP4i
JyMcg03QmuLzd87NmdfEb27+B7Iq4UwS/0Uj3ITXf0jVTV45CcU8AOjj+EnsNrJm
N/9Kj0QRVZ9P0u+qo6aPcDoJ1K6+4m3ivNZaD1RKgaj6IVkQMfhYYYjEezCcZlHH
6/j72SYgOqyADSIpmFtZJJVOrDnuK8A2txvvTjyZTC2QTU8ftrXRpnG84rvKjKTK
yGySVScX38edua3FQwKtpQXY/eGOrxpM3sQtmlbslsx8FxCubfKNaEk0OCXuKqIa
6iIis+SzqZDqOrAiDeBRScB72+9PIU4rvhB0vIvEC3oDWza9TdQcIPStjEkIwxur
Z/fO9sNzUThsMmDJW1cv+b38NbJmafdjoGYmS/K5lscmz8YS/CK5njznv07p8UH3
Lvmb/i5rxHb5y0JtNpdMB5eUjFwq6fVScTTEpVGfzrZ60/P3rRFoXZ1UIoiGfOCN
ch0uCz3n+CxOTW/33PWx9JuoG0R81dMZSspGGzHJyGNdqqoiuAqoqb9WvQRWoLDZ
W6Ize2ruvwjW20qQJuvHuTLmTsnQprfH/gthCxkknbjvh6nBV88d2eS9Q1vkHRcD
/LoxiSvYq5Fub4GdFexa+EdqdfNxrH70+Y7EmFQF8rdyrN84vACh1Apc4cmKTLKW
26cf1/Rgv+yJbbqr6w0Jha9Q1xOFWz8TpCVfM1VilEBq4wvwXfo9qin8Lt0J8jge
iDNiB8aNeIWqpY+WFT0sHvwl4wEYGks6g3y4ZmYAb3Wp0L32MPJoOP7l+owJWHRK
2T/mEmHFLgle0H9GGKpWbFBXvUTBRsETxtPrtbU4vELjWukcVcNTgSD/dOg2zrJh
UtjgstGkRngdypxUuBGTcje1cd6/R0td0UpSvCwoFqIG1bbCc8g2ERbaFOB2ZDfY
yydPvDNb1El2w8E3xfcj5GJSH/VH5BPgEvrS5bHJh1+9o5vfd8kOjYBGsBkuvjxx
0TeSBwsBaIdFBRu/L4HkN+69vol+UsIV3s631TYud6n1TCUsTNqVqN+mTsxhwfcW
t2yseUUwLBpHvSmAIFr3nEIwA1y+ky0RVEpmgrB8QU30y1tsr38qkySI1R5r61D1
ZPsblqbo6M0Cn2//OPsrPEmlU6/kK2pzpdo626UIPxjR4gqe46hMnymUj3WfIdVY
7jcCrFBk9s47NzG3GAZkjjvylyNbnnNK/vC5KGMr7SqAbFB92lG9VX6B5fdE5QMf
1iG1fC38C4a+rJy2CprFM9iKE83D6cQ/5LKkmEnLS8dh8e4Mz97QUlMjWeqpWWjb
Rs2gyeyI1dUV+Hu7UFTVBMFy75DOGY6k5CiamehrDcMllpy1dVA6hn5QxPr9774S
xyFAQVf5LsfDTj1LGfkiK8JnhU2EoERMLdgjZSjBBQLS1SXzGnntoQ56CrsLrZzf
K0FwIjqKG1BX8qcGil4Zold4eihB2eppvifzIYYJkQMh8vsRUsGy+ucS0remiP6C
dJrlnybrtf+DoEX6KbqmbUrBtKFygkFkvucuIcUJPk9d8fIzaxI5QKWxB+FQ3Umy
TGbJtWRmZpY0FFyJb9ZZFeJyGE5ZysORNmDCksYIZCjffMeLPkjMdNb3UAKBJRtP
rX5zBR3u9VXkzyGp+w1seuuPOi2oyjFh2Vf7khNE69OGevMLe0x7fpoyRXfdl0G4
uTMtP9V9cfczutjkBy7Xsv2F+P9/0tpmNqrWrHEl/Cm5Ee60ak9nqQUg25jHqvOm
Rp3NCocGN2NvZUcS7LH7FbyXH062iUuTPolEfIsAlbsMsvNU0JQ5qCGKMTqTH65n
94ydOeJL5SP01bWXRw8A3uEd6bDeEteB5ugirPY8BuG3s/KVMsnaJeKz7R0ILQG9
UeyozhhdEB2qQIGspJ5hF2BencTKQZqa3rYg5hi6QUTS2fELaxhyvtZNti/5C8cY
bIaheay0LXnN0KQQCB94LQONDlm7P43tzcgs7jvGLRq/UiboihW/i9/qi9uxl1gc
Dz/zciMB3fbsWVk2QDIEJUKAmbvJB+gpFQlxPh7nRAxCcD/4dWBcChNW+KgSjeOu
pGfIaVG9CGYMhnUCEOfK6KRiDgfk0nEKtUnLY/+vDq3GhFZtEGTU6oD8odJFLFMm
dnaI6d0AxImEWclwP8jK9FhfkD9OuAYHT+/m/+mgsGgL1kHobAc77m/5bYWAVCLo
hE4WAVVh3JWJfYX5K3KaXzerKv8LntNbFOeB96/NKeYnJuvT2vUjE7eh+x+XdYYc
X8NXS4wtid37mbcI0ru9lFiP8SXUNUUx+MkkDRNxD0qtD7hX52eTM+nYyIux9OV4
vG4Ilr4SLo4GHWlEcWMO5WfnzD0mh+1AY/DkzMFmdaq3HOQd+FMfs69HnuK9L/0A
rEBotfdDfc3pPTyMhf9lsOVkTVlUf/A9ZIRg8iUdjYFFGnnacwYDRc/TrwZojRfe
M7NLFJsN4K7O/yQZ/v7ZlR5b0SaK/50QPVtDYn8cbKy7Re6KUkDaTej/ymjYQARE
SU0h/mzSdmkJgepPL7zDrPdFeLX0Mci+eGFy4ErnwuaNVj6lFZAb2J/GCvpvv1AD
cJ8tQVLhJl78NMbnYs6KJfAmiysPu3KqbVUvMdwcjZtFPO6+jLeiH1XIP0dOtO7M
VuKnkH8BtvMuQMTKiNv4U2AVHo7QbNU8dV49ex4c/2kd5e1AHMyt0Z+13lSlEUpq
Tx6ZtdUUza9Oi/IgXm25cfiY3D3lpkCa9GwfwKnOp3Wmr3vFAC+YFrZR3Trwlq+c
DtecWgfWI+5BEh04wKHfBcOaYn/c0dBfaKW20O/91C8=
`pragma protect end_protected
