// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 03:56:19 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jz3131TYG6ZI5A01YxSre9SnG7BBSDaxA0YcPjYZ/N5jq24hTM3t46IAWWxFoP/m
fKME3zFVthmETCOa4WGqdzAp/jDQKXsRS5qzvBSvh1QvLL2hUV43YiS70ClyV5DD
oQ62bu6JnQMVYRuENsuo/G3H+z2kSQ1GxInZKFuxPm0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 48656)
nSNQ88ejQSzOoqpJEg0ZMvxKe1Cnym+4HCN6tnp2AIeDke/Ppw/4EP7uXWuGZ+lZ
74WaecTFyCOiXP2qkHlJajX4yaiV90C+prEFLrgzCGp86jy1Uo8Uky11K1AhbQw0
hTjbaOIhz7y4DY0NJRKYX5hzHE8WovZ58S/U2Qp7bH6SL/z/MAemUFQZFprbIUJQ
fkDeNILR8r4gxfLV43PBRkVwJSEG0udlg6dxVU9bi6rczsLtemiiln0d3dOrInmf
V6vRFAZOtRfiXfP8DrNecXThRjjcikiXfaRAKkkRPHjM6P2yjlPNDOn5EWdk/EOq
1aJn+Xwd9wyQbTWV+EcjY7naz19jR2mqaQ1nVp75hb3b5a3WwsKAX1yzQnX5hlKY
ufatJ3ppjzqKffajFg1ytQHhaKteZ25pSlrnE89flw4tL0Sk302pvusomH16kEX/
GZZg/Bs5oLZDVfhzBJafdvTkBK92H90N4WFuc0dDcmWfRWtWdUmMs2nMzuPhcWvz
2UgdSwq+U2lfLq/fhFAp46Iy1qCc1u50Nhz7MQZom0g2VAm0CHV/0Iv5rM5/UsIL
xIvApRmGdW90c7s2qTWRd8AWqHIQHG5PAbqMc9Qbn24KzSCQuCyxOI/sW2rFt+hi
f2ER8JPcFBGAQPGBgqljNMkDVgXQCgS5jUVx+/aB00WTRQEZysWLhUKM7ucw56c5
76HGfYJ/alLxER/NKHzxCeBPlk7rcRMBf9KxE9NnFJZImvOscYgzon15yHaq9kte
ikRo4wnzihTdgmrzVI67/Ki1SqG3Qv0TFTc2A2K/4xAAr0XLTUSzI52RfPCVVr43
9OcAZUgOJwscxmV4InUXgSwRGGQGVb7sWEo42Cm0BP84YWyUdo4SzuilOkynRNXO
NDI8uRUbKRtepeDC6ShXPogKFPSQNCfZzEmVQpQzsk1wuVrvy65gNwpeh77+NuZh
3TIS0PXlpUnTnJ9+77RnxvcRgCPP8gyitR8DGSvrYdIk22KeB1eTYTbC3T8ILdfi
YSSXV/WyxGGoo5/zzOV3sTGeB0RsdwXvczvwnFseQaZNPzuW3IrN+3+iS/FsznCZ
4Wnkcyw23bNIyRlywr0GFt/zwJz+mfKbWDIND8K/G2BFOI2Zntzxe6yiNnQr5M5K
0W65KfP6kUByHjh/AI2Cn/XCQuhE3aeUZNJzpsv2BZCohjZqEq1C9Eww+AeDEAf1
IlW3oP33/dzAEoiJld7QglmGkJ6exsVopy1vYxe4sqPJ+nyZ/JU+GJ9TvoJTrbBy
Nga1fcFvhk9pFeDjcFiqPZE8zxRcIzQgx7w8z6qTUZhEQ2xA+jn0tNxlkBbSpK9K
wEIhpPjmVlf0vlJj1i0uVIHMncLzgm0P8g/JvIaeZq/ZJKFT73AbQU2QvMjfpjGo
Uu+hAR8esJFzpYTNIrM5egmPAykIbaRJTYUSKUh0wmwcNhz1RByH8BtUtJR1Qeew
9fwndm0vG7RCk4xnGsz7xlVZRq5N1LNWuVZjJrQOHDRFsrSbmp1Ktcka0Opvv17J
w7HAz0QD7rPFrY2s52DpQQGdxjBrUXgBYQfjQzi1sG8cqZQi8nnUkrp5muVRL/Bs
i78/yT4RlqzaDoA5Xrkp5WDt2gPnnd6h8AKVpOOmMiDqPQlSWTP21uArgSTOX6ac
/0LkwMFM6zyJtcl/rq165+Rwm61xv0YzbLBM/UIP4pXf9LF4EjCqvfk07fYLi74I
FTY2xboa0LE0vAc6fbAQYJMtniAk8QzcuSkKdhHtDwo8oNipVaC0OrVrkCY3tFEn
tKV5p4Pnv+2BoXinngiSGAUUGak0AYT6HjrfgtolLDS/W+Ib1M7FWSYtFItS+WrJ
/7zo8BMTQg6NajpJvJBV4+wxteYQU6EiKg44F6hoNihEmC5VO0jtuV12bKYypoVC
3BXxYBG9qkV2lOBhIFch2ZjvcRJPab1g79viyG2uZ+a7P/VLyFU1vP/sYfbHbhEe
CF29XMYWSvq7EDKQIKU+rpYEaOj1fsQFZ9LbaPq++T/MiZrzVehyHn493iDQ8Q9b
nIWwOtCwGad8eo//KE7NRiuoe83Tpf0oY/9ESIpx6YBdHQ5vk8C6fU9/RGdkRQVa
tbkU3ve0brJFPG/OlNUS5GORTwwhY/q5RN120vmAwBMIl+hkAodPSLkfbJR5Jfea
ULnIrlBfuSsctTCt8HkEw9xhibxZdzMLlbY3hPyb+2qSH/+7ME2RCyRTsZG9qM7Y
O4fxFb2IuQDxv0cN0TOmMvk8lHr1CYvqN/ZtVuapHBEyPXgwFQEbBTGE3y5DcirH
j5IzN20aoKBFL0nif+1hdq68Jmt6YI2pvy+Jd+XH7kWNNPtOXvTfv2zrUkXWZ4fD
fzyps5YezMOUuf2veK+fAVKrscbnRJFGE7ONw/Wz18dS6yBWgxBwwVUdF+Nz1V7S
UlWtGjyirEq7i8dlymjaqYriCVaN0vgOUDG6AxgPNcGDfJRRH68/vrdB0JGuuM80
XIwDQzUzPdI0imbzJlYHWy39OBqSe0b7kQ1gRPNtTWrLnQ64HuZ7O9SzQtavpV3Q
Ob67496sGRMLVuauJi/CI1XBrxNBfE+sINz45xkR0adExGoIo7tu3M4P7rCF79pJ
Mkuvv+QybH4XaEiqBqWOgbt89X2KhfV1nN1Yuz7SnAxVAAEItKb//L0t9XK6jO6R
vqJgVBUO0kPTI3UtvWud1oa2XM6WtVkQhFa0bXOLnH7X90Kh0Q4A7RhjVmGMbv9W
0jdSgez3ORzs1BhlW5AmAGCq+pUXvwvzsZBjv8+m9o0qBPj7O3SCF//LpA0o1Tzn
rAgSIpxoVSgNfTANPM3xq/WxDp49s7KfIE3XKD2Mgw1vvVOJkS2Kw92OZsG9LR32
wGBNvfWwTCOLQKOoa/FZ764izclQJDoDjluzJL7vkBU4HSS1m6F5JjTf2b4vzBDA
/nOwWOmmdL+QQbiPrp+dUXdjNJZ0oSEtlvM4/ksU1xSoEofYFqt89+hl8iP3vdcH
MBhslEMsnFP3bTRP89QhxSntjEas0WquKQg3Vl9cRMs9Q74Isog+hQXAp3OHrLN9
PB9cBX38/ilWZLTAIuULFozCnw7KJAt8K0AgzFwHP87MY4VcL4a8T3IShjNK25um
WxqledfL+fBNmak/71sv4oamcJ+Pkk8TthP7/w+O//4tUSb9yGlVkCNkN4gG4hso
pO3OTV2+FfMiskc9TZ3DTJdFYVe3LphE8izEAQQGO29D3984DgMqi3ot5I72+as4
cdphxu9wfygHl+k0SSG7/+aWNKUrx4uMV+f0B0katEkwBOQ7n3Bgx9zE3efIdwzj
FN0WUU+1DSHDnI/MXMW0CkHNGWQMzsM/kSAn86bJfFMKv4JGEV+JrBrff6Obn8T7
eZLRCk4F4R12VXN7Qkv7Y3t2+fmzyU6uu84iRcRXi9zWqSA4IwczmArx8YJd+Iy5
UaWbrvPv90cCGj1ZBm0eg/VQq+u8hLpeHy+FTvQO7g+dD4TuZnVv4W3gKuvedt8y
dNrH7pvhq5Qy+kgxxyqtb5D1vRU9aw3HpoSg9I1CmX3PoV0orwrKvRV8G8kfPCHc
akdV0LRzPZLu7dL4FcalVq1u5lEhnyT+/3fhwXzEyZNFGyaD4PK1RG2YedyuSrRF
0XZdbEXEBNmZjAX6ojkklgxKRWfABPd6HboFeRO3uxvsrIxOOWEVvy7cT/sKwOVK
+t3CLlq+P08YRkIw+g4/MxcyPOX+k4Hko6gZf17hAV5h5Z+fk1I5v0PVFkTpANTo
Vn5wJ3uyJclCwx5d33axyC75o3DbO0eitQymvsru8Bf6QPNstcBZpeTp/T7iE4Vy
GtS9cC8/GgoUXNSJRNBf/zrGqlPQYVJ1g4mHbfW0oJcOv9wVyV0Qlg1G7K82HvTC
7PZM3gL+0H1p0Rt6j4/wY/9laoU8/fdwPd7yenkBR/8jw7E2s+0VAg1C2r6YvOIi
L9AzA50yRdo7QTOokdARj9S1AgqJ9000tPbo7YQNVNoyq4Jw+LhPUgGnTThwZEGJ
0oxduGw7H2ouebwavdeO+b2WOGHKPHWTz+8tZkQBXn4qrJ72zBO0e7Ns7gphEWE5
PNdWvjdSOgHHVzQzf+B3K4RKiY5CfDdjfyOn/cK3rlrT0mpfAliGVU4AEZQFRZwL
mwJWW2LannKgOVkIZZJZqjVpLIcAl6v5bS4889gvoiKWO38iH/8gUxD8fG9z5ZrD
CVpDvI8EcYzn4QgGfiR36AdmPDNhS7bE0zOR0X0ErTGhMsp95c8oPc5MKE9coQCu
jsA1npMV5YfJ98bXV3fcfGqT97vArr6R9pRB6ilxfBCffyCCxxGogTXrw/SlYb0Y
2Uwp2aOtJLIccCexHBNN3eq/5acfev39ciUuh2g8bpE4jRv/007yIubkHdhQSgfc
tIYagXUww2nl4oknplXdX7LeAj5HEkulyi3NMC8SrTVHtVJc60rfE1/HHKSpemTm
W4oSGQbIYrVrp9PnuPf74GHhvBw4izAR+r95lsmZlUyCfKFNQSGXxu4GDLD8CrM0
Bps9mp5EikvGpFKvzq+MVGyOnE1qaaRaHXAvHzXmjrieQNvw26PzmE2VtHf08HVM
XrOogWBFT+oYjUJAkRv1qD9O+wmQWqIZ/Xs2w38fMg8ZwUrQzyQxRfsmTIrCiWYH
DvryRFlV6oAauuMaYPwZAUXQVvY5wbJFOI9trTxc54bMTVTfEOS1w9YGyiE3ajOi
57AD7fpOiqy9R/0I91lpLUQT8om1Y/YLDVgldGvNKx8MG205N7zV7gD4qFCrvDMR
sesGHLb8/cB07w9xaeqwcFM76B6M/MIZvbjfkbcZDwwMat4N3D5kzI0lN9ueG8ft
5KHR/OOQfZsRLce4EjcdUjdOnjot7o949FlhxC9o2eJWJcGPre5blUY2G2X8cp62
Y1rrrrR+QqzAz4oDyTDd7ZbP3sK+KJmUlPNBsRRHn7WKf69UqkvxQOYYOyfYFQT+
kwh5XWPFnHhnJlfSkJIlKjCpEduDn0hiymZmHFBlO5xsrFmLAvXjWxTF0CiNd/H3
m+V5Hw2dyrXCmFN2j01aSk/DqyqcXj+0R29XLxmbpuHoPSQnxAYiRqLp/k9aHIy7
5un4mYbexektG4Wbi68cvoCJHP7vU4uC15kojuBXalln3xc3/sxsmm++k4tcGao6
y2eb/UoAWP6XSFzaSZY1Fxed7x2IEJ6i1cfHTS2U7LuSZz477BZKGwagI1gOYXjj
IoayvD5Z6sVAiE2FSjUB9MIwqDP/6L1LP0L83Y5/yAa8+cN56bsDKoAswcBAKfAm
IkpbF61aACyl9J0RZGpyRU5SNrALNyBfuJKJnbTIIVlop5S4sXKyK00tQKQywGa2
H6MeyzvOGcphft+nSER/C+iEWbOhfxYe9W0urqdRcnrzVqb/NjOnpltM/qDLM3X2
3ssHtBRhvL28VNhe7l/6n38cZLs77cFkCGntHGpVxTkafyj0pQFVl/pNlmD9u0Gs
9GOYkzGVVTepHyZ9Lt+2szj0isnSo6A5f3HAjLcRWC2I4AX6Fh+pX7tp/jU4qH3n
2hB398xSeoGMzlgDSfO3R3mvTZX5vjdizk6WwOCQTd15gFmcSJsp1/9pXjcmFJBM
4OD9VR4JhmAH3NGqmfPds1dI0F9L2nZhJuUxSRBTK9WHpkWMXSkviOkq7dHkywRh
tGXBgO6MfI0pnFaSPmZv/BYzp3xdT/McRA+/NcGTTObTa59vMFG2aCM5y9DdKwNP
wD0b7iABazL3WQ+PgG4yY1yIdWSNtL3th/1ABC5HM0FeW8Fa3cyefqneQerajalj
wACxp+AiPgLUAVJeiuT44Q7IEp9GJP/A08KvGbivMY6SUVYsyX3zZwOLUdPozKVM
rTGuru2dUxpLYDVta7lXQyT5yfgTZQtdTIQ0DHh9k3Ijyj1O8U2HcU/hEoI57WkM
CgvEHO4jUF2zPmB90MOiq3q73OgxjcW5W3LzOHH/jQgnipJEavutPy+nWQz447St
JuwUmrmksRNIZe+UeieFaxT5r/uwfR3AoNZjbMx+91rJihOW8pp9TFZ2mfuVSxlX
pIq/q87wg4rvHWJkTqb6b3LXCs+n1SkQMmes3p6czcdaKDWZNZn4hG3eMP2yzmQI
R5VZx05jJ/lHlQ8rMtR4M5KbK4yXoWtW1DJaX/CvYelZ+/gCK30ck5Kf3peNtH5y
ztjGVg6Us8McHi+Q/rKFsZ7jyv7bmd1ex7lPbjz+yHYxrMAwStL70j/Q6XYl6QyH
y+1Y9ZHkwfqWWfqfH96XLYVykN7bg7SrqCMYRd9WsjJaA/KbvKqRmtuZHwjZBAOA
vYVBAJcdwr2XNZnPDt/qd2ZrU8VbSlA7rFxPQpCYKsPnJtjetYIj9Y4F/IYEC2Fu
pyFeAUVk18T1q9MMwpUpIdscgBaCpec0NopLEyJtMb1/YzzGp9I5FQhbw8fGLqtU
ih29rfIaRP9l5JUBhq7gx7rc7LW9dGlSR4p9NJQ9zHt5DuCWTBTMXDhW3527jFI2
8wszxDvS6PfCBR0d0uhSHEGGI48Ag4Bg2RGqjSjN2iLY8lD3xMPRJ/30tM3C5Qii
KSsLeXr5clsxDiUMbKiQ1pfpA0ZA77ygF1y3uoTxOGVtvX+WTDqtZsd5Zm9HYPTc
rHsXNuD/LU8gEgTX8lBycd7K61Rp/pg+EwzJVGE4ySQt7VxoBq3lSj1jLsDs0wV8
6FzoBe51TK0LYNVNkKxnW9HfT/xA9Aq0yim6o3NkkDm9fdU1j0AhjHtTpmtP40Gb
HL1wIKi4gy9mf4y3JlMxK01DNlEm2Og1xQ97bimsonmRuRbcUMZ8Q4LMVkqb5Oaz
0g/evQb9IzvS/2089VGRqkETZ8J19rmNaMJPGmtJsZtN5mWDbkN6t8T0cFN+yM7R
QzwDlz9KSpgNjLWfCHnZseHlnVLV3IjyHbFaPUONq1c6jZsUnts0Ynnzf/iGxAUH
aiihpjC/mBrDtkHe5GsAm81AFRo/fZFL99fh9gHffQXSj7P1wchCqZNEqa4cC6WR
4c4ajyDySIp987bvYo3IkYMkNefZy+KyxDi7T3L8btJp7m3rFEiYxK108JBpTZeo
ehi8CZM5h+nY17gvEecyPopiXf/dFub8ARXl/v4kjhCnMZl4ifoMdDJUCAfBjNNd
bO8eN5wq5+u1JVPG9ho+UCephnKB1puGfu6BlkLd497dvFD1Hp82Ng6brR2WTww6
ONzvczpBKA/TimcRYpbkJQGb8SodCvlnqYgbO61ta5I0KOxHak1Ccq62NUDh43w6
BBSo1zMx2OeIDmIcqSZ3w2jooIJv3JA2OKN7Z9/H9hiKMmSkMnvX3fCWgV6rCPrD
KThYT7o+ByiWLhDjpcucoLOhtGaA9FRIOyGaj45g2OPPqUkL0kRcotgGIreW9e3O
Y0xuKTqBBTIlT03/xObcd6DLlHhs9KuSbC1qjkp16iuEqVnny4Mvdw9bISfqMMtt
P2x6EnM/fn8bRP6DmSvo3Nv5j0HmtPkDUUtEODpeVDEFt7KM51FWXkVMtO4vnd86
IGVavRTneWJrJrxFDmHo0MGPpk3MJuBIuKC+yhbnHmcjB17CI18TDszGBFdcaZ7W
jVHuoruujCA86RIOf76ZNP2WchtTjnBeK9TfnpAv9oMdKh7b9VYEf6dM2NkMj1Rd
A8f+w0KbYLa9In9zLf1ngHupx29EtuMnSgg1MXnuKgv5v6lIxWmAdaHsf8yr/0qe
INQElKOEoz58wEj+3NfJtcm9p/BO4bRSJNTQ9JwzGHA61iHr3bZVQGIUo8idKqF3
0Ust411Ic3+2U6CTmJ2Vw7SXlWY/uyWeiYGld3cqC5ig+7R0XSRWoNPspSERkmQx
5mxGcZEST1zE/TQQq/DnWXpAE3qs5CZchQQ5IgB04rhqyvPRxRESoY4OpHFpc5uW
RCTog7V2uevB215rDCq7M9XpCHuFqm2lqOPMdjikNPGJcoVxGo9SRGL85XoJ9Eb/
hI6x6WEADWnoZJrNlBuFW3ucO2Slu3vPEV97ND+KYbpXk2T80VPBXVKUVDcfqxUh
6Gcelk5Gqt/l2PeYJt3r1/jWByjRmt/od3wUvXEBNRhezSulnIgJknXlmQFV4vDS
L0AZnvNXxOZM+E5EeAuJjya2gnFx3Csggk6XHJUq9e14rbwAJF0uGAFcXDcVIgwG
BiwQ+OfcKFRQZSMGy0xyFl2W2yj2BGdQEiQNIdB38VmRiXZ9biimQcC4oo1ZlZUb
aKfel7dB2na9eRlLdBoMEn0wKPnfLxtjpEP34aDeEQOanpezAxs0fvtYr8UD5QtN
bPJ3q2k9gicrUbiNB8rg8bgpcS216/8+8bZc/IW+f8hi1ZmVSubodbQ4Yp/ZCpX4
I5j4wGYkgslvtdDPIzgY3G0R79t+AlYtAqFH2yPntLfPQ3p7ZcuOtvWB5fRKxwHK
NZrLudDoqkLIfbNqveBWSR49adHbgzVCz8Iw3PjVaBWsXN0lEqIlckx1NqVHBG0f
3drVyvyrOj67ok9j8l4KwerZHolYIPBFeEwW5pN//QvVALcERDIrWDCZPOY3Rpom
DuBLTC7yXuKF81GXgKvsREeHmwO3b4WYSnsYbAMKPGCrlvlY6pdJGg1tm6gD6cHu
wy/y9x8IBNFZbHw5GdJq/IrzfAGiR5lvlCqz1/ZTsDqAUaefMIXLyqD0DM+czZjx
YstfQgY8RgVQD0dSG5cITDbL08rQWBDenIIC7u3L0TPs+ZNDD8lRo3y4kaMBArfJ
yPs3gS9udUKbP4w4mJgkuISkzwwNF8oSE4C/LQ9wzFVDIUIhMsHLEX+Ks354WQUb
u0KOYr/Muw0ZZA17gVln+oyyEydv8F5EpgsnZ0wnYapZzqP6cS/eKCGjZCukr3oB
mqomN45AzQzOtfgDPEaZPalUBt6Uxfjjc5J2A3rMAPvIQZCa/B0o0TWeL4wxRLgf
8sRqQMHHjLe8m3ZvCzAXtSMv+RAmVddwlKWUVu5v1yKzritKNGeWOrZyF+h5bVVb
6mo9Lp0ZSDKpw/LmuQ4r8rjVDNZzKdS7nSw4KVs/ejluaVUBMOIxhDIEKkuvKgDH
uQsNYePx98XePxsTE3OFC7lI4JqYk3NZOhbpd2euVWd/E4KO4pY8qEYdHYvGYOBo
HuJJRmCLhcQxGcDNNKOpCCu21WTUY4VJmfYpxs4JSGhIJnZD54RrtBSIGaVRrF9H
PjACGZNk42x1NXhIpkY2tUOFaDBN+3l66bF2U9AbADaaz08iGZmWqVRuFmH0mF0h
r+ZvdsNCiC3DprJQQ12j9BNQd5gPpiSadYsTOsEbDC02Hm3l4YOhGS+JfLgIuz2c
2079Av/4geBS1sf+Q6jVKOOFpmhsbZU+njrxp2PMU7BLWeW7b0f1srCXZau7Fybe
Hh5to6w7yINO6aHFOEL1DGxzETApbvEJN/F9/HZT+QTn4gxQ8BcNUfpt/RwIBrSp
LevcEuTjTMEoPeQ326XOn4O3Rdc2bRSHfjAXScJYuKNpJj3wTxfAfWxaZ4JXD5bz
mtfkBbRVd7sDowVahdA2yraxDujzPwPIdoC63T1m2+XI7spH+hy4ROfG6hXicmie
V+FUP3PMw5U9qVPDpfVkutueAfa9Zqza/7K/KyubDSpyPNzyUOszscRd7iQBeclO
EfJztCAWxerGRRDI1LLCwhNAK7DV4F1LJde6ipuHGG8R7BCYuOn1X2j1Sb37vxTh
/iBs2S4ZyP5Qn5bZXyh0wt9JhN9NKLo7IAQkGeBKP+rVJUsFAqqVKhsyu+lISY7G
ks5I4dayoJ2tK2OGkLJmBj1ZKOlZieVeXCZwb9ffZ7NYcZ/TXlM8HXXCvNzs9dif
vYZDJ1cspPRPva/zkyUu3XT99WfxBfLhg4GxQxMlK0tL3CNXS0VlyaA5juWojPyR
amctrLPb9J3KroXjE3s+/TTvsZJdvqMR0/FV6ogyXqjU9KMyT0N2FrQowfQn+WUY
Q0ki8RQX/MTJAe+Ij8OIYo59ADHzqqw0gYQOyKJenF9yPBy+1yeIWBbTboOeoZMV
lvQhcG2O43WhSI6ePwQ6uKssKryIcPZL5UtS+/qDzMQo3QpbvhZOjj+pdsDhrOFF
94t+rJ5oEZhjbqHIJoHcg3mL7t/Q2HuOKXxm4JihFDmge394CutaOeTfQH2TD4O5
Z9Y4QgazV9VMWAKOG8wHZArSLUOFxjgTxkSkbUW6peLTnPH86wK2OzsuELhB0bUn
2y3kjyN6lVFzckgQU2qm2SZjmH8/7mTjqEp+WLoVn3kBtrKsTNCJBJVqj61VZyHP
nKrCRFItDBeqL4PiUX96JumsTAnyNo6wm5+01imwQ1VZb0kmdMx9E99aWwivEiXH
kld83lnHSzto1cwGGVQb2/8JyToGCFvHb/jlW1vrzUFK01Fbqz2QakQOI4zdgO9A
xePk1tqd5Fw5Z/H/o4BQXpeNMLMLh4i915xiHl2jGATUaO14Hl46ZYG1UWl56k8L
ctxkE78F3KCpXJG3iruJ98JWciMcKraBJ6QflimLkzPpfbTaDHCu2tQHvqLgHnJi
q98RZkH9/EKOIOyuNHA1cn3sBmNJCDzBKJayinbMZdej9FCFG1v7PziQpkUpZdu5
Ms9HYabUwRBZreh7OJTNFUoy+Zy++uJJOSBCUV1aPTh1ma+GStic3wpnRomZwshi
Ic0cnaC9nkNV29bnjxtNndfKb2yOe00XLlCsH6jAqtchkoCDFYOprKKnQCGqS2xR
MsHj0sR2Z9W/Z4DHvjX+l/ut2G3vt1cgrOJApJuXLdK3oQOu5J7C6zv1apRC4cGC
N7Kjju3ayhRYimeuFlty9XQAw9+ShkBfEnjXI+wxtsMBYDfo+tFHH21SlgOb+ElF
2UFoniNV0uX4Rwgti6wjbU+yNOIcqeocuH3QJbJp3pDLuHvQgFWhZFG9iX+wr+jh
HeIXVcxa5rG1Z22lqf1Mq+jR2vUre1DmaBTDN7s47Z/hGZedc1PHSd5/Mg67+Xb8
3jukW2BZylzQqd1io+HW5s160FSjeUsvYxu7wQDpYPG1c6J2banQOX6dCCvEJS0O
/Pvmm4waqvArW/1qO2K7r5GoF80jmPXFI8uw2onNmbXiIwidGMAvvqZooSKa/5Dh
cydzcIqN1M6XVdciVi+bf5RRwKQTB2WvIS1qPZj7bNwI0hZtnIUiqXExH3LrE+Gz
IfbUsSXg2tQCw1NzKOzYW1GjVjoNYwuP2inobPV5mzbk+ofneVd2SXDvIu/SBmCq
5BCT7nl1Dw0XcXundBrGu3blP9Ds7mskaxGjsx1OqOmEtspF/iKb081CRj+gO076
SDBWQ1eTJ5PYvLXxe3ggfKnSAENa/D1gVnIngvLxs2DufvLcvCypjySxJh1j0T3C
wzx4OhDvwFQ/wAtLjMm2tPqsC3Fbt/pU46l4jzGZ5zaU/QUgmR6tDQyR7OqEPAPV
gPa6S5TAh5mx3+3oprjB+Ek2PfYARI396CoEV7bWI3bYL0n22Hqu1VzuQQtJ4Pc0
v57cRHrH0tff9C6540wj/NXNSdTW2kRsrWH7rcMiS8O2FNWkJ6ThkS/P8GSVaPxk
1xnaN2wRDmDp9HD5kgyk/SEBpwh1UjaHxuSbXPxQtnkQhs6kwu2D3Vl/r8wzqWDT
xvW0gCwuir5DENPrdgHWfNJmn6oLmeoirbPnvaCGIkLt6PM4Y3jgOVeYBTQM+fz6
3bfsya2/UsrrsG9XnNQYVuMlJ4pIYogN6KNNMwgUwsIu9VbdzNmnKrQImnKAsncC
GFyxuc41KHLFOLzMCOsFBFhq0Xw2N77N1OtR38iDdIYGfZf4INk4DEDqgXumU6RW
CTa54ssrRReMcyZdRz1yd5+n+f0joZvape///gtyUWM4bvKabwVVUnqNVxNQTRwL
nGJkFOgLfPh52Iq8w8iG5iBJZWjPURw2SBik6qLJe1Hfa0QBWnRTHGxUJue893Dr
45GFQCItjEsblTnCSHrGBU85LOEjV9r8nyVPl622igUTnmCbRb6BpkMDrTCDY7Q4
dtDRQ6cVMEHIu78F8jc6hM8ChSKwCm61QHNkRHfjN0X8Hel5cJMEBBDW+DtlZlXT
Erp9amqfYY4GpS6wtgqWAATPnr0Shab7HK9ZkeBmtSOC7jj61e5U9m3k3rWhz++Q
nmP6dNqTQ7ac/JIbRbNHl1jzYV/GWqiNo9aCWAJ4RIzm0omJrOlf5XFc6hd0/Szs
bgncGUcBNRuRiCzmlxnhtIDTzgmlko0MPXXq+ZE6ddG8cb/zz0m4kDPzX/DnY/w4
FEneKnt4PNRcmEJrlvi8/G5X9JFJauBllRUaMT0qq90m34lzEmDTQ4tHFyGXl7aQ
DsfSNaGrILXWIFCBZXGDQF4NPSyyLAzI6TWNRRt56yYnRGDkm9GB3Jt3yN7BTGj7
ggC6x/M3DJqSqAj+nKAXQrJTIotqan/03/tPkiecyGx0LxRnOV6vWWqvLzFefS+6
3VXtouEbdejP0sbLkJHAqugJvUxEq0VEQmZPgtQyziuBpign5nRxIv8RpmKkxHPN
eU5lBa1IIo4EomL6a0ZFpwvIfRwZse7CfkcdqSGTBqKfCVO0FOCqyb7pohzANNbo
47EXTheAfsWjpkU+G0v4FK9LSavRY0M2Y0rL/vmxPogVTtjKzmjUogay2Cv9BtnY
Yxa9c/LwRrLaQJLAcWsKYR75NO9GkoWGv7OY5XEOzjQitu+mCQspuHYyDsH+HhG6
cbG3B5QTboio8VZ/CV8etZd2WFglB9mns8UIye5j47A/zJA9LKz8CjvppkE0f4sQ
4RGAMdY9tL2WXaUynBCIhy44ZhncKjhVUho3kwvJGQEn+SY1PwYJdjr7jPP3ZEmM
wjl0Db9DufGjKXsFOu8a8pNfieCHPaavRpSfLUZzplQNbM2KL0zYiWo64psOCP3x
eGqg7t4a8F/hnGiTvUsrWtNEeFbD0qfV4jcL9q+ztme7JDDcAGmDJ+rrOebIMXqX
1LwLBnDyT5/txxQ9rz7u6kdajvTsGw+/iTY9EjVxQtwFsEPJiUhsKrss/igjnlPr
xCcDaXTHX6ueC1Eb3AsowpKO/a8aW0WpeTt8GoxjDO/MFz2RAmNE7luDgdjXp0Q+
184hgDb5zj8jEfEGcfcQpPG4C3itf2I0pV2SD1VQyPBz6dH73BRcLsmBz4xEFWxS
JNrRtAWqCrA/ycIKEPoSgLzxBHN2w682c0TcG1zNwHlZX6jF/o2uh3deEqDla2q7
Kesgt/r9qsKHvtEEO/6By9AsbDxyzrTyqh5yrR3oPnoM19EX4dag1j8kgnFSyp1S
yXFXRQSHkzOd9MnxQtRDsXpfEQSO7N16sxcPhRoCQuuYxhaEv/5nHRTkgMDwmdCi
8NIkPPt32uj62S7NAPiUsLeGrH93MrtAT3xduaPTGM+dTd0EHnp6YQqK8jigQBHf
+qoJrxSxL9kog50Fv9NqW1lwkP7NPfgqFXIOA+E4ulYkWy8J0CkNjreO6PnsJRQE
3RMUqTK4XUuJ9uudPqOG4pz8SE99/If2PxSXLkt3cphZ88mXiyCBOKqxBeSUIhfS
KvufWAmQdN0PH8w145RHiQtQRhTxtCZNI6WTl4k1YlD7EhrMvyzVUJ2yl2kkuUiV
sg1IywjyHqeeDUsbseQkOV/vcgmVgmPPTZD4uPm8vv3Vfr0LfM4xCFgrdLa8HUdk
FSwLfT9OSYYr+h68KxjGKRKjaROwRoa/cwhJ+/KkVPtMm5ocqXWMg8SJEf9/Uv1S
gJ68kkr5zUQe4/YTf+twZMGfvbnnpp5DDzs1HEO/bU1P3Z16s+cZ16KxEb69h+1R
R+TBx6npmJnJfqeqD530N9GmKYVVsfEEQZnSSSubiHK34Y7meSan5EW96i9hb8Jm
OQeDAXhsTX7dI0nhvaU93Oi1wiaOGwQ8VQY83YrS1mefGHKgZxpSXqHbjWV0M6VN
MbrKtZ+LIKGiWl57Lvw9kD3bCBs1CbHBslLyDaAEgT/D4PMuJRjYiaw/2Pto4vcc
sZvZjdACIy9lblsGLxKeJPru8NHkVHOTi4HrgRxZahuSCfWb2a0w31/0e9clNo82
IGtRPg4mdoAC7YH1XqPswY7GLoqTpnHbVYtOLJD+nJlFUI67wNZDSBAUqGLkqF6L
Vh8gXJR92qRpg+c+mnwHbDtyc7r3PRL5gUfhwyeTazhmTLsStQOK1yhYvK20WAZI
e25XtdSF8+9E0VPMEK0YCYScYA5vtaR0kf4+RLhSpvvJwl0m9uf8Ii2IHOl39rA3
gsdh3U/GNqEdAPGDBe0wnM7Bb0fFI+8uRjFCht8ee+6pm17jWEhjK25eUwuQF7m9
vQZgoNcYgGaEvhKqFlvA1bUjrk5oOABj4s0CYv1z+np8Y9714jgdtig1EaGyf1A3
ECUivl6H/F43Ufd73cdxcap0md9+f/Fwac+h+Qqa+58QdqblQ9cipy1H+8su6Mvh
MQ60dw+mGrj7bsnBpEUJecaulTjVbcNgKjXHw0bPjJ0WMpPzug2vWGP+5Mv2koMe
bwJ1vVLdqN3kYHqVFa4BEAH4KDpvGCDBTjCLnPt0xGSddxprEFCT+ZZN+GO4QUqY
mFoqZHlG95cwbNE9DZ1wDyVpFIGKP4u3Kd76hxTBUKEaCb1HrGhOhYUlQL2QXt+4
vrJ/ZDcItXFSePrxGrvy6KimA2p2tu6/ltZi+NJ06OtDf3a3QakIP90PuWqjjLi2
xYAV2WHFpKXzQ0rrhCcOZ80zeC/o4xKDs+KTvKwVOsGTPKnkGCwa9deCS4y+/mkx
hNTqEunnztbKoINvQqr5QlVOcomkZsuuE/HdsL9ERDugaHyEPIAiaXn9V6TwbY46
KiGVXnuSBmM/yvv1kmGKNfgvL2YbhJTw4T1Pkv/Py2ijzExJDS5AyIMV6mkwRLF4
LeohmPGX3bQILIzA27CxLgWYphqun+lgtMfBTqDveEn4S76CjpW9lPmJ9rjMM9Ot
VhOLBnZp+ptCykDjXCFn+W9IvLkKxz4lk7baf0WcDj2VIOvYlqsyQf4efJSYXHmq
9tY8VaK43YxhkdsRSv5jC5FZCdcFVXSFXr7yFCvWz9QA3i6HEk56DchxrfjKZM/y
CAiX6gJQCppilZjTALnlPCYWmREiwx7Q4UOhJqoC8JC3yTKkAo2JzS9ynMYkWEcl
JXGHaaeqwz5J2kFjKywvBoOx+zYRlh7Naw84nT1j3svQP1YdrohuVA6gWvCFlCiV
ON0Y5/0ajDIhuzesaEgjqWsfLKdaNExv1j009tN2p2mXEb2ud9+1ovBwiIIQC9Py
D96VgHyprIyM+xGDzKqAHl8CI2KR9OVQkqUkMwO7VZ0mZbZPsWZ1W8VNwx0FDF22
zMQYw3jduiipOLLMmdrPMbmipRT5JneTIDjBy373ZiMGbXCQQN8k++anpptEvgZk
67k++E9aOBSEnT3/pbVdTFbBL7ghi+ywgIjOgJrXGtWKeczeGEpBmFpSLQZn0CRv
+R7p73Aj0rxLR0b/A3wtkg8z57gM7txG/LmboWnTnh1KcFbCDQycnIgfXTIhadez
XPa4ZWHZY6kBzuu3/x4y6aBqKpvYHMHsOzqbwHqYo3GkFwHxwXeSJc3O6KQuLZHk
2Ud7u4PUTGarqs5Kt8anECh4k+1XZqyz/Qci8K9tE4r7zMntHvgZvxqk6vyKXt3i
klFblHsNDlW+ia2/NGeumHoiDKqh0fHdfpWjwYV0pffFBDZb3YGAu2QWrzsqdM8w
x5N/xis8a0vZ9636tAnoD7J47oEKQiPs9ixfasZ4ZO1WE7DM1H97pLJh4ynAnvCK
U6KF9sl91gcbp5DCIpkHDMfV/BByuVqyyhkuElc2+Hj6iGsm0yq0qF6xZqc9dw3Q
+BwKzvFRf8AQ40wj8vM/ru3WwihAkHnj76DDn+NCk+agMsDEncEYkYlaHZG8A4sy
GUlli/BHRCaLolMVBQDHgWnPnD/wypFIPHRHx/TMUDuPIfeu7TBi6wotYHtG9f7y
dRT2FwtvKPdRhhvtpAyPgP6ULjyHVgRWCxQBK0h6q8EwzFeotZ3qoPM3ig2VZUZY
Qj/wQbPdKKOaEYkjluqXn/JgMy/UtgohrQ1wcZz+Xcpv1L7nVEH36kZ/i6kKJAcP
o+c7DmjFZ07S/F5cLNj0Az7w+I3XdfvQSpeyQp/b3/CdRw3RqWkiTY7wQ3NieCs+
Y/DDwhW+DlKoK9vy5sYKgntjm6ILha926dLjkXWF3BK63QiuBdkgGc61BIhZRvnZ
snF5tpscbOKrCB4XePX9D/pyjTQZJQzN7AevBVxob1cYSZdB6xi2wdV1IqGlRKg+
8Ie0GO4qr5zh+GI7jEwXn3wxcosIghS9ZykziNG9DZUBj9UPGrwHtXH11yxWagHd
L6/0s3fBZITihV/bKkuwKZod4uk7ElKvkr+TwPpjrWVxo6X07MMqer3XNllEIb+g
IE7O7VP64X8FcszngLLyOkSRL2DjwB1jtrLs4uuRWUTUbvaF+k4ndFUSu42GpD6H
qV4wlZwBFCMbFkSR2yhMA9cb4mADEmvtTrRqMtYRVHfcKN6wrd37ca4WprMt8Uv8
bYyuNcKXFslsAA+z7e9BJ2ctWqrFV4Em5KgajGHjzPdmGYAupJtDzDCX/B2ZJkdm
4ie6bka13rlNGlaW7LfQa3y/UNHNtbGd4q7F80FckeVvwNk5PcjV/taoxMQJb1MD
6ERibq4D8w/+jLLxgcfmNVlHnB7zOmMByBJAgMW9Pzy/C66KZ+fgrLK5B1JkFQs/
SHPxcOlF415YNUbVx5F+pDWzzdmYfBg2RhS4crH/VVf3Fl/5b/POFMiCStzJ4oxU
TFnnmBs1AQOnFfoTP91J3aC+0WUk7oER4QVLB/BTr5HEdp6stwSdaf4gGSlqzBY7
zR6Wka3CWa+fh37atUkivii2vhm0DUaCwsVuA8h7RsQxmx/iqXHisHCAzKbfWHJm
riggwJqGQcZLPS1PHKYuVyMtZsEGEutxxyOqt4OXXfUYi8Rde86asfc9u2yIA1Le
G5qyli1w2WWUhB/W80mzsDum7ifBZOJmZMIlVJrb94qzgY31CmAJ2KAsgi17ZBFQ
FH3DLX9BIzMpmQVVEFdbZKwzor6iqoFNJi7nLF4Ys3C40zKFRg34dLtDFgn3eODb
4NL181dm0ELqXQtHlxYZXcpSuWfx6E5Qlidv+0BXU6HchI2TMNkZGRJABdytx2kb
rY10a6cUR294ptwYL0h/p1mUl4rRf+C8hyJ8ZzLI98LHDiyaMZpTEz99HKxPFJZm
+BBxDuFDParNm7dorqOgO54wizZ0039sjmNGaF+l3EiSl1bUsLsDWOolRqx8ENSu
cSEkWJqShD0rz6BnrqCcuGdCtofpzsJ8Z/XQf+sjO9JPtoVd5edOBm90cv2LWLdE
I5OofUtkLEQC+F2EhSB1zLi3haIyww7NYG333xlaaQPgeRsGbCqjdVGZfIH9+CGF
+B2qjCqZpHeaMTwX7KsveiogkJ4xCtWqo/U5rrgAGSh7g7kNSH6rl/31c3hsSIdR
Umw98s8zvriYj9wcX32XSzdHU0pWHELrk0a/Ks4ewEiC8+slvyrb3GioDVnUJmkp
a1fJto8++zmwi9gA65q5vQwlq/sE6nEQbO9XjGXpyLbUwSvtwWtsHEsYGO6VLX/+
wu6YhxzmnjSUdBcS30XhlkbEj7XDvQ3runwMjioNzanli91Ato1hZMjIS6lYB5/u
jKINmkcRubSDtVO1tuUlv7Qa2u0C9EXA0lzE8EARCNoxPdwPp74WjVmz1R852yRh
foFXZGuRdoFlWfn8T2s8yUYyNJqBgHKK55YTIUI4POlRA4sbQWJMnQU74rLWBLc/
7QKbKfeqFQbpylIcVZFYlZPC5bVG8nUuK7xq2EukA5+cOSLLdcqIAZyizMQA8VXq
6XD2wL3dRWIKhgpuZgXHL82psbGmJYVunCsgRGEPhWRQvUCyVQJmIBin7Vlw/JZf
sxVypjy9rhQslg6JXd0wapXjvPAX3EbKKUdU22zKUhCcAZii7dUKbSxC/bY5R2pk
4KHe5Jjw5S5qRaDcghCp++zXfAeSx8NcYVSCXLcf7S1gXMFJ3Pc05LR4k6vqsObW
DB/VLjAQdvhlBS8tsvdCllzQBteOsenvtQnj/ZZLpNdR7AYM6pky3v7L2gU3TspL
f+o7r+2pPvCn48fCaRasZZkIJ0rdbAeV6moapyBwVLpiEcCJkx/DKzNEm2LuIhHc
F7/LKMR7rXI7yoUe/9JslLm2djASGD7eEeHQCousEOd0QBU8fgOmJ1ZO7pLuvQ+S
TgeTTDAjkv5vyNewzs92CoOSmMyHVfAWZaVGCDqxPFbRJMui7qFuaYmNKUkibz8G
0yFGDoCVcBOqH6wPHxxPx0SdJUU5dRRngurwxfQMBiLYhoXn+XwZyGx/Nk9ewwrn
t1zMO9qXoMFmqsrZqHg8riYqZ2cSz7XEBkK2mwlrFXGLj00feGkpMRjxBKF+qkh0
8NUKZrALwy9QRJBlfh6+BDNaYhxWcxWHRkxEXEtyuq9A3vd4HZu8Gqz4s+dcceE/
r77uzgxdYWBKAjtmsI6vAuGLRc2TgJYmJeg3n4vcXwfRley+qu2f9gRhLW2Fuy0W
At2LaJgf++pB9u0bLL7FEPaxPWXG2qbKjhyEroEHSk6iiDrXvbdFUVmfOekqm70J
ZePCpgQCjZyHoP+PYaCRhPClN9a2TD8jfOxeINMgWUjk0gVreCwgrjJbxEWBKJcP
WTo/ALmFJNCfBgoBfOgzAOkLylSL36+A00qG14Bb6xhkYW3y8IxcOdipIoluWnAe
x6kfYc6fjTSboiLL8YH365GofZpvwnXMWZWkMaENdPGitHmRlTXiX6H+lN1MEB8W
5G75ckN9mA64Z1usLqFVZ6ouGx3Kob3n9v5+Y7zoOeYx/nYspN85d+ix/RFq4/c3
fp/aci3KYUgtHr78dKSusHMhmc4D9dlvJ7ZqjBsbzrM9aoeoZz5r/4m2SDeR9PDc
a2MpBEB2xBi6dYe2jAi1BQXqNYhd4hM2QAVkKjh4uisqgxjsNiemcJLIcOtYPdik
6c0wwpE3kpVx9rXb6wzHBYOBG8S6ooR9qMaDG6FDoRYRVszYU4xDLbdUNC/n0mDn
rjz8xzFuPN/VgJ+Ry1Jqv9qDrGf1sDaiMALe84pleemangxeIbFD2WJMqSgv0dVc
83rcC0smNaUglolipCJ4XkFdF/vOvTgRzlzP33OzoiOInQ6c8p0grUTQxY9ROYVp
xOzTShbd7h2DGiNqzRC7J8mFVIy68/JWmWLIywCP8J98vf3vcwBbB+iFYeaMaL60
0b/HqYbKrEbU+WSvhk3x2XVFbba5b1zakrVuYz9KO8P6FXmui32SRsRk3izAW8ME
XSl0wIb/hZnC5b+tr3CvF4SSMWfhMXApIrmHS+67epZmTMzb7mcDjS/xDDmY3mBh
QhbabsE9ipFhNUTdiWAzQFMCYOWPTHnJ0euIutCkjs+Vp1TxnYTq0y+Qg2D0K+e8
YIqmdZmkIp044rVjvzpMSkIcSKTsDYKzh1ocuc2i+9Zif5lwSRO/yYGIB8KTSNgn
BDTtSj6cNHbAYp9VuM5iG1Q1bsmor/HOXBMJB0zXzZGLOtoivmr2J73AUwkqr5RG
7MFYUWwcamzKWihoheVr1evbuKbKZ27KXMpuiG5TI3KSOqRDZS18PRqrCnyzuYkq
ItE3QJmyfNc1XSkGTHX9bdvgG+ERiJIk9t37OSIo4VTuP96si0ynM2mGCLk6zwze
jY3JCenOj4xaOETbnBLtIkZvDk+n3giI3v2jcg9OdDAl5khQQQFSEiAY+Di7FgLb
3h/OohiM57NTMQGQX3PG1QWNqvv9Ci0JB0LGFEz2+D1uC/VlSV0WzWd+FFhW1wi0
fxBKqjhpY3PQaaTUiaA3oQePujt//HHvJSzq0Qcnhb54TVpjHuPgpCWCFSFfMGxx
k/XMfZfL33oM1tHx7p1C+om15KN3SBnPQqW4T+eWr/efQ3JxXs//iXYEHWSpExAo
lgVfjoKDYaKCcgo0nCUnepD63dzyubkmkk0mUBAZCKAqtogXNeKteioakRHwLvd6
aZ+7asq65+jhs9rQHp1t2wAC7aAnctmtXICHAZwuwxiG7NFEPgYruxl4vcUvdvX0
yE1QzT53aMyy8wCCWYIFto9Yei8XB9U5KXGNYMGs8SW2v3MUXTEz/Yzm1suuxc6w
l/s7RKbLc4MgVUKHx/mDProsMW/Ms0nEP3tJ6KodwENFQdiH3/7CwM38V9FYkw29
i21wwkJtQN2NewIn+XNqGJtsV0yMBhCL/Xkl9stJm3mx6wp0YNOBKqN5yKptJ+VZ
s74Oe9RBzGHCKsmcl7HqcPqljNLt4lMZrheJBnP0Znaa53/fKA5zLObE6O6JHDLu
Pn2Nb7E7hcxGfuvsoE7JgbXxZsVswHD4Eua8F0U1Kg2k94meQ/w4ot3FQDWnyUC6
SntE9M0TdWr5K59T4fviUm0eD4cC+2FvFpvhXfulGXCoGWx7ud6Ljq8r5fmZjk2W
X0R5RUDmkb6nS8R073HPeEsQM0nv21XY+e4YZw8C43Mss/A+1rUGuNOTaTnTPXLM
B+5587L660gOKycBlBefSmdxOQCM6Yson+5aFO/5bV7RIvZmnkWy7M6bD8CLyQiX
FLP599oM9oBPLCqGYBX4PiDdJEoYb/0iAxHcmdf5lyNAOzhLt9peL281Ri6bKGc8
YOSNA1L0ub7jU5VFO98DyzlB4ILgSOjGXdMFy1l7rnBMrkx9Z+ctglqu/s1ad+i8
O4QUL82zGMplzxR+z/5uoirRHbCNdTC3wb8GMpjkjt2B53nGcWmKb6VirAUGTeyP
Yv3bdp9SKdfPcZK0aaH/7yu//6xs5a0r19dXIjaeeMVLVKtnnsQAM1/BoWMmWSse
ajYNJj491pDyTFWmXH3AuqX/wMD8mhGLVCPngT3wKmMv6KeCHchI918zPvUKpxPr
7ibgyE2IVewZJt/VfYJO4o9J4cpzyePo2nJJC8nIiDM4gOtv62ATjd1JsfQ3D9kU
yJA2Ajg3pAScPFaM4HQ2NbuaJXENV52ZK1bWPbIDTjNvrw8TKhkAlfZGyGGt1IRE
Blj8fGRy8hKf563zZ3JvpHnMyTb9T9+j3C3oUnK9/agbfYd0z/HXIlLOzZfzih8z
IxOvsA3E3b5Cnhm+PfvgDzLoySxemfhu/+Rs39VZy+Yc1a/95edQGvXdUyPjMKSP
QPFWZiEgzDCgZYW4tmnyQa1ewKW00oKEqJ3eW8Ri9tbB9o4E8S3B8qmxo2N20zUV
3/ehEbuMTOzdK4Stkz3i6w55UjdTbh7HYTY78t+IoU1SpSleKMLKsusQ5dNzKgjH
J9tQ/AucAT12iipv79Dqgzw7Ii05LhlIH+4HHC7nJvs7iUidoWa3c9yjqjFC2eE9
O71vsTJ2Po+LtoBnchqOzgV4BDHnoAInqSWpZItAcR9S1QeaNyzN9cFvLJb815cF
hh9oEMMOUou//M7wcixHcd+5ZtN86Ry0117lYWrTifs94dTTBt8JzUsFwkt4HHgl
mLLGLwmgGsHdNV7iLuFo2U55cnfkjQns1o4zT31W2LoyuUD2k0wET/RIAATYSTR2
Jg9HIv0y+A6KIfqRqheysv/7exXwIuLp5yxUFRzH6+4U/bHeu6X0MKJPO+e5G3DJ
VCUPtj5sWwu4DYi/iTqLqKa1ae2jFLxsjnJV0Xe6F2Ryzw2u1hEKdRk1+prTy/C2
DYz1st48kuxh4755i/YlbT0HNWjzuSx6/Q5l7NPwhFGc67cbslvvWo++G2JavHr2
2E0S7f/OYkyruHQ2abRqiOiDiNq30wAYo0FYj8xYOmfu/CB5fpq/Dl7DhJtCTBIh
+cB0QSxlv8KgL08vgze6uwu1EpbXAfzch/8v5AWqBW7zU5mBSmso27k5R6AjPuO3
+woPUzU1mxHyCJsxC+6Uawi5NLKL04DrJHVu1fJruWz2upZe/eaMSfjCOxodz0fK
iWeUCUO7ENW45w5kTRfdH6Jx/I2gMiN4MQpbAthsATunbHsg5yGqwuD8URXiHzSE
V/0cdvqfrFjBaH9PGst3QHptRoo5OmoKFASMplMKc4JyQBeSjMH12u68iJDXoGnA
fI/0oqiS2490qcuat7XjqlyFxewWLyB+fDhYZYJLaZZ0IbG5Y1SPNn9y/IUdcIoB
Y8dU4h2HUx16wAuH++Qf+ZO6em2K8ZkEMccUjL2Okgbem0yJltKcZmFoMaJXXtRO
aZCGMSMfTcKYjlrbtCYTMTZzyaK8mkMLcfHkhGwoxFhmxiD9/brs1MOzLzloj7Gl
UyjC+vboG38JRNLTDfYlh4XSfA8zKCorVd6GAs5mvbOStWj1sykciVkVqc9fhOa+
55EWiNwqHVsz6/8U+LmK8pFI47JIH+1quOPYtAWEiRs2hJNBBFdPb9uIZ99atk/w
eN3Y6Iu9JZlQmfjdRNWNVIcNM7/cYkKoMfde+stwB/yXGPvV/3JwpyOoaeqFY0DZ
a62OLGCjHY1S/kojC6VhJ4ovjX/peg0jsfIXqhtHPVegVX0hvwpec1Y3zE3q1No4
IPZFXXLtIg2q7kQN9iHFGbNJrOXadzDyKXcWyjFczM28oX4mUdWUkJqNeY2GudOR
VcbKaTrQDyiolkmAGOmg3UfKMvho8Fjrq4zclfbjUttnE4CErBJh/VIpITttmfGx
DhsdLW4jUmQaDaBYZCHuzvWriGGeJSR1hX43VZqlf/b9+9AWg5phJFYbMaR3Rzca
2UI8deXbgTEslvWKk1AR++Hz7j2aVEaDIYzGG5+dvtHEzBr45I5x0Mn0nv4HuF8U
HTimOYsqShCYckv5oICdPPp4st8StZvlSglhnwmD2cRBoDCkuZAENSt2akxa0ETy
/+jabfpWrM49p8kIFpVu+R8yw+qfaDAIPI1ZssdGcOzyNotiPssC5gtGvi4UiYZ6
sRg92KA0OOKZYbY1XFbGvVOhAn1KXTXlkRLiJzQhbcYNDgOqoA1cTwqDzVci8HGI
ZWMbJctIfHzGKZP7cFCWx7xWQU6KYvUIBi0e4pUkuS4JlAJbZPfuFKQ058ne1v4V
DWcWoOIoD4pVWNJ9wGfANU9VuPh1AshsYJE14tLVsKKBBh0St5wmcfM9CKxIE9Qq
uh/ksuHTGjzxwv+PN+L6koZ1vxDJuDQ0JdTM0CxVVDyCnO5oHdtUHy1gHs2cIOi0
OGTK/g0JNi8YDQI0B4A6pLzjg+4omPsx1f+uvuPAxJttAHSTFmtqwCq3oI0BVuWL
BZaLbzAUoFOEmLnWa50TKZ3PuqBlCIw40feI64FmvC7LFIBdpVgJu3Vcdbs88MdW
l6qfCf/s2ZhqlQIGkv+GpkOJ3Oaidrx/nVC+cyBzGdHEoXethnKL3w/11A3jj+qP
JmsRRFJFV6pcu8ecSBbELh2Pviahyby910sEjl/difvVVmrS3rc4pEwU67c4ohdw
/5bI+uznesKGdnzTEeIjazky8zBxhKw+Xz0ecqR61u9xxczKRZZaI5g4MwQsiGXu
xbRRliRGVNX+1QUwh2fWXDVYx9M30V48wG7hWOUvHINYuqMdo0vKjNFeITnIF/TI
VcR76zyaja6c/kO+fZM5kXBkTRVLNfhh8teMDPs8MJLdCHnxY1isDLLddsRdEasl
qyrtAJXXlDHfXj/jGDBBntJQydEuVTQCpiVm2j84tecI3mNn506qd+23O0jaVoGX
J+e81P2bgkaroJsJiuBhntPLKRz5qy4HXpO7YpNBgMafDVAVB1z0ayDwpJC6NA5W
nIHz+ZwVg5DKCr6eJaFs2tmWtVTsqwe+p6dJiGqZwmSPo4895xZ05GHBPo1NMaN3
pNRyI44uEpPgL+Z9iqdz5slCfl6oo+343VXOtFPhhfty53Fgor5ebKs/0M71ZgkC
5N+Pk5zFZI8+O9KN8BqmEji35yW3K4c9PNjcfqjLMIqgca+gHWM5bqxxkkjI4pPV
LQ9d77lVhy177m5IidduvHOHSw9xBpmy171VgrvnomTLeele3ROxPomvpchssX93
095r9oFMWmXGn8s3spTjzdbjR9Hx38IAqomD04Ee2MRF7qxVOBg6TjhGdDiON/YM
XrC72ayra/PYQw7yFuvSIHV1QUAwwZXcIMzHwRjAsHzPLeE4rcNY+j1Oidintb/4
zfp98T8zJGIj97VquHbR2OVF4hXtWYlH5VuQlf3POYTQicakOVmnvP8TP3QVdLyB
IR/DJpRZoAUipfVFYiuXsuWrUFGHjhY2HDY4n/XU9dkKEreAU3fUSRm+PXexkrRB
mYfizQud84grn5Sn7a/uXahcRufDQMZyOErnKFxcJ3vGUVJUOrlIl0yPMgV2mJPq
b+5nbbLBRHI+RmjA9Pf4VAI9MoP/z5+V1/WFPqZim3Uxq1sTJ6AtRu0/gLGY+kn2
lUSfuXNfTSS6nQfLU0G3NbkvDDoVALCcI+se15tUvLfTppumpmE+BiTkZTiVByCl
P4IGh1TbgFWAfJ3LdvemsfkEkh9wC1vosa7VTAuZ8rTW/WGx0G08DvVKQes4vGEv
yXsXTQCViWkgMXrek+O6SP0RKdh+SURquk4So7TtSnsJJw83Njs+T7HBe8draS6T
Kk0Jt2zKPMQKsK19Ew2xg4UEu+KL4S6wlSmtwMy61OfC0P8A8virs8WmVrUjECPF
L4toV3EaTV8iZAntUeY1rGWUHN1Jm8VEfDL0nx78u47e02DmkwNTyLpHYDex/FBQ
Nmh9iOsdJklp2sZTYZ56/7/1dT1QVQaasgbNzVHb74Gpm98/Bg+0mE3LZVoDMHOQ
EruIfAz362vSf9Fh1IGBrqvNB7S9F/W/+WN31GuY9u23B9j415aCNxCBf4yYkkTw
0xSMNlxgxKYg4p4ggJr7gjSRP0LI0AN2lxJSBSYcpy3BJfXWkzMMSpjJ/zddr57E
9wOnerstb9RpvBb0OoW2BLOF0Vq0/v30vR8GstDdIQdN8W9zJO+OHH0CnHT2/+qE
aXis8s48QYKqYuAYo26mjnjdgEM2UKxkolt/35afVQLE3tf8K+dIV0W7s8qCxtUR
8xgZk/sGBy7eAlU09UBbRKoqC8L6dAjjxkx1Xn7Ku+y5cJ/U5U3oVolfB5ED3W/q
4NAGlva4pXIYkY+qUpx52ntJ9zjKA0GS0xLpC6D8ep7ll2gVon5oRYmzGCVjln76
lre+r7qWaRbbb6lO5OWmOA4hHWrKLowsRHt+ZZBW383dzw0PEy2TNH/F00ZruWgv
5wSsJkQ99OxRCg+a3XfItra0HxcqAY9JgT9NAMZXaFFOH9a5PIn5Ozd51PPb5yj2
Q4tVKGrODIm21jZF9005pWGB6NE3dJD0AW1kZNhSPkXMzyUGr0nqg0LppKmGZdIx
QH94m53nvuwOmdXSC5mOqezCfUUs0G5GsJBJXd14sE1Q31sTC8uJQQGKMMXJDL2p
4daoHwuVVuDWJ9lsf5Rj1QWFdG363PftUe/TmfIbMk9Ck8m8b1KnDBS/qyNLLv9y
kAZDfhiaRBhVxZsc/SoNVw8K36cDy9DEJL3CvS8vzDavkeECMzSM7PzGi7TGMbRi
EHNF8KUAx7WUpYSq0jUMFxiEBcm8Gwcted6GpN+mOLdGfZu4mHNJtJUSF1oZ1m1m
o9nIoMdtiRyOf9i2Mrvr7s6KdULmgSoABpTpqDOY7VAq4IhZlWsHyCIXuWzLfxbw
N/jjUm10OjldAjpZlXKb2mskWfwDrrglqJEdmvSSbFPoy+JQgb1z6WbDeGXpa96h
UPZguxpLE+ga89TP+T68l+lTYmSDtP6dHH1qmuYVq4fNXyJ05rNC18LDEhQv6+y3
jpqHVDx/CaqNDM9e4u87h2cPGlTuCjbpHgVkx9EPj8vyoD4Le7JHDvtCq/mcB1Jw
QdTNWySRh7efD4uEOaek9ACWPBiZ1CGr7b3FljIrAMPqBfBbWGCwbUwyWCbXCGDJ
D0+NQYAd0v1ILT4tz2ZFCflbErUdu87licQCz49BEHyXHeSMhaFXHywbvwlPLNzh
so8bAS6LAHEEalOaRDLHX7Q+7+UCnOSvG5Ye+ObJfpR3BDJfRVSsxnsKchbj0H5B
o3xRtIezefznUFCQ1bzf6c8RnTNk7Nj8sDuVfA8/7kJbt6TdNqnI0xIWNFgoPokw
gswnIrLlXhL9S/QnJbWCTH3gFt+X1TcbvhxikQQOu+7aarOTCdeyWsY9e4oawiOz
HYI44ykBlGw/gkTF4HzwsMEZoUQMDkidwvO/RvA1jQyC/OA+p6SFli4DkB8TJ7iL
iBGkbXk6u+iwJ8g56pcZL9KqadRrdY98sU3vGNINKqq5KOwKu+2aXHsg0J7cov9p
KKf0DpjBPvrViKWjLhLGo8QArj5SDg1pkQ+x3wOcpCloLyWHtRgOlWAUEED6MfyU
Umz9/vzJDZnBlVc+7r+/9PZrmCUjncorz/86KhJQ19Pw8Z6jZm6Zh9KcXBzDFXdw
QurfNzHTOEJNVLoHYUNuI0elsZHGBW8xAaUpvV9VHUt5jKmhhb9yfecKx9pObpSF
T4JSLtd2LriOEy6tMoYXNsAt3YwFXytWnjzlTcjR+tY0t/foHysZZ9RgAl4zmS6b
031kFkp0vGWgG5o6NoG7L9eghm4J3gXHBi/TVVgBHeSM3fgyZZF/Ik8jODxoK4nc
sO5T+9e34nsMOokoCPLmcOhHJQUQT32N30k+PPa3oOqpWDTPXkizaIxmTymS9bU3
+Qw9yhKg6BWACMLYxh6zBwesN9+35R6YrFXzsbvmkWmqTZOz3iPbUNUt4ZBc8jbL
9tud6LSF8LpCfX/aD+O0uW9uA45782nrrniUsje9lVxQeoiHduQtPOcCMH8MJXhN
TonzOyMKAwpsFTKb5aSqrXYlyr4UerVe5cATb9Zo/Gd3i9hWdfK2PVIoS8CFHGt/
J6gh+gofabhH+NICWg6vjxFEVNSMbCRGA/dmE4iopSQdWz1U+WPECMkfrhp90c1U
L5jZzFZyqSriZJdSvTlB/SMXFYlMhmrruWVSQdzVaztcKA5mT6UHYOaYDnyW2CDL
pnYEcLr/FAz3yE0R1ei8qnnbsDovpertud0y1rGiLlOYZcak09bLNLJJVCxUJ2IG
rLfzkIzdkSpGchYqUeyqHAKKldULBfOD/ErB0Q1nh5sxw4IVRxumj2AWn2LxlXEj
4Zc+5vxQvR8Zg3+DfysJ1QxLjmm0j9wTsI5gsm6iAwV2owdysMnZBK5USWXgSRHt
5qkNE0dUEtY5sF4KzlzS5JbY5qHcQCU9jVLlggXzpwT//WbZEqJJpYDbtRb28rY8
M3SmXhyYKmSKvsiok/OvO6MmozbHODuZ2CKRhJLPxmvaWWnNg0u+oeeeNYAl64BY
ev1ZjPuHTUa0a+EI6IA1jUh173EP8b8RPzO/NQBxo4BAPhArxrjF2y/yKRgYULDp
jUYhbWqsOJEMU927KE2jzwOUreOZxw/ORfxhNP+3LkqTDBBTl6r6VAg2iqBkIAcN
W2eG7FBovcSRxYY3+COflwRL6pXm8o9MbcNMnyeQaXdFCIXZt1zJ8W0+DUxxyEKm
xvO+YhMZCs4wlPhhSHHJhci2QILUtdfU06OphDaiaP73BPFD01zwD+o3BreWSk0g
QdM9N2kN3f/b79Fg822uJxare17cOG1cazn/CygJ/nlLhM9/Zqf+ahScLYQWq8ad
0UvYj+FdQ646UBBhrAAWf653bQQ67ksw4HwHDxV4Ke+A7uS4CKyk6xz2U1JHaUn8
KPsbi5zZbmlwkgBT/QnR3V0qtMBXZsqvWC7qCIdkVtl7PMTSry+tNYyMehtgssQb
NZoBcqLU5C8AnCf3D3WX+fO8xEjcHSgdRHz1bMmuqSfK78HGl/gwonr+6PwGo/7t
CTSTCnfKyvIMU5zAiu16ZTWekh68o9le+fX5fnCC82lCcM49LAWo19E0KWLi0HTo
x0DWp3dcJvbUssjJiQA+PtYtiETCUQ7cQjcnKTkAjSbStAm75Z7yQwZwQ5HoDeY1
i9dl0PPsvzBAAJMWztkap+N6/vsrbeM2j8pUCVJkdsrA828cIbE28gNHCmp0kSgw
/x+g92SaMSKtwZ+B2+soSMEeTmvZxyalH6RiZRYQSQJJBswB7uhmz84zPZFmzNbi
3CP+Z3Ttan7icO2QIjOv9ZFAW59htMX1lbqYVxlUR70HUiLLBt4kmzhKFzFvbYDh
FAw9riK4g6by1Hf5cYSjM2o3/jRR1RyTTX4zl3RD5fwS5Uyo2yKmeZUjb2T+1SzF
LHUaLItnghtglDMtoHuMMRrPIRoCieQwkjLENCTOgiglJeld22vky71K0v4Pi97e
cZgp9z6vJzDFdMKSfboSbm/3L0pdRuVq4YuYJNjVb5bLFpRF44HtiS5qFINWjiTI
wnJtuN1V/OlMwhji6rHTHhrTBcQ4oJkUnMnBDaBN4uQ2cRtr4iGHUs23hvhRmLTy
uHvP26JgtAefGGdkovE53FAtSY3qcprEdOWkvLiJUNYXxeONti3ih8bZAJhvK3bA
74l604sRExQetRfCU8ohU6K/AlyO+VBNl5pM98PGapssTpmNWxcdc3GSNMAKVlgT
WGO9FqnCo7McXaxYl6cpbi8hyWRobQAqtKtpg3ktwHQofH5oUL35L8ViDpGeFxak
RKKN5ETkKuGT/uzy7CltWjJS0mUaGp19JOR/lbR4XbPcuJY6vaQi1SDOAoT52htl
0ikFX9oCacnyWS10MZZEVkev84TzVeVOYsHi/HhoA+NVrfEXPQqg1qa8UUEmPQpc
nZDQ7K/wecnTPTXiyTuG3VB72LFAXuFrt0uLR+4VDjNw3q53ByuLXf1cjZXZqxn3
yiijf/Fn/lQ+MLsQ1mzpE7PWcYMMaEZ5B2sAuzOzburN9ywH9rn7UpF6fd29dmIi
BcN4JntZvxt9IhE+dyUaqqSElC6krzvz90g9H8Bx7op5YhpHGmyjlgc+z1nwQiz0
P2WqeTLP44GcofbNzFTIhgG8SoEqWNYTNhf40+NjUi13wj8J1dRRB/wVLjokE3GN
/wVdA6E5Vc2cAb6OcCKBhX4lbSt33lLQyhPqfOnNJD8TtRUuHrJn5k+PLE8sxfs2
tSekOS0ldbQHs/k3/oxXD7rCxE+0wJjliBcJBeShq1LJS9CdLR4Xzo4B8uYzJZp2
gIAWpJbG7j2SmGuQ+NKVS5TPU+49AvviQVcR5MC0yIaxm07MFYtLy07pckl29jAd
sGVOB0tfxm+6UEDiL56qE1/2YDj2TXXa+irN26EO/Xl8iOMVLtlt41tiHe0eZP/x
olBGOI2PoK818WuMHquh7ucLaGQBCl57OQze8fnmqQotDWMSU+9CMCY48rovKgBH
It3IA7Tw7Frob5+XWbIVCxyNyueWAKY0FerIZtTMEPGNtJCd9EHeE3PlyshOmzIU
5k3HhB9W2/xYpk9obLkpkyWOuaQtH3flyXTTavvKrmkCr/DPGBvcPGlNekI1SUuK
l8Js2b32MxrYypi65nZQMsbFnmi2Y54SQ/Dy6mxG0htuI2vn5W2bLYPjFXhrPZvW
+EVj+DW53dV7CVwNug85+Y3KBl+lCc7oZUTdo7RfSRVTOd1li29FS8x77TLXYPhI
SRtKEktJCJQy6BZkizDRpld7IK7aWm8lRyGjs59XM+8ft7mjtfS4lppvRxH3lZA/
9XpqAOvNmbeijYuKFrtzsJ8Tb2eVyPFi+ukw2ffZ0uh9IVVLq/MnyN+bb14GclgH
UWWY5agXKaOg+k5zMQoCOfLx5cr++4Y9CwEiBOkeZ2oORwYAdiQ4Xrq/VUASJO6K
v8Wpci4YYNj+sA1uK92O3d2ifxqNaLztx1DlwacO9ujfIVFPxRAydemxEiqXJxyl
oUBZNdPu14CzVLVnUf9Njbh95fZUVPdCXJlzLYQyEB1/HSRL2r509kRY3yOqrllJ
q2aXnKZ37HwGBI4uLIH2a8lbeK5HV4YuLIZnjoX4Fd2QC/w2HaU8J83ESR+coLgK
dp+AeRFvgPAyQwB6+fZF4MQ3NNcpDW/FYoA8OM/npW8OFd3GKEY8e9h9+72G0uPf
12l0ksJ9wbu7ZAB7cUmI43rFJnOCKTow3Sux1ubpLseszQ5QvgAKchLEKhK7TOgf
RrAm1fDJ2ZBjw0O01hOEBxfqFJe03f+tdy/WoYgU6aq3ZSmWcxjyTpLfl19y9aeI
ukTvd+xNeS7CQZpH7FYYc2Y6PtFQXG8EELY6B6Mx86fQZZ5+WE74qqQejap0cJJ/
YbH28Zy2giaUzz1Vuhohh7SdWMtw1z7e3GEq4Au8HumXMi6+27mdOZGUQPVri8lH
IilQsz9927yUbWqNWc1oz5fAe7S3M/ucfCPdZnSuAHO4nMSEypwCv8MplfVPXt6/
vSdfOTnlRb2pdFp4w3m+nKSQdhpUf77MqKcYgZfIrxUh1yyYYNjeaDn845rFWRHi
SATWsuBkYqGVhS/UEGJmrmdERK8hQYrIWX6qEZLNTi47sEDaceSREJyBIHen0obO
OBFNtHKCgwS03y6dBGdhg0QvAhOG81YLg4FBNRrp9Y+ooaMz1eDtaknTfRoLJw7U
rA2cWqgZ6Mio0XZ9Jx4KsaHZ5ckgA6gH13xMtftBkrLqv1EPvBEQsz/A7KfCnPgD
kzBgWlCTg+G7EtrPHr8e9WD2s3R9e58V5FF9R7gAcf8Z7DlnwXrQNQkTGu4ems1i
ZROo5L+isOfsJ4Pt1+VR7k7+8DyIAljMNLixzIqoqOIQQcUKVYtakidyN4QM7fiR
dFy2Qsw4FSXgla2+kwxbA5h64K3hhcTVvi8CDP28hL1ciVzJJk8cePhycoW4QM/2
yoYE/+otcb4vTs4DvL/0MMWBuKIS062JAmpKucIDpq9flBA1W0S7WFsKmYCx/svN
G9b2z3prr2oit6f5rh+7vbSfbs+iTgH0LomTbPHT08tQ1XJuzu9oB/n1SySvQJu3
QN0o3FPoOrW5CZGOC8Q58V/3gkVai984V78O/CLd6C+3rjtFZJfoEyrcQhS+j0K5
7vyXS/3jL4HekJVfm+NFIzSoqTeVLs9Ch1wttcHn3krZLag8Eu/D1owFjMo7Zx9A
Ud3zAGFxilYK2Nf5gAxWEhKZFXFZMUqreFGLt/qwcA8RxnMYT3cWBlVmxCnakv7r
aVN9+B9BLh7KdnBfEvCv0UalBEpvNMYU+WIpSMMi5oyAgDcPcQL3TzNYToZviUWX
VlhAtd9P3c6fAi2mSQY8e1OJmBBRAG8sT8dVDymLLGjq1jhyFdMXb0pULf87uRLI
GxEugxkiZLRIn6QcuWVo0UyiUWZW2GBZ3MNdKThxP1qGMtPu3aWOc6AVzsECEODW
FmlaNL9/pBrYikxsaoOj6MMxL7XPjwA06Yfy/6IOgLDu9GmvL0k8rxpZrYUxj1x+
FsbLpWW2aNy/wmFMifQEAuCk6um0o3BAVQuH7WQpPOV9pq3uuxmrKXHe/XOZ+BQe
XiiBGawTdb3h+qeAnAz3nDxLnzb/wW4oURj98y7p6SzHh3xQwhogQf9r7XPougPw
FUzLP5M6k2/+qCqvanZNvRnsU0V6iqhC2m6J9q/cz/HkxtnW3cA7bXwfgPCJFyZ+
dzpciYCAjQXAIR1/lDSMkAyaRZHij1bdf1tG7VGgJwXyeXtK2nk8PE/JmpphkcAQ
MNcnRzThK+MhqlUYzgenGwPnHILhJx+pzFPE0VbzoF2U7jvwvOUy8E4WBX4M7KAI
9pmiOpcFtp3D3Ew4fzVyhnm3eitVm1Fhpm4h1ROne4NGzu7lcxIzcFrVof7XuUJo
SZD7rEG9uUXbl4HjrUz44GCDUZAXdJWHUbh4keOJA2HUHhf/O4c2UPZ0z2XdNVTq
jGknwOnVGs8ovTMj5waGjwGtCjpdRcYcZOtRPHKDLmrK5VebeaJflnZwG/Fs047r
inCyE0S5Te3uMzXGBx84JoxVctuH4CBRLd2sLFa1guOMQsgO6QRHi1eU64gpf9LR
pyuHNLDNk3EZhDeUJi6dvZrmDGxK8nJ7lo9BYRUvu8E9lQ6kFrpYvmPENdK3S5zu
RXNVxWL3iQ1TfRBrqOt+Eu73vpvnuCq/KImHj4EDL7idLu1H9emCiSY5GBAK0yq7
tf75433Oo5rMh6bwOHBb9SsABf/gKo4OAIz3Ov5beErmN3u1nshPQiWJpLJ7NJx6
Rrhs1Z+Gt1M43ZQ8/aTw/PgQ7CNytkCxtXljidfYaIUT/jwidzgchNZz2GP+jlUJ
4AT0FPs6KCA0c24b3j4ZXtnAUbngi9vPLkqZPjyQ/Er2TyVucDgUukhAWYSYEuSL
w2RK76sxSjWDL4987FRahym78J36jN7+DdkExyMXIVkns93cKxJKYfvLu8ZdfExn
rYNfX9MdxALR4jDbj2WcWk9N5K0xrDjeDFWB5/f5WhOXspQ9MhrF0gvhzbB5DcAl
LCgK2PGznjl22EwoHuQNIO3/obcDHa2Tokx5jvbz3mwF/+tB9nsepAushfyeiYTV
A/yfVZEJlP29jrP4hLdVa6cf364eassSkFh/L0wZxfdwisgssg8N9LvPk4EAms0y
WaFd72b9ZhI9vqiUOP63pwtEqGpxordVsCGAtlqNHKDiBrqEf6nCljqm2IlI6ngT
EUu9sldncJggyq6tIBM6RHi/7vmMtY1lGVk7rHEj7mUnI9ZWrH97g3ciR1XXQ4hk
AGi4lehfOscVwFctfYRopyorYiNwTsVMffqNj6/2oPsP8QAS8jkaV6K0HOysS01e
YlmRnCxT+JE6hxocctgpz8PNeD7CoEN0Tv1sf6G4t8JxSruEg1DZeWckxWZV2L/5
BWDh7nSpPt578/tdU4N9zCweQFwvXmmxud8pYckkx5KiCz0SkofFP/W2VfnpW9Sm
DGUrnBYq9cSecBTY+LsTW70zK1VJfLlhdJ+C7enQuWkEfsID3q1n2L+FHJrVltxS
ng5eI7D3tC0Zwio1gmfK4Gnqtu8voA/aw1Ea5qVEg4GlkZRF6JxSChp9NVtdUGud
5t09BeeXk2nMVhV9ucZuE9wUkSKCrcvY8z5ntKcylY4wDwMWqHt0kx7bLbZPoPQE
lNvt9P0kTtD/03nj7H6mt6PovvXrFvWs8A/S1/O3HKS/VKIFd/WkWA32+h5PSGtt
AOK6ljj6eNdXnaTxi4j2xsgEeTfposyLRWGEtbunLGcwNWNzfwjCm5/AsHyfKZzS
ss/ATdNvGhcJi6XHUt/vnjLscKJ6Cyal+nkBfoSiT6B2GzxnU6qRUnDD6pbBOqB5
8vKybEZDcRqhY7+OORE0bjx0WFMTEsLgADUWUxWD6ySzauQv2ZnfrU4jqFJHptWx
nsirznB9Hg+ifRD6FEDbnb1fb50sWDVidNMqVNOX4LyAUW1EqbUl+mmUtZ45491h
HpC9bvceTACLGmI3L/sWUhit84GBH+vOzJHD/1IZTuUXJgNjc9oW8j1shOCAl+hc
KgfsiW+/HnC+8DOgOH3rC6TzMLdB9P9Hdc9Dzblwr/39e1zArzXCwvi9gltdymAZ
kVHK+WwHouZlA5wAaMh1d7SHHMSd5pK1N2M/Q981hMR371fgJqg3GAFYSqKHxTDJ
Vl1j4d86e5OVQtpZ+l9rCEG55CBL2xXbLGCnLkqdPGcyhqWIbduUAEFD9q2qxyKi
Cu3LzlPlfSJlq4a/Kom+xl7zbjwXg+fUcA8VtOCFN03RclQpb29Rc9ccZ+v3J7cf
EfQLVyPdIBTVla2qfw4N6Op//fnZ/OXQVzr/G08mngPGanHfAMTkfNiwA0amsc/k
S48NjreOaso/u0mFJbPb/naOU8EE/vRK5Lt7aL2nUtWYZr+V1CCr8uaO96UyUR+J
I9Oc4lw9B8Ta6rlYQOzUxBZUHtW1pjoNKoKTot8lHOzLlNx3GVjOwdQTy1XfL77L
qUibDRHdtMfHgSdW9XjujCDuLechELemsu/HKb8gxERZl0cNio+NajgDeNPSPUBL
+LmbHa5nQbjvAN68o1hCLEW53us1WmZXxuV7iNwVbomu+pr3bn46l5IT5TT7+wVq
QrHAXHkNJhLFif0oqEZQH6+Pu6mJdjJl5UDBJ+VpIUMWNgVwKiycNXIqNvkyVO4c
IQEhHQZeh1xzOVOrx0NYaGyXeu8KsidF27pn0yCC2LKBUosc7SCJiFb1rfkz9hjt
YoeRflkEL8GFZ0/u4q28mDyO2RFevFGNuixjh64tAxymeBicUOtYitCw3hS5Qrvd
uPT0ISHcPS/+j76s6h7Xs634oFYXb1fVSdkx3R+HS4XJ8FGP82WCdoU+Pbvyn2Yl
RiVjCowq0dRO2uHOBmqWZ3sKZFpgMhoMV21QrWfxaFDTpzQckdOY5MumY8B/xLlE
ZWQ4UDkkH8ympnFUpybzUJtWl/+f39kYYKzuNU/5mL30VzgTXooze02rfbMgDLhu
qGXuUpKvkJw2IvtfNB+x40tRYp96TtQaHs9/4Iym52P9GgmREJHxlJauil7K8hn8
8dbAERF2A2rMXnxBzPApMxOhwaia9sQaF9bfmvUnhpR+yGDuxKcYRdF/a9xgfuBy
qh419Pqhtagm/T4zMPgPXL1JEQPZrm490IkXuCjpC6m0XM+uCgpfuriNynHPl130
TpitAQJCt8tKoiewB6163LQXY7wYs8N7Vudfe0ec94eDQ726k5FKpxHDslwPmKvZ
vLoxFp+7Gwfk6KoDZRN1IsnpnXoBmLJxVHmA/vMiYPARozg4idHk9aqAlROGLZep
0Eh3P4TqZZSnb1p2OBKiXksrZeVTQolx9FUzb+LrpxHFGgjfgk3Tm/MvR0zAt2jg
R4zo7lZgIgSjSJPeBNJbOPKq6EFr1mdx9AInyha9SO3kgTeaPmBottrwSaZd21A8
0dTG+GqQGwipmEfC6BB2YkM6vepPIGDldeirc77HK4FRDt7wLJ1ENhfN6OD7TheJ
k+cQEm1FcNAM745Ez5fH6kldcKh2/MMxII9cEbZ8F4URVR6imI6aYcbq/0RYI+2a
okcKF2qYSwKGOqfC08QcoA92Z+PetK1fNf3j7ZwmjKldeJzIBoJS+iEUHbA584h/
ikpoW23l+PoGANViidZs5oT6LfJTrHsdkr3eCSxHwls+Kldoogu2RTX+S2Zh7ZHh
o6hPVWr+CbW/Xn2duIEPajyq1scRGBLvp+6Z2XcT0Pw8CKsGHKf/Qw5VAw9kiiat
fBvIROXjaOiL3ttFbu5LRMdSkbxlr8JcJJmoIax4hhWzjRZP786DY33Y14JFZ+wK
pn+kF4i/eOaWMkaJ0f57BNmrZiNW+E38O2PVA36fPYhR+xBQ7WLEJ/j2DglULYZY
uHI4Hiu6rzdeCE1NFvOCxVqJ2n9UrO5wth0QD8ByrCvpCvdPr9LfBzH6jAOOXvNh
oR9hxGZXtQ4YYDxy8q9VAHgkgvF3D7yQPwS69HwQWOSFriZhm5ZnAgIu+n6P4ML6
1lQluHWue73wOBI1f+x9S0eZeLQLEDRuuJ3no96bNdK3wDF0HuSVPt8BMwmlpITB
fBiVRAiW/heteZk3ucNBDpWhFdU5RZVR2ilBJpvhdij3xZUQ+nrKUkOCJPOz0p+E
96RctLGF15+UEwd08m2tKpU0aDZ7k+9YDWvmODEHYKTUsXIrWDgnAq2O07yHczjx
sQaFWiFIRkP8ju1kv/39gTYFbdafXt0cFI9wndHycmM/izhaH53JNB64BQd8AQHe
t1BrR8yPiOdb/9VVec1tkEcAXrCzAQ7hFykipp/tU69xK0DztmRE/wiXjp403UWH
gPRecTvR23namiPK3NAu1Mpw57zyKmrEyHFhCKAkz5wJlvV4t7SFUazQcdtw3KG0
WBkeY095t04yTUqkuNIG8Jrf9PRToJLEI+qNKmDpdlDaOndoD0pWucsBGCVfL3+0
HGXkRclHrGwX5ekfL/FOzRnLn1dC9fz0Vyu5t+pyPVPkz+q/vtkVzxZq7MLFfwgh
Izw6qIpSy6DNpAiOlKEM8IVXwxYt/OdZ0UNwKFBZHik2x623t9QfkzTC5zezsp+n
mRpOCQlp6Ts20WQJnIkmf7DnC2FvrOZEb3BsQ0kgyH/jtFiSF6BrWpVQPmk/mgRz
ldY7HpnCJgX0OtDC5Iapj8yzdgiTGzxx8cyyYICXRL2br0Kp3Z9pUTM8WCLpqXak
s3edKJiD0gk7pDBF4gdEfZLNWzIG39p3beMhrRvtkPZmJuxSi/6nWxwC50dV5RaP
zSVux0lvNCasq1sWFSYT9UExwdLpQtfK1v+rwdaB7BCTYmEe4cz0M0Oz1yfq5DnX
AktRiknKrqZfLSlm0Y86hT8E5R+Wy3tTExGvl+dDvYGpccFa31rUDvuySMXmyEFx
NPj1N3x9mNLIZthUzhnGJ84xf9cPs+68imaBm14ZIuUjsUZla6DeyqYmbk9+1vkZ
OgKB26uAAPijK64BWaqadPm76MpZC/QYnFEQ0iDjTiXsE4CtlYYKRmwusrUEy5Qc
r6m97RCMllYY/WZdfBWWY0WWWRO4gGvcclv9IJ7SM8I5BDVoRotns8CJ94gVyvQO
h4vdxiaxnLHXD7+mS99D4LJgvy+Y/qZ2GWMfJa4zdYtgFW9fxNdMQjHtLQTrlryf
I0r6FVFTINbd26JoxVl/dZmSK3gVfJ3LcaP/m3lSbY4zaKWmK/tUr1lAMVDJAAsN
jdAfyhUTeUneGUrRddrUqEq1ouBjR1+yftKmhi0pLEQhdOuk1oW+2M24gr44aOxu
ADNjt0zBug4JpUKjFoyZQsxc4JVBZiWHAElyuNeIyHmg/NpBXXr0ZsKylXCtxCKB
lIC39QmEVLjGumIr9LdrO5wyxhaeZKLQP/8DZB8Kcwmhc06niodLfz7KKkcq+p0J
KYC40wKIqfAoYfZ6b2NttQig52XLOsxyHwWgKmQPgCzlvAzyjUqY8gH7dxaZ690l
yAcCP5da1ImxG6W13/aOsl2KaAMtnj3yL7FstcWhW2yORgJHxfYZJW43AaUid42s
SXbcYFFCr4RQfd04qnUGRQy5/h86t1Qxc4VXYQscjQ/DNEMSHUFEgV0B/lvBgWkF
HO19JxkFABeNS2PwfnLFGJSQ59G6ziRFq5dmDKQAfuDt+hWXRNZAHD3kZ+a3GwV0
zMm4Prsheqj6sMOW4j++YS+U7tP+I+jBP83ofKVFz+BUOquiStj+WNE+DdSTeKTL
MeqhpaBdWxP3NEYR0K1q8u6YluHI/oa4qGyCKBZnDtfmUOZPV2Tv7NRK/pk7BRLU
whZJjD4qGdUsxEYeIVbPMPa7o4GiAGzbI8xLm72A3gjY/wyaBailNzBXYrjOf6L2
gvOlRkw8Mz2Q/OOKKjKI9ovLGsvJ4mCPfBIIb7dI/mePT1YmRQ9lYfsrNctC8lmo
iBD6INqBPswH+bOR+2qjDgy2grk6CxnlXaEnUSq0gSHgJTKtDBdan+Azv7SBOJtX
juQIqRpNg6RgBBaHVw3wBBfh+kIX5jg3M5Sl23n13hfq+8dUVE4RI0hEM86Lo6p2
xb29cJ/Z6UPMfv1HR8RE5tJKYqQDXhL18CpfgoGE3SiVsGlkHscwRSPAvY0cFe9h
nPIwpNLw3Ovgtkz+EzQmNhewSHuVaZvEr4LXFFuiZGOaQpTF5CKTNxlCJ9GMQqDO
qifr3piUAssufri9nx+k4+xTXbFg8m87XLbcl2o+76EaLpUIZ+Ym2ROFznWkpNNc
Zj230gdTeITQK8V/RYrhphJXPX9kLkNpQXOoOhj9NAjJH/qM5R9wLPqZNUMg5JZw
6ECvTsi2bcJT81yqMmnUvfZG+MowTIj5d7xRj0cH8nFUvF/++ajII+NBCUTO1/3n
XArxV00uGDqmwIKDCNe9tAM0F5sknRkAa8DckDw0MXf9ASZZlw9CXTuBGoXiyxpd
7k55j79hc/vmJd2yGeIOnyokjRPXdY9SmqXfLfOwWdTXx1tUipxXD77nZkiKWPkI
umfYqM3uVa0TsN3O9MZM86YEdxxouwCGtOqH/Xo6D0/UPcDVGlYS8u5GLYpxM7pH
0HGnTNX1o40zJ9hGhcJGndiXXypi4x8D5WUANAFiXiwJU8opUQNRpdHMBMsLQ2vr
nkF8f3bdQZ/UJWieaDuAQM+lzzePeZ9Onr5/FDbQurAfwrBFPj0MRyPMp6Sndmby
oRFG/uLcU38GsEQ4P0ImxEpBOPxLQ+HPhSFKY330IhcmPP0fEErHuN6BDmrcDSEc
exIf02xv5vV501VLNWWrluGHzswfv5krhmZLYvj43Fswf94z6N35TRrdy3ja7WTO
mWoYsNwWeHXz/3pvTvJ4724SRE95e+T29KteQpFtVu0RF3JAzTTAjSAHzaF6czW0
NWoMcp8/qtMIsuW3IYAcgqCpQTl/U6vmKLvQgzIgH6tNQgv8UaCCfVdHU0O1Zjfd
Hj5ez4WPMBydwgwgycBxr18u3SuwygsYxPAWprjY0vWAgR/hz6gLiM9+Mic6qnLA
lVyalKyCuDwKjCw9cG/dOjN6y5/asWfIspBilFgXaWJqNtMuzaejoBJb4Qx19kYj
3XEqrukIN9aKC6RFbU9OuBG7Om+WhPO7CGqvFmQy72WSir6T+XIagAOhOHpowuAF
WxdhzHTsqwcFYEjot5QzuPpku7YIgdJR2wwWRSDU0mRtQROPMD+QJOUY8+XY2N7V
CQm32AXcw85D8dIxU7w9EX/5abhx3fDHVkW4VilVv+gqlGJKpXvbGVFfJvisD8xn
3UX7A9+M6ggLiCdIipqBfJaA7T81JBkKi8/PRD9ofpjPqS7DiPF13gfItYRdWdte
YV7C5qQZaFEmKLE5qnb4pjIyb/oL56BQhtnJsPHGQr98XENGFD3ylb6kuX2qkrRJ
HE5OqohcVXUq/FDKy5SNhVw9zZtKXn9qDaVjwcrod6vzGVxHyWTskvPtIvYO3zFx
a03v1blUYGb7IOv/Dya9GxW1om2TgbEtgeeclx8xCE4mY/bitSfaV9m+7syLBmLF
T1M3h9y3za6jjU018yw0uMq9bA29scf5v11BugfLhFWgDsshScwochgAHf5j2KXn
WWyDmBrv4IwMVsk0UPnvYzNsFBz40CfsD2k3302WWT/IWd37DLMhfvpJ3cAsG8J9
6TH+lOmj4g5Q+IhOmy50A/4J/jN7q33rz8Nda6XC2V/3JNx0lWDEKubWm79K0F0C
0bDtmZ7QARccLXcZdmeEnPX8iMYFHYDZ7qyT1sqTk2Pg7/uoBk0VV0nWYeG+YXhg
fqeNamt2mtjlWgiY3iY+RMxOOeVCnuTAm6FqChtDlLvjc9kdWh2fmJFNGORq5gPw
Q8WU83k2a9m20udb/+jLAGgLWh3P2BBEeb7kawxAY+lfUZ3rF2p67FjQlt0OwCmj
s4VEG/9OTNnRc0UOazy4O5diOh0FehuPOfvrZzk96ZR2h/A2ROGtOGMdckr7Ua+h
Har43WTXdqr7fMIkKs45z+1+OcoMEgZqnTWSow9CZjvzdZuEFhdYwE4yM03Msx4T
aSBDKieCf8adBRPHN8r+pIPvy6MrHlvmEnmGsGqFNNrZVDTsFKxSAry+cnnVAAX0
YNofkCZZEH4tfgiuX5f+hpvJ4OVEGk5VEWHewdq49lFbuVfTo7baOBGALjyk6l1P
lJKTxi9wwtjONqFOgJ2VDGWq/nmuq+ZsTZ+1vngHv6wbZ28TkdsKGcSKKGhpxpB1
o5oxFOAR2oz+xjnoKudoc8xDPfHudAclxutWuMFpdNuU/s0+mURRX8yDQJZbKT7T
MglWhFIBdtJ+F8CdA+SWg3RrmDHelHPp55u87KSLeQvhgNShHOzQPBQjU8Pen7Ut
MgFM1JgTgjo0Ct9KRgzkxYI74F0KpL2eVQ+c7DGaMXNH/utWo+DXBlEf/Vzuv8Gw
D/bEbJbO9k8kfyyPMIhD84cc3930GEC123+PJ+AfFshkI8oBXBimMs3gqgUEgnQx
esYQuDu6A7M9VTDUS7dGYiQYCHTb77bwIq8u97PuygXD3kFWU+EBEHD4OSj5D5XN
nqjLR+HjvWXIKJnFOM4MvEAEdkfMzFZJ9AQaKPnOgDghlHe9qMeCQqyGwCS5CRHa
sDLoc/0EaQ853Dr4oARCIYWBrCQ2eG7zT1rS04JbAbLujGiAsVUxSuvJMbF5zwbU
vAxwW5IV6pEbX0mO8gPwiEHpaQV1RQxzGHIDjFZW+W7oMEMtYtzb2p10iZFOe9WE
NhFEIHbYAS4WQxZpCUmPx/qXy/Fns2d20w61ZqB2cCeR9vUT6RDUToDGDLkfnXxM
Cdu6aWoUVOfKAay4RY8GQ1OVbGc5TxYNStATeF9dF/ejc8DCRN5o8dPSij3RvXmi
/bUprvio3l7FksJtbZ7/uY6yoOv3tH/N1mIomryVyQ2Mfv33KN1AOyXwWVJOUpZb
WGlC7UBpml7DAS94mp1J144GOgnVXL15i3PhQ4BmrfwjCb2PqPNJVenUnqQvDuI9
I0+RL3soo56kTtprEaz1zzRYn4OMtCiZTHacygFjTn/7LGCQidB4yGvQTDJM+c5m
NlZtWRkiNPupWigS/3ErnRpBUv2JkUFCPpGmGuSf/YN6JrUcTqECds4Get4EjGlf
SCY1xTit9iMcu6ihhgsEBgJl+HtoW7pI8yyLyfDaZ6ylk81Vxw2DuJHr16M4u/x4
hhf081hdc7qQCRmuaLkbG0Er2tywnG0dMjhJjAW9TMM+JIpwlNNCivW8PNqSMrXt
4VLtU2QgFhC5d66mT75s/2gptHjC/kTFWZ8nMoHGf+JbczeB6ZE6VipO8OXahzDH
E8ik1oxl8CjF1YW9tCaKY9F5AfSSuY2iEbDc5N+b3Tg+f6xQQB0m3gBh41CqJ9ge
6IYHSjQN8U/5thZc2A5HYuFbKUXA1eRe06UjVaALyEDKG1glr8/7voKMimVzYjLx
QSyyGnZuTZ4xk73q82PIvEN8kZ5xxP+viK+9dWnDanwyOxHAvx5C99jUtCOW5UEn
8L0eMMFwFxb2soU9wregGWD45ro2C0eqPRKUVgh00tcdGPp76wwaFeTbJZcnALaC
sauVFj5aoXd2WxiMwb3wxPOgGspN4R7nRBdzmv/iHW0dC3ucwp7W1J2A1LtoDFFF
FF/rKR5uBPENAbCCLpcflunu1+Rg882KGiOhATRDADpFap2MiOcsVy7h4pVi6h5B
tLukpkpArZkzfGebVtXtGskDfePm2F5Q9e2rYUo5/oQCtj28llo5hjYri1TCVNH9
GPm9EPCAgcZXsNwMws6AKdEeuav5uDdfns89AG+BvlQAoZkeS8qLOdoWrjDAtYO7
+frbpoaIF7Zj4uMT0PanfLuP3z4JbFv5SC7slmw72YQsKyAuV0PWJi1QWjDNuNxz
w+zL/3mk1iHz2NgLpCaORe8aOjws0yWht9YBJG+rwkTYpl04m2WzAWCpMlEVhYHH
6j+xADjdZwoyMCiyc8h8ufyA4jKi82kvBQeuMBGmZTEicCuFz7mW+XUJCoF0iotm
Wl8KA0CdEI4J83KicV9kFrjJEQpq6Fa4vFbGjd9aSopFgpvXbG8lRntnZHFnbaIB
E4iY3ruyrDIECexaTXmLXl60hK/rxHY0Hyd4t1h2+9L1380rz4Gy2V7AaXEhtNpN
/8Yza16rCZgLLHrM3A6fcB/4CzYt7M/ThfWrTtYXUQ3021QV+KJ5rISN16OPfmvu
gtyZAbepgLaYesSIV1vj8ee4DNlodCiWsA7jdfYVEdDOVujIThjDLcu65HioVFTG
nXSyoX8ojmyDd6wj1TLJjeUIOsG7zxVaKprDI+7FEatA8lVbNFNvIIY5CivhN6Rz
krKXXtDH1Cr1KFPR6q/6o5i8sbiHm5IR0Lg3ibmevU88VL6i17nimBMGXayqkoRJ
+wcBTUN9+ewvfdtfvsLIJjt9u6db4Ld4ZHCDb27itu1cyrlR3aR77as5vBuVAKO3
t6tE2HIlFNtlPTt7fMeM8+FPeoWnLcme03FRP276mi3w9BmVMbEA3eCL/hjemtae
gwEi76n6JnDLN33ICme4qJ5EsCluPktliIRlrPy26W108DYcruBaQjdfdWVTwXHD
+DCNrwPTb4uqp6xgP0J7g38Wz34QoFVVj35WyShbJfdUTX+I3rpIDZ3ZguJ6ZVLp
RYc/RMmfVIJ3n3hKN1mDd4nbh4F1AkxaLJZmDAfLOU/qf1TU7v6LHdTMMQzavar2
2Ltq0fU46t4P4WAs7wPztqQkDwGyxgMjBCz826HvwFGuz4eJ5Sst+8qUTKaRAzra
Q7dnZ8VVcTvUJO8f8if4uQGeoVgtsORYP1osZ/05vdwq+/Ax5H3LfHIOjxZ0sY9i
1bIiaGROhkSBDZAIpBI0Cjv+PlLhvHQlf5lWiY7U7txqIPoinarXaAFTVyo/NX+Q
Tyb0WpQEDtNX/wzyevIxYNUhO2x6SFxxC/b/cuahBOJ4qtu9HIqwTmVdsdpS8ATS
aPtNvJ7jdjFTt+bz08KFM+v2E1sryJAqtoCYZhU7E9bOJhC5IxsXk5MIFCd2EbeI
LV94f5IzBB/g/chjBfv6d0mHwiI2BjuWd2S/QdjvCvjoAsmaf50bcU6ACnsoSeSg
tCclNQVA0REoeO0l9h9w6vojleVAaW3m9avax6fQNaWL9vHhggbXsMwfb5C0nHgK
Xpo1pi4cUr/rwFkb20rWRoQDciPQFyEY96x4TxJXJ0xZQBFQK2fV73RX439d7/eh
xspLMBNea1jQUQlNTgcXdi2pVbvPutc3pfhl6H8c8ulmAU7De8qMLDwrIR52OPOw
Wv6SeHNGbkSmeC1m+LdqtkfZaNUbR40bLO3g3sDDSJVV97AdJBaA+iK0oKaM8tWg
BeUfGyvD7pZvZn17Tt8zDuEyhvPb+hQs8uKh9VLh1hL+7+S977kbz1z+KCjJAaUa
lTVVFP+vuQhjGvrPycdQHoRbVfvn83INOJXwhhxn1sVgfzgX4ZRTerqwr3aeSsTk
9z9pb1HF7/CPIzvwh26IRb2nl7Lg6KmVHJKnlfUEAeIoUXqPyyKNlZYue6hskgr2
7hTcqMSf0H45ukUVM+jgwyc/yoTquj4ntPmhgWVrBjtGXFCzLJ9Hm2a8SsLJvyc/
jwA2YY9++V3Gi1AJi8EYUY5lZLV1pIbAvhnorSG02FtSFjX1GVpmNZEQfkcNKXj2
zEpRacVZ9Tvi3rBtmlj6g2yl2ZfxC0Bxz9YTN8rXX5Q9cwUYgXoxXklj+Z8Kwq3w
OuTG+EqdPtL3QIurJcL9NcvqtY25duPb9fCJ5n7w+TKQxoWQ4l0vZ3Xftf9Rchd8
YMCyBY/tOlIrVUIsWWJlbdBmgObAmp6WiP03FUAtci9+lBe9KAjOCj4sDOaAYICD
qTIooWrDSRt0plRT8n02VrxHePQBpzIJntIaAfd572dAmy39tLQFkGUf129WHojO
5Wt0FYh1EhqTpGM0GdAPipxD/ntyWA/1SSEY5GP/GQdTxJMfh7pFP2LIllXBtZVj
LNeWTSP6Dy7as5cBxu5O4oE/Qr8OOc0L0FC7gix1xKqJ8r7SDuprAaozns7Z+DK2
LfY+pbCXotLTdcYOKhUxV7sjCw13/DEOX+uf0DoTi56rta7npDpxkUf4BDJfJ5MM
d9VaqCAexC2erXdfbq+XM6AmbHZdHTx1oZsPKOWJKuea07WMjQRkZAg+pVdYyveK
j0JTyTNzn/8zQc2ho8BdBt7XmBdEUVfhwKhYvWB8T8Fx04cQIEBmk+ImqKqXz8l4
IxPaMk96NKyw9XIs6yEwtg8VPBIp7c8wUYszExN+5j4Esbv8izVlsC060xjDWG6W
YvPx6evXRGgCaKKRjLf7lSsoGhZ/VlIMwjVFEtVpPW1oVJnl1x2OI8d/gP9SEsjn
kBdgb0lhvPwS/0f2oGCWzGPWqqhq4Stod9+ZSlNb5QtdG3fUtfHjs8bYAXaUCpig
T5V9Jp57dcVKLo2bykZ7wyynBEueN6gUuLf/dhVFJGEH+Csa0/+35bIg9OXr4Fg2
uqA7tT1pTIc8TNIusrSdekLECJGmzA3XtvX1VA3SX3MKTs799Xa3XldDDb5ZvY3M
v5W7cBva0b+ax+NBk7LfjoCkjiGIqi+9FxyagIFbeL9eROFZ2bOb2lafsnIWZBw5
KXmy2k48Aw4Z6LyGmY4jknBlN0O6KdIbMXlL7A9aj5eKHSUVebWQRmis7GW6MC1Q
RBsMUmIM5/QIEmYWa6H9OVYmYWAZCND1K/MCNCwTcGVNICkkQGebfc+hlTTlcV32
QgEqKdCxGGDYtiD22mavRfQXp7iQ+oBVO+m+kYv9h2No82QrfzBJz/A6mUUotQau
pKGsU8WAM6+e4RisrK3CPbJDoygN9qVrPkjNC5N3uN2IrcT2p/RrPYOqigcPbJY2
5r0tJgYivamaoMrM8Gj3/nzuT1mfyP9pkA1FeSaGyLpFUXxfUVj3s31knrdBa+Fa
gHIPn6XtzawgK2SWMKNK0SD+iYkambIZEmPT9N9i0k/2qMtQC1M7lzwIeC8XYgB/
klm4vTGG4uLvxJH326yEoaiwBv/FuR1bUM2OW69YamtNIh0xdUqWDweHsMYFmH87
Y5g8AFjaSU6TyMtfmGh/dpFvm1+Fpq69X73xXkvE/ZZIk2yGJqg5/axZg6d5/K7+
qJ8vqUwruibX+8N231FwlIMtQZcM36JRg2/HI0pce2JXGQKZm1QvZeYIqavDRHnq
1AEHUtIbORAcSVlwOwm0fip+VmBuCeTygji6ORSFpUGVUW3nuwedkIOpwJ50wDlW
OBBVQuKqteeu9tiqJYRqBq/T+WNKu+TUYfWApTOSCXyBj48WQUMvS40zRnWKrl4j
vVi2g6pYqDpitp5dl1NDOkTAWYIaXShcGQyJBixUuIkVMMTa7+q2a5Z946YREx1x
QzPl7DbP/HTJFFshKXZV5eZBYL7j0SeBCf5JaAKk+6a9UQfSBru5/pdboPfF/DpF
nffWHybt1yVxOTGvj2CqQ79h4JfOpvqaRmUJdXvBEyJ5Kcv2WoznNARRwjIU73jv
f5ObCnAfN7NzTvRJCGITsq0G6riv13GlWyKkTbWQVIn1M5MwWCEs9MU/SyKc7GDQ
iKf/5QbZ0ZrSdoPDUNP5y/fk6tyugkZISMYUln2IDhPzZrfs4rfWRKzMgZ2Ljaqc
DgnoPvl0HuLSwQVGiwRw8Vxgtt5Ik6RjXUx1rqBdROhW03kgN35HqUj+rJP1PACc
0EsOKZmdhqxrCcdpitwE08XUR3uFrf3CLChwdjAUH8bOULAW8V2pWv3ByKZ2JwRv
r0AbFkMBn7JPsoy6tNzi23rh+xEGvnsY+S5keHwYh9ZLAb+Q7f1EmW0SGcleVgbl
AxIWJ7otse3jY3WLcHRfFLS5p73+nrMyxLeY18vvAL8+wclrNbGctAF/foG2i4B7
NmXAQ0tdl4LNzEQydizGfHFAdmIG05Xyn0b/wVTPsog6NrSJfDteCTqVKJQhvoTV
wpYn83cptphPfscoM8kRSinwA7ridgWwJujNEQMxUQQOfPst+5U/FfcLA/uKZUYt
JJjy+g6JPhJi9bvNMkBBHjfeqzXjJYse9Ty9EvJV15jTFg5tQWcVvufvfgN4jIoS
uzxK3xNIx5Rub+u1n4xwMyImtYMHgboBB+Kch4dgD6JJY09OUOR5WK5A8mi0WlyY
Rb0oyEo/PiwZXga9ole67JORLdFBRSms5lOMYLIRKbL23uvSEVATpExXt9oL1t1q
jLc7JsXuAw2lS9x+7Trq6VsAaM2+zuwb6LTK5Agf9wahpKK4t9vOkkVgI9WP2hif
fW/8HSL9AZzgZ6qFi1wfMuSc7G3/N+sboUpL6dQdPf6e3nSbtgEujPzwVpMdaypO
RAEiDknxE5O/MSkcovNvxptOGnTqsPjOP+ZgmyxLg/KSSIuREHl6rADcF6fZU266
FQDHOfIjAjC+jlJ6dwXBa7q6Am4GTLTWfecFcRwNRHtq80STNE4frag7hUoIwDXw
ZBEd795N7nWj96OsujfVyIaJcxc6RttdCscvOacAXlLtX8/VMWS9thk8JW9bAPDH
Z2yEiUATvyOIEbFbq/wAhhZYEEoiNx3hWz/HLlXpErPByKn3wtr9pdFyrF9G6Rle
7YHpc8ymWkrz63YRuUyQJjdRWFYmQp01Tg+vbxT1J3D4aNxhE6QuISjGf7xMbGFD
AC+jj+i6/od7nsyz9MDpO6LLsHTfz6/wAbOrXx3+Mhba84Zqc7N5bdpctuLPjF6t
1GR6SJ+kv082pvRfVxQsn7QkU5K3PfATeDN6iVTpak7cnJzuIfVLVgRSZGYbPjRY
vIn6yk0q6RQuh20E1CL7ePH04qwBmo/470PceOx+XecKNjz1sTIhupVyXTEcIpS7
prGFb/WNCGoNdgBRKst2QJszFxnKoTnbxOVG2WNU27zo8XPV31DoP5gdfpclam/q
2aMrngiNTjP4wV8AqzZ+RDTmRDj/HUwqAyB1fZH9TTqgYb8WOeuB4JoZbEBPO+ni
HaKe6N/sIhNrxUh9n6/TXu/CH4RGMLEC55XQ7wv/3/+Uqrd+1GnNFdV5kxkVQdu/
CIOZfpn1q3Crw4swUD4aQ1DYPOKm7EI8DJobETYb9A0q6ClnlXF9WFEB7g117y5y
2dbcUGTYiwoVtv/HQLH+9tN01eqQfDkgCc0DU9cBNc6xA+Af2CGA4Yqd3euFGXoi
5K4m3RW+pLmet/fcHAAgQjI434FFnfns/mKaKwspmO7MO/6IjbyPT6aZmbCrsRfy
BIm6PYYbsa9xtaLwsExvgoLu8U/0MOjqkh6LBTlKhTrySYIxYuYqeT2psdbxaEFs
FqfCStDDv+nWJB8BjOjZPMhuxw8EofmOBoZPZp8+uuZfC7/VSMIIdckYF8OP1DYR
NZ5hng9f6eYdGvIQMr+wtrTsSTJr+djG2VMKiOZd1EqXIK4DXRBiJsRFRzHRw5Cb
bnvlAfrHTOviZdjIJWaSPkXLBGHrhm+Lcn7xnSnUAux2WPMK3c88Lf7pU5lyIsUF
R+6J2Tp4wi4yqtfRDcH84oreG1DjmUVMQGQ/9KjhEjPoeYxK+0KPm24N3Qx+/rj/
Bzdl81VIIKTnewhubk5ECLS7IvMrDFCfej758g4yR6RfwuT3ckmHeIiQChcjNqdt
lAAo5XK7Wrfouv6uIur+DRZkefNBUZMkKU9LmRPqm44QkHWHPQMTm/c+Gm5/L63w
FuRrl1GefOrHUaIPgJp9jMhdiSRqt0mP9s2fy8t8e8mXJ8DS8mCkxbG0/aLyPgif
ozN2HE/kfrfvgoSc6vMTHwdlq9dK7pPdz/0XaFiENx/9Mq+3wKEEuzbBzqY9Dhp4
zEBVbe2xOk7oxJlebC6hvTWTK/MMiXq1KvyNow6GWQWrMK6FpK4mT7YZ8Z8ihE/9
YJ6SQw5PmzO8h+vBsC/VDSlF7puOlGqjfH5NPQTa8OyWur5Fk5k4qI0cBqkjJPN2
12w5i3cAoYWBQQQ+SWowFPTnSx5iodN7h9ZOK05I69v/4h8/FGU9ErTFCkI5VivD
FTggLcb+u/sl76kraKLrvDmZbeCme5Yq+xB0QI0MXT2CT8MO7MKcSezEqNWGeCap
29UwnvVqLh1JTPVKih9w/GwOXLUKF533+Cihm6xXZpTNNhG3x1sKlO91J1t6AWGN
MnJRT/6rH7XokM401B8teIoZ2E2zGCh2sZpEOoohXOe7zR4ugs9DTTanH695Hhv5
lrxkVpANVqw4jJM79Q8j906WI+cd/HNm3mXs9A4/LQasG1AAcOxZNEGlCo8qpnOM
1gDpRJwSZMrH6MaJC387KAKjVS2bXmQCeflG/tBsLqIFHQZgwjuNfqWk4MW20jBf
oxiSbkZqDyI7npmjPdlxy4k7PcQdc9nt2puReHFgCf7CmLS31VLUZgSNj+n/SakP
z/9FV3uOm+fwfNzhu1Wc64jbGLWVJTi7CYNV0NA/EsG3gRxwd3TWryiouVXTIHTa
/T8G8l+mjq0Nvz07lMs/1FGKQMTl+AxT3qoG9JOM++3p8nClBDqitgWyEcRC+RRN
lnJabCyFmxDCFMtDXgQP/XSShZcSlspXhS5C8Z+mfO7BxSmoLI25cB/+FvJNTE9v
JdfT21VplM6s5gKudOfqmSPDyvtyBiN8zUNgsQ1Eay2bk9s94pn9+MkzjLCWMKyn
7eFTJn9kGqQ3jLxwolVz9Y/o9AqZVJFJ27fCQdAHhrSafjkL+f0v6GQUD9Vtg17N
O9lrKw17BrxvNLrAdjHZQMD6RVjRZPQdyoxHDoSVqU9nM7d8e1s4IUQx7ZaSgFHm
S2Yb1OKesXSdBVbmDPZtIoUj2A7lCEXCnwn85Pt0aK7JGi7GaJa+bYN6CdoizGUc
V4eL8smU96vPerVjQgrSAs+1RUOtSdAfTS7+VuKq8JRiCvuT61E2Nq+bwC0/7dfS
H60WfPnDDGtIK4oEtU7dOI88qIDX4UurNYb7fxKEPKnEkOTE5vJjklDW9/hWX5D7
9QyC19dktesYGjL6vgaA8pMESk0iYBCtwaTjibyuK/BO87Gb7mpfk4ncny81HeRK
ZMKCX4LICLH9ijg4Y6DAh6aGIeli8DNCiVXSoBTRdRJWwML4RGUD0aqdQzaF04ic
ksp2UqfAAw3ak7ufd2wd/idkHymuTb100QE+FOORDY0hLzNASwBp2ni/v0SN0Tx8
ZpbLfhaF0BvlO5mSoK4+amfP9B//ta/MG2E6m8p4H9ZP8TH0HLW7ys+kDpGQbuMd
/14HHszeta88xKQcG2x7c4mpnu9MPYXHDPkWCwgsDdsfyBVh41XrUhGf15XwP/xh
sSTZgG6zP/QaHlg9LLkCiF1PXgRskpbjCxd2nCmle0Irsw/rZ1ksdJNHCyAaoaEF
uTRxA2oFM7AKKn+PGbuijcQ7hjXsmJaSa9QczV3pdN/gcaneTdn7dh5TszQNuGbe
nPgLBWHYMSTFoGnpsW7dX5NigT5o1tH5foSACr4XD8BVBs1JohZtM43P9NZHPZtR
3W1YtRGmP1OWAgkufj3QBouRczl8MpmWeuE9vV7JC4ziuBDqyRBBLxPqC4/9o8in
gJOTmEtORnV0tN7jIZDuwyZ3XjQfK12hmYnfadKy9pl5tGGVL06jn7ZbLA6RJKfa
gvzovuT2fjlMfLZl/uL50oFVNasaCMX/l4ewdBH5PArcUpJRsZrnpe4VfU9Zn2iZ
LRH5MR+dUT+tIKtlbVcwhCQRxbRuMARk6iBC/0MpTNiE5wYj8n9vieO3Y793Ap46
1RJ5kS8JVM3FmSNHubMj3Cu/vBEn8rUs6tBUGY96LMSW7gitXNFfa6ZZR7NaZb9S
uILeZzt+U4xvnwLfxg72eyWaQVPYiyV+5nHxYI0sJGTtaU57x+Gz6XOKwzJepKJO
eh3HPDwRj/uHImTvOiZ//7XB5TE//cwE1i0dQmHdFE0spI7nReAKXZqIjm4cFBzp
x1XLn4P6tT/boDb21Hizc2UuRGuoPaeinuOJ1CAEQ+e43AsPZJtdCaAn9Y58o09i
XX13frRfnnnz4MkQmYBig1X3sfdLtEao/kuueHk654/f3bLGCgswBV66khq6om8E
FU7EHrEUxySh2NYm019nJpp0xpMJFbh7gMSLhdoNCcJdDqEK9qGU+bdMjih1/48r
/csfVL/jpPxxEIIA9DMth88Yj9WgtSv1DlJ5DrBi0jzsiAKvnb9bmgP5bSRwXITo
um66n73TcKreqZv6j8Q0MDXIcxdLJI5zEBRFPqFEh5I59Ka4Dxizmo5MG8mFvbJM
eT3hsl5llGRo7OdfBqgZPiJ/2p9WA9tLP8ulIjL7hhiNfVY9oyp38ki3wYd7TkCD
sqq8f3JmwoFspcXkVQL/Vv1RtgQA/BV7fUzGaCMiFRFLv99mvc7351YP4pXCACqf
ZoymLAyeErbBbVKGJdzQeebJ9QWes5JKMCN4hbpoFxsO7oK7BQhbdJZAEk8JJ7ZX
W0GI5OBii1xl/i9FXxL0e0AKptoUNs2M4QEY+gJZ+1jHi9NgkNuinwbsx5xcmTLF
NmpIEKO2SSRPUHk1ABVh2oONUp9RDqsdHda8+h/nDZeyWx7mwUOuEUTdLt0/PrBG
0UYIKOAbIvidKuBQrkHWMLy2UFzQXzjtjUv9smfFBvKA49zqNnNjzkG0++AP61M0
h+VxvKMrH644L9vHPoAM3mIZMqEP+fgbgxuzF55+421l2gFYZLnz7KyfpA5FsEhu
U2/WLsFaCpMqJJ81zU68xKAyGgB1GSWExkhRa4QTqQjZt3xigDTVrmA13Js2K9hJ
vMjxzVW9XqMrtdh1AFBzlmhisJxt9oEruLq5Ux15ImVqqXqXYShWaqBWSwTdRj2w
Qv0YL3UNfhLd6LuHaJkYKR6RPdraw5r2mkaCfkNKO7bMwRi/uVtX+7TmckenOHpm
tpnIwuxRORAwkO/ARvfDWaScFFhw6Dc9EJPyYjvZdaCqI8w/5x7vj++oLLnBqrRn
D+yGTmHrkHKMfaWpRhImyEuSPId4ug49URjgKC/FAafmPJTEYYsZC42Oej4KR2sI
EyNtHcUgR4I6fNoMUhgkawWWz1C9P4xWrN1mOIo5s2U1V6FaUUyXiCrSELzN00p8
P10moAqDdQCOa2BnqJa0s6JUpmUXQ4bljOl+vxIvTre5BE7ulE76UvDAF0qtDiU7
7yZXHTYEvbBro1ZX60tsm69KKzOpurL4/qIdgJ3W+W4cVPPE2A8UJ1+94f4D+1Gz
Nhjv+RhHbdkfugRNAw6jsKGhzoghUfCwMho+PR5Kfx8PhluAdr+eXPoCM7MnZOUf
eGsLLbuXYNh3V7WNrz2ycAJC62RYZ0H1AJSOfovPQzCqbS13dDRn/QvNk3pubt99
+eEBv8hHyBYSHj24tLc3K9D8t/tU1OGIzlvPYetFZnEUodGDcnfYdbU31W+glP9+
kJ8XeG+GydYfDTUP4srd8+bgSMtFHuRaqYNPv8h0L+7aotzhjgAMDZbQA/Fdp5EL
EDEeyqYd/wN/o+FkpwoY2Nz8yvc6/AqvIpsuynMFNh0d+BqxH7zaB45orwInpnkD
e/4ad9+5m/+/1TV41nfK/mj1/dIb3QiHQdfMebCHQnrJNSYFQfv9fzdxBUOyl36u
OMLiC6dQmpBeHze9h7iJKPTYze9sCv24eSkZu0BEr13SAvBwl1CSRpsfiex5FhJe
FaUGrq55CsVNDtzP1laFkfUmtmdcUX/1mVD0FKfXUASEpFC7c98oCKlC/wB5DnWb
RBhuRJQDhvgdRGs6SBAccW1LpskvqkEVzvDrUH//60fjofA1UaIo4fqhq6M6pdtO
VlOzcxJWPrL6ULESOYDNoxEpd344ffrgkILaus5n1zsmxO9y6yzrWihyiePI7OlF
FO+09YDzRyQFyWo+1sMrdV5ZNQhHXCw3KwAkbV1q5BncAREM+9YLXmA/kz56wqBf
duNFe36CrwLcecAY16rAJ+ZAAn5W1D7vbVW/7dhTntaEtJ4LF/eJrN5RGnZGCZy+
E5VMTAkMDZ93t9UjkRDD6BCF8PW84avDgbz40Jn3D2iuLeWCWuRfVboBevz9WcEV
mwzG90njs03uGHxSpM9BXVMeTEgb4PGtWKO8WYXhh2GQbtwp7h7jJPGvTzJsxWVS
9dIPD983a+nAWtyIMqrJxedK6nEL5WHien05ViXINcKDkixEDvSXRb/atx1JiIt2
mXYNCitmtkm1gT0EJAXyvrXmVXzkQNTmp3SBGWaH/vi2ptwvO7/nqwiWgPzKai85
AaDuJakcJ/fwHXBFWGQWpSWdXesTGgQggn4f94uSOGi2jiE2cRl2ug2kgE6Fk6Q9
Fomux4ChbFv7EdvUcjtuSuJQYk+kHh6h+ofjocJgBtJWnomR2YsxCiPvfOfbWcbq
i8HqNGsvJDKBR+N9BWzGtI5KDny5koaW6sprPT4XrOUSZ4GIF2h/pDcMo+qBDWUe
TTwQNPn5z8cuYOcr1mBSOgHns8d7qW+A4clB5MfEMukop2518p1kSE3tIWXgpH4f
a+7/vrAftP4S/IqxpYm9/Zz8OF4yWqwQjUh1fqdPUZjmK24SWghbQZ8X4YhdjrFH
QcZtk5R76SiTtsZNyeE/mgMXZyxgujMBIEGE7gSHiQb00ooHTozCRubS6K4qpF3x
kLQcBkILVJcFC1uRKLOEy6uDipihwYYGQLOf2XM1V/U9Tj3dTWvlKQgFdgeDOkQe
brlszkekpWv2q3dD4Wm/uDZlg31PtXh1N2uq3TIBV9ygAdbrRPS5XLlH6EPaAmHj
FwHAbNkJcbfZC8Dgk237aiZarGk3730Hr/PfSJYrdORFofQRM/V9WwEsSGLBoYMO
TvYdssZGfx4xqc6udpac3sob0+UrXr/qzOSpxvb76b7NGurYMg9ey+GZsx54bjTI
oWJYJp6HqogDRjsLVHvEp5GQA1P33w+XS0CjVckofBb8yo3Re27YID6H3wm64M/+
GuphIKK4mGHoUnrp4K7WhM8RMGfY8zx7rGAqfDAk86Cs9lXGKd/yb2co5GO6d3sj
jKlsJB6HQZhuPIZ8YPWQVXlAWXkzZCjt3gHC9a6mv7WyGk9SfmHBP8ypuoKkc2pp
gRqrV7VcIUmt96jxfYDn/1R4kirR03M6S5YdO8EaNmYHzQ/HsX7HXYe1kCsuvWZa
aT/CaGPRZxVKqpXdKgLEcMm4pYibskKfcvKdyobiyxCkkdGt0tGRgM0aQdgv2xEV
C5TMJ9W1qy3Dih6IisZhRNd8PcTdTYcO3dB14v89RnPuEYQt9sFbwynSeKzhoqJq
J8+woRq8MOSlf4jPHpCHTqo5XxFZ8uWDp4Yh+TQgIFGjlT3mvQUz1CzabmXIwf/l
5i40hCCso6jcelu/hh6NZD6sQWiwm4PfSkKAnXldYgfWJfu8kaNNfbknT/Ztqi1c
vE5yHNFp41jASrC5SNTx7eFggUNJB1o3fJaOpNdPLjy3+pl4YmgSTJi6/pexQMHE
rx8BmYs/s8n7Sf7LL4Jh4/TSQ+2TwbpUduGLzaY60FHom3LDQXF6DfuFLkAk6+jH
1dLRfNiIaHWT89PSdK9qrN3t8NSNn70NH0fEdtDQpRKtZAUDN70Px6jgDrhQ9ZsM
HDd0pEgcYbZIRi9tI69cKs1Xvpun2Vl3JzdS+Ak067jWSF8vcykSHpJqILJht7DG
iXKgX8sJTmBen3bm8/7XJp//9R6vFo1TJcGHCoXfcwv11ZNDA4aCuyZlkVGhjxr/
qR3S65XKO90VPZjwxQNk8W5rm6v0PEKRvE5WohF0DekpjddZbLv/ti0eFFIN6Wm4
JqVgSoheb6/8GoewRN5OgocxkOdoMsv3eaHqfZ9fHjoi6XFJ5TFScefO2orSLZka
eL3ubAfrey9kb2gri8t/RTf2l8iISxRVCd9L6njlBsR4RNd9k01HpaBeOLrzSZYY
SbDHrP6zCoWgf7iji8nnIMmHPHDXp9Pbw/Jn1mXRUxobxI+S1HFng35KknmOOiTq
ElKpVbov5VCSiG9zwDBFbsym6mCJQbMr9HLRpJEBohuvI2boMKwV7XUe9t54Ok+c
zM0Y7k8jlHAVxpDWSkp/lgeESfDJxbZD3b6c/Kp4uiMY7KDERz6g7Hwi4hPMZ+K+
HxmermAdJX+L1USbmlsZiH+a08GAwyojiXEqoihhZi1QL8nffQr6pNORIq/XL2UJ
5dUlhCixpDI5nNTL3patO91cfeGyyTyK79+HV8ceNavCXA6br8IRM0J2vgBkCK6y
WGlDKUvWOzmJfZmJrPWGskDBgiuqTUUxHgMXqsBdx5fM+UVKIXi/pL36hYCPZeQE
5wnUj8EcA8n30Dv4iyvP10XfNI7RSnG3NMZh+XUCKJo51O+Jl9SaW6tVoQJpee5+
cwNKkjY6+YjZRR+qnJgWWsL8twDn50h9YjAPj9pcPGIGf2RomCCgUCO9RYMflVkK
frMD9fflnvZHdGmL6vV4rupKn/Y/rVg29lLDxq4BdEN2hmQeQc2UMMQPqWX2l7nA
wvg5p/MxvpHGNnO3od1MWJO+QqWqKT4U7fQSyq21650R+yH6px4hjBUdaC94pfkT
dYTUdTG+0xeg+3u7XpbHWkM8CRsiMM6sFeaHz0+bzeavMDMNlKfJSsoWUDyRmMpA
zKUkrspg8snA0FAmMRoPXMoIhtNZvi5xZZYcn9SesdoshbFjFiBPtdumU7RXZ9dJ
uTCkSvrPnChqY12Wczs7MELxd+AGBlp9nw0gpGdLqiLUYx9afuPfXONxbwDTNnLK
6cvXujrBlKbIGbY0WTie74sG9GchKEXebPJWNdM45a2XBJemgenW5qTUI7hzjgYG
fihIbUEkPl3rqMQEzoMYWXhu9iGPz/n3gHtFos0qy1I/VmoHCPlGBwVuYlEwlkVi
+DCJFrJZcsXk6SO3HRinHhGZEBcslrcJpKW9WfBIJJVjiAr5nKirZgNLbO41d1jf
sq9oESDNY5XTUHs4Dk0oiyI1spUwnOQ8mFXTa0bc7IRFVe7kxvbvwjkOBaANbSdM
UhCAFcoxgPeaZ31RkXGOwODqVeFXfRr9orExc7SER6sQFiF9RsYUBBk/eR7cq7bh
+Sx3SfOQrTBJ+2fQT8tmC7dxx5uwDtb2mwFOOvZWYAbx7TjUyr//s4SGKbWrRyr/
H9dj6GY/HmmusUOI5Y2ijAz2vsx3SFsxYM5J/6SYyzy8nIwlz9B7ZiUFTW18Q/TT
mfrT2E6PD9uvz2NdEVJcGbX6OsVswZZ3e7GmA1YNtyvyAA6dZIZ6zLqo6Ax/0TVg
wY2PV+kobSSMaRqwa58biS6Q5SWoEvBB9KzY/h2pLt1FLDN1x6fz/z0+9EFV30Pi
ew5WvntwwE/MNHpqYjGNO9y06G1d6U8Ys4HkAbZyEWwd8GHr02X53cA5E4yldUUI
epYzwS9BZNpaudNnfuU5fISPoumG5iTg2c8eERjbkldc88mS0xAmzAAgcm55dpk3
irLSqaZ5hFZr8eF4pE8TnKGSMgUR3D8f9wXvbu6l3hQ4kbLnkdYEl+XH2H8aecOL
zOl8mB6pKvQ9es1Rak4qrWHfVQpqprVrmAWLvq6UhhcCSjuluAeVECtKhZqDpf7d
oX0FjH+D+UoK/18+K30jYikZlMGjyX1YLq7iVApBAXXRhvXU6BK1sawq6bEOv7bq
8SfdOP4yaEJXvC9XJnLVmYwIs+8G5U9Xrq8HbusopCpvO8mdxLN61dd5nyxdjV5m
lgfCz9loa58WL4/aYn6nHqA7W072YQphKIgq7jMrkd0Af/iw51zVLfU/+KG0CSHM
j6xFa+WI56aubUcK8jNDhDTR9tfP/fvwxKCtsAtLrVyUHolzOMADddqHPRkxxWQ3
krGinIhfziGWwl7FpQMB1x2nZ4byfk927A67JH21e0Clg37HSx03Hk9K+24Ncbjp
m6EOdv4nvMDIFV1vgIPaDC6v8mC0RzuAJdAwBBj/1V5A9i+QOTLWA0X5ERM5Cy0Z
DRUdxeQgoCl9btr4Ux5EX8ctLE1rkdWtfIzPx98V2r4vwQiveDRPxzwwvOisUkoG
lHZZLRVzCMz8LRr66xDoGMcADrJahO3p45Uq5/iDkjmLFnUewSQhJLvtryzQvJfx
02eAQ1UKv37o6tMNGwpbDI6lyyS4EPcncLqdWt561fIkeQKDFvdLiih8rDWPF4Qj
YBTKDhCO7BsXvTSnSLqudb2jFDJ1wDW2GH2JjN3bLrixDC8LJiOdFCjo4c8lleW0
XTndS9hHEGdUQmF4TKpipchpoeTXbhJXPhseG+lQS5pcU5XKQMZ6DE4b7OiK5WE3
dXqqzgGEs/uE8y9nh2s47gvz/U6i7g2KBGq0OqMXED1yqf6OKsIkAhUk6viHjdpO
aGDrDDcysTntDU5rR2jDrAFLb6Qq4VsI3mezLmEaJoKWG2QAnrn9K7+gwHZlp5c3
gXNyULIhes2+/bbAPV8cRvCo0AO1yDzVkubl9fDDkpQjQOKgWne/pvWR6n3EJS4q
HzqGWsoCWRrJt5Go6eopfGuAr2EOWWfFmsLk+FOBACyLVtmLYqk6uYMHYXW8pmz2
u/sQbv5SQcseuBARqwK5qU2S0lw0KcFBAt63w478/+6At3iPWGsrYfNN3lXNMd5h
NM3LlOTZZaFHH7JT3IKg+X1UinQTV3GoNkNfZPCRr+/IQ7rhWoWIKn90F3e4laiU
v5DxiG8PzaiH354dwkmLusr7dunBoXmZ+QBrn13nJFgKpti0CLwuhv0Pi9wWNIyl
UpA/qXwLuioZBEo/ZzWb77a0jD5yoqTO15QoSc9iNiTqkqBsO3p+Q+IrZgtz0AY+
/D/QFaM0FqYNRboQbjx8PJm2pooYQwryN3stkE5dlLO4M02fbiXEXK9m/0QqO0xT
WvshijcrMUt4bidOnm1e6i/UIy9NqsLcn3gxj5TeXYfshPIsXhgqxSl/dBJqOtPT
UY2jjRdqAlxse5UKrLX+jbm75rtzRdfNII4Llp/3ab57a4bAdb9IAfaQE/PLdJ1a
DE3gGmHTtccxkhrRhKBC+05kzgAOZKrQMDPWQcBBrZDzxbzNIEHEL7ZdL61eldoY
kLgKw/uZiWdVSlabICh8WBunDKIYreGgfLCN0SSZ8na4bask9tEp1QmPQtJMQzRv
HGZRB+xr5l7oStBE/xonKqf1U+0eJacUhhabcst/wGYtF14B8KQ8AxDENvvpdy4x
OadKSEmbvHVjrmUVpbZ3OXCHurSfHxrAh1iGOwdPnTRvmQSH4M+LOunsyOdOlRZa
fjB9d6LfcH97sEoFIFUdBpuq9Wep0/QOuiinKcg9/WuMGsyZ7iUR5dzvGCLi2IO1
q2nSn5S26D5HqW6OT8Uy4ncl1l3eK/o4gjZ7Et5qGCZFZVYnUxuHFl//cS7y4qh4
F+QSydOdG8i+c5MSEWI0eBvKnoxm0vqefVBw9aPHEHqjtM7JkGwCAgDO/4SKhRB8
XFn5DGCHT78nOv7IdCa5FUM8HyblMOc4buG+YHa6MdUkWbldhrULTKJ8ykpCZv7O
SYU8Js72Ez1c6RuO7Mxle+ohQxtCoEhDGSHfYKtvV5v/vC+7apcMBkzQ3K9xxjyZ
dlnMqLPCeQMGYeeNxH2vqfKW/YGI4JHAAdYUDVZ9IyalN5cTCOZTWP312vBRKpqw
H1z2OMkH9zbqh0csNas2Ngn3zHDn4rk4ZYjWgFQiYRL/qwMV9NwbkJqQ5c1Wk/q/
ILB42G4NRDWGEfDQIu7T4K/88wF4+1FSgXg5NLkofd0n9GR2L1nThQCnQosou5Gy
yqw3hhoS105TiiTNbrt1wg2WkMrGXRzEL9hrDBVLh6XgHXGmDW/rm/U+Xic5uRGs
719TizPqBFYG1dIrVLakWERcZYxcsmAE3DVcUAlDxK4JwcJCDpCT1nR2VHHH7AKo
tprIYE5+/6eoHlPx7f7/5gc4DClIlHozrVFYykyFn5b17cLcF1M/XcIDS1iYwvkC
0zmSBr3REKMq+fkV07gwte8uFs7tb7G8rQbwwagedVL3rupqPJ7dEJqKKqePPa6l
V3E6MuGsPrK7UZfIzuh39Z28Qfh0bRI6Sf/ZdljUmvTlKC+ZW69yAYYdGK+u8RPd
K9XY47SKKpsT563xdSkLm7Ww5sBrzEPvFMuxdE48UoJgTza0A7hp6E0cW/JK1wZ3
BRkWg2oH6gpLe6jlovGoQHx2tPovK65NLnB4AAB/3tyaQQLPNUv9eHccorhOpUk+
jzZgd0K6lrgeMnIwxrSJrb3DSmaGXxfP92cHucbYXK3yK6PEVE7c1gabmT+5Ozju
bS1uS5SOXjem0+nrkhPFMv327obSPNXr1b7lIXtpFCmKzOKSZvbPi3aIjzfg0GG0
gUX9gOh1zuHfPXeaWxleh5ie7Tm98ZiZLeZSPIc18u9kW4cXscXORU+Qh9osxym2
Y5s0evbGOKVE9zq/TMorPUYe9DbL4WPV0rBlRgVBYxPrdFZrndNWW7xCxjZ2SP6l
V268YkhvS/QJ3DZQDdber+BM/icjHplxfaYHEz/wdjKzxYH9aVYXb0Gv+5+HXVbg
hwLWE0/Fs9Q4T7FJxz29Gs/M6VEQF7Y5ranNSoctYfRrtz5NcKtn/VrnXow2pHtm
LfYlfJ47GawwoTcaOyhY1Fb+Nzt+hqCBi/WbLPc/R5H8wTo9WvyDiOV0jlGwLPxO
wBS9aO9pNKbGUT7e+ApYMKzIsirU9BPAq2Fd//KSav/6viU6AfZNSRlSLvb226dN
5jmGdTV/y/YsTDCqxXklshV86xpEZbTLomndqTRTlaBYpIziFZjpaZyigR/k3/Go
XBdfTiHuSrJOxmx4MgHrN8ZafGG29FgqEl+7AgxawoGPymlc3+upcbVb4x0yUf/0
UvKFLgws97GFBMYLeOHWeW/5sIy6XyR86xUnW8cH+RR/p33oapc29VYQZ+Aoipni
vd2kkaC1QiDAIlTRcZZrBpnm7CrVoUiTZE5GB6VJ/3GPOL1gx/Gizi5j4CbQAVef
uHVY7hCeMgROlfbd7X3ANEjh0cNfotBa/xd8tCbcrQIKyiTVIILtHjRO1HrQQwRJ
x4mtwnOgk/enJySfljlxRbTuKUbOoqPh7rkim/UaFPlQ2LQ9bO9It+6gOdEuSHFR
h0RjKcruHtsumUd3vS01NfHd8j2xiqEMSTG6q8QePZx24ezkrPnK2ZgDzyu4oujO
0Xb68NE32542SaboR5Oo+NevviC2oySULN+wIe088/vkDKbIk6M0CZ1SCxLjvhN+
9tlczQAcIEXPO6rpYyH3rhs39p17FOZLlx63DgsWD7YplZL2ptGs4+gFrmZY7oTk
vbUEtMcAm3UzFboGPAUY2WOUhoXUDxc2HIztX9yWNFCQIPdvCpsdkn1HKEqKjGGC
mXFe+F0ZIo2yfSlif+j3/30KokN3PXG/6j4MvMEyNo22oG1GYTSAllQG1g8n+Rga
5XSiQxk3FZAEKGX566c2YpJ/gCQsXZElvI21uED45fDPsjmk3HtJP19EAZq5K8NK
0Lju69TwF5mCc5DuB0/+/pvC9EuTlaDBLdU0CAl/XCTuKkr8pglae8tGgGJpwx3a
BBs3QQ1+bF3J0mW5Gp4O5ZDYTqHIA50qIl7JXqO8qBWJCeWvAIr2ut/PVOx0Zzs9
I2TjvPwK68Ms8nTk6/mxGo4vR9QrMJB2FsvFo+CpwXR2DSXNTNLz/9nD3XN/PdTq
zlyrh/LlbIs1c9ObLGA3qtxO6JYYwNOj144UpdLOzfwsCfY49kEq/01pEl7ja7PY
rEx0692wLTgaUIa0M8Xlb7+bEFy3NuLNE6vDFHNXUEDlj89lkOhf09AZYpLfFIJL
bxgusRjMFouKGl8FlM9OE6Ggo1ACsrc0r3ZeEU4VXCGY9Wyjos8t0hKiOePOA94w
u0n2XbkRAQhDyQHHolALsVJMk+ayiKHksnd6urCzTwYfUxBbtUp2QihyTlcUi+xw
l4VQkAXtGe/FElqjXGUInzEdeOxuynjStAemWirMaLrvyeTtAWK575dx5f95XHoX
o1k8TZCB/s/gIHQNXEANZiUeyESQ4nZNgXHprqk1VEBeO9NRfW/7tpNic//wF9jE
+WWXFcNjtObBVaGNB5co9pU6skR+mGtbvHKLFRUyvunzLOJHjYdrP5201MbwAuFc
b+u37eTfiBXLneyjLa9jB13dd28nEaGhtIS2x1zG9nyuyx9LYOxLO3y54bvCm8eA
uZ00U8ORLGd4ZG7bNCnJ/+vKNj7JkSp2kCD8hWoypuTjgOnZiv2fRnBri37fL5F/
kfY/z/YYxSowp6UoWhFQ8v1kUnchPNEN5knoc7oxpicMe6i2CgAfPt54OVvL0nFK
7QBafDYlru3yEMimMq5vtQmoQhNddg/Rv17al0cbnRjY7wmGpCtF6iAQihzg7RkA
ouhYnidP7Tu+nczGq0phIlgeVdjOngWy7zKPxFKfRdlvFOchly/JYUZrfTynvUSA
ehoXddyEDhsGbF+u11ZPSyvmjr009uLTdq9x8FVzrbDf1/liptQh5qc05g9PA0Ps
/B/SDsk4ymylrX+pKqC7uIzZZxItw6CsLnRx9Ca2iyolx3EEfZbQTW4yE4Yy0QOa
vso1uB3s/2WUt1eIRA6nzVZaLiY4fv/+2Y15wX2A/no6J4Z5SKVYqRgvwU8C+AXz
m7Y5pI9MTGqt3hy/BrQ0b0+TR+soP8rQG+/4bIWzTo47ylTlxTCnaWgL/qZFPEZX
AU/RSTHHtiaMbUfFadZhPNk6FdKAUYe/EA6cL/JZrqdCKqNypiGTIfe07s6vuEqM
VrjSSF9Rx2p9bs4orVivx7VuGdUw8QowK5s2ny2242ra6dOCaQ1ngTVU2DRbvTyq
zV5U7keQ01pYPowtH+wYWH05M7mpqtsysAfXZ7dPCbW87wSHhju1tfu10RFHMFZI
wK/Hl8LX9XHgxPlxHw31dCLXykDio0Noi2BIIFC++V9Xt4FE3CkyulISyo79mVrG
xAH4kWaeo+yxNf3DP84Sj/f8baRoTgDGXmEjSydPPhAIosXb+7SmWjVpm3CH1eoa
Wrz7uKCeijEGEsZ4IV0IbavY24TOB3t6rpdoBO1bSPkAqtJ0PqVn0u+CUSbJuzbA
+gBFhILXDF3agnCozPG7gND5butn7RsVVk+TMQ+QR65wTpEvKJVE2jeaixzp42CH
OUQrxMX+nwWfvXSVxPg6sT60EJne00Pyp+zQr5vSVsGHburGYfwWTkSf3VcdPMVm
VQS6IyjoYZJf4sosRdqRMIgB56MgO2UEEtlh4kc0e7iU9DJpvJ5SPbMffzbGBwFV
wmLdEQSR7EOB7s5aDqe/PwXwSKl9a+1oOELRJzPc7GJizWTv1lBlJicInTlRQ8Oy
rbeBAGDPy98F4tLOHcS9+hm5TouAr5xnm81X0UQoFL9MisjeUB27QfMtetxyVd/b
tSmXhV3f9apVdp5Jpr/bTphKajg6w23UsYh9hER6gZFnC797qs3dLaTJMhuHrrK4
g/dNM80R/t3v8f7e4gcjKL4d5j/tKPAUntXCt+fKOKw3d2s8l/Rn+mikFwa4KxL7
55sBrqtYLRqURNE1sjvn1+X38Htz+tFTXa3P8VrqjlQ9/X0vdR4gh+22BcT6807C
mfrw7mpxue2g/DH7NR9f2aRj6rFbVeqLaYP6Afih3jDHENl3/51z1W/2gnGTCOqA
609zGlfoytMdg1SDR0wxzBwx52BhT1/sz7KRvaVlyOuRI7FaOSIpEmDnjlJ9rxlq
8jwxoMQyebjuK+cicZ7mzoI1k4x8jEF2d4eta+myc/o66cV7DLRkr+3tli0fV3bl
e4NT5cGe0PtbK+9qnzcESa5cmKZmUaFqkjI4pza8Ru+hCeEb2/MqPKYw56HrhTQx
NTuGEhB7O9eN1t2CC4Mr6ctVtBUvR7ZE95cu1h5NHwINegs4qSwBIbSltUJqtrqP
IOYaQZ/AkF6MogYPGb9jg8usi7eP4AlWmp6CC5+42TqQ8SHky61kjlE6okF+z0hD
1H9RR3zHa+FaqizPHRrORQeUQ2OsiUmspGBpYy6o1DGd+gbIybfXdDaS1nRjlfbb
WVO0zUOlG2XGP4PZDG0vqkltDndT1UZKpJyGNA7EXfhQTc3Q3RfufcqdnnWp+2Pg
CaujEgZxlQO6JjGKEvkGtd3JiQikok87ao/7bH7y1qbPSh6FMsA06Kydbs9ER5rP
4AyZ0kukXrWocFgxJmL5g4Fn7bMgtB8qE3e/6XQIhPxQoM/eReA6EAY2XtBnuoX3
OWDmO4NJ8vLbFjKW4/a21GbZoBRufZmfem6UXv+UHgBRdAsI5iy8m4IqEmrDfkW/
n0seanCRTMtc2/EdIkqOmG7d8fFxlBTFgvG3/EELf7cmbGxQlFgTpFI1ce6RDpNm
t8ivgoZF1/JATW/kUZ51T/nxetsZFBrIMG7ohvcWHfngC7mX/RuxHmIOhJxApta1
5sC+ESBFDkRrG+SphdD3jU8e0INQQAKCQ8cXZvYtq9hq48W3FCb5nu19cI3aj9du
ob+NHT67BdQvID5Q+NagrplFGrgBczqQ1nrkfnZs3E1AXWFSGqerc4R/8D+VPB+Q
stMWs6NPtfFLhKhyz/dsC4BGRcgbV2/sC5VBwlmOJVMNihSYMoXw5lFJKgtH0MEZ
sMq88Au2LO9204M9x51DkCk4PmYj7MDES+wI2QS/bDMKaK49ESvaEV0Q7Frd3P+4
Ian+DabtZGG/82PPWFH9W0twzXPe2OS2+DB15jpX7C3W0CDhXicD64nO4zYHoMN1
eljZpG9JfdRcvWnoE47aTnCVbEKKe61r1umXoot/YxOza/OFqgWE/coOnn1tuW2L
KCMx47atIhYdOf3udf40jyJypwP/0a8AdHtJJrEb2H/vcK9Zq+/psBYteFxjiQ14
7r3i2UIsjItAUu+aBUa3DOgEQpKjxuOYgsmTnLYYctXLVf5dSmCx25fa6pNgXSM6
V9Ec/Nyi9BUY8VBlhw35lsXvkcilZ4dwMbyT2i77GTHZh+Gbbahf4ap/OdEiQ9iC
PEkYlaOdLwHBSj7ERDoSFd3HEEgf3sCnit6coHj3avjWQI7E8bP/EwsHdmQAEnHz
OeIRi7n7HjBaBLqR3LxOdEhmt//FwG4L97CAhggTrq2xGK0zjzvWlVdTMNWJMgxg
Dutsc8GPPxSDqHyfUq6QloNecvoH9MM6AVbvi43xUI8fMFQ5lUFvdCcTX06m6Mn8
6YRCgpgBumibDCpc34ZEvKrBUYOuw0bILcFYz8TxygjfLE2w5DmPsEuEhvhkPnts
jP236LreEE9TBVsKkp2Fqa/ssDDjFtjtio26pozvD+F7upSCH3mhcnwrLQxbRUzI
XzO/v1bVf0FaJvJgeQ7+y48rG1fj8ZtorT0eT/n/XXTAGKg/kJ3625IqOoVN4cNq
TJH1y5hwlXTHnUYlMTiOBI1bJr9FAsMJn9DBy3EOrZzuLsK7o+u4bmE6oDg7F5ff
NzVrZ7OTolx5tf13ZcLoaFGZ6Ouy+N8kOV4rs95Rt78Z07S2hSZSP77SxVirRCwl
aPX8ol4+5MjDpt2W0fLi3UrgKkKAinIBWKNrDm/5vlz/S7O9MR2demK4Yk2D+lKD
vMtk6baecl0bsitErsbqlIEBIvNAyAmdi3L1Wu2OAIbfftleVDunpGeq7jYqTsf1
15fmNhI9iEqVSTOCj7bcEB2VKnqVPLt2Bh82XT9BfNkVGypsjCRgGqsO1enkRJ6P
NPQVT3c0QXJGuKfG6u8CUnF5YA3CHq6AhBfki7fSIImIFr+JMhN6Nv3ha6SBQCnG
kjnV88uiA8W6PT3x+Y45GtOnUh29D9F/sX51jlNgBknYf4F96o3qJPvP/YSL3DdT
aX1GC9ksCGcdax8VuSnngpV06RlFqMcuYyuUdIx+0tJjzgeGmw8/5bQNw5zenbAv
D5yZV5yCagBgxfdsAS1AqgVOZsKmX9FRozyqUGgerMUOzcGY7xcd5GniPXZr4w5H
XE4JKx1oTxY89vgzZHOCN5ZGELuu1Z1FMPE6e20rcOLNbO/kf6nRQx2mNvwj1SYB
Zz/QgfsaANuO+qFZQAhN36Qrt4x4YBGQcOn+RUWjqBxdBf9w3aagULmFEiVrnIyG
qx0KhTAmHJTMhSO3nkEo0toKSdVaQuHWOLbaNz9HoFUrDOfp46czwqIZHk7rRkRl
R/3ljssWXXUGB3FDNCa4HVz3TYcawHncmty6JRlt4DE/yNAQhmmhBtn4SDDe0xLK
dJQr0QMRDbiMy1dPdNpIYAoVsMINyKZFf67IF4WwKP0aSFzDN8DyfSn0N1K4+9l4
AlCKtpoOa7RjDek3MnJaC50xNWLzkdRriUgCa0uHmoZTUQ/C9+bvu0bddcamGui7
RyU+cE6fdD23Iq6glEvB0WAUZNJfjJ8X+GlJOcP+22ZG7dDBAEy3LhwvwHex17ug
Nqls15wm8oAdiZ4Xq2l0QsL9ha7Resv7rX7VC8dJw9JrNNG+B434DsORxzNrG8Y+
8tDZdPw4kJt1S0WJtwOjFIgateZ3mTgmXQZ2CacNXHgDalt+zZKjrMLZfZ9QpBTx
ooJ7k9mllt5DJmlv1f518YhT6+kbbo2lpLWlZ3i/TAWkobibIFn9J/inlQ0pxXDE
ohNLDXedqKMCJWNj4nwA7kYK4tHEb3sFeTQMtKlcxjceSFmp2IzqGlVq/tQWBjlL
N2KMTvpwuU88O3qf434Z9kS3uVmdzAWr2R3426eB/B/eTnzN7TH2+G/uJDV8Q36R
qYkGVUO9paHSzdYMdsgr4H9n3cVIXSfX57nkZ247PylBl+xmnb2L6vwmiGDyOVvN
U9mcaB51cOJ11ApZEfLNQRP9Sro39EDqvsM0+nbcCBuYELVKd7HNBDf2o56Q+1LX
mwWK2YpecDHKPgywyx6Q93ORi/Od1rdWhxOkPxDXhBIbbEB27gM+Gaw29pgQ9pXJ
kkdQuTiXiuk9qIkN33gmQmUbQuUtBuwu70UE1cMb9M4mORPl4BULqvJpflB21OGl
2Wpc2uro2nujwhLtcDX8BwlUBZdiGjWJo/sp/MfHltYCs1aXYEEvxSqPU3A+864W
X22ZjYX7o1c3wj0mVZi34osTNILj1XcW1ZYRgvneEXoI1N/KCSTFE7G/T6w8ktT5
mppIOCzQ2fH67nWEVSGppggPFHTkZb6Fk4pAXKLmcvaxk0iPCrThNVUm/Tz5fJjX
0YvT6lnIwvlRvsy9PX1TzolkTrzYnEnLzHNSpEF9IZnNB7BIEQU2C81+46tEKOzN
wxOFyL9X0ksicmZt8wUzWqfWKvH2tYsTmieD+0X5awWb0ElWfIsCTX++pSISwPxH
nNezQtkEZM29Qz76DuKYf3JxtuywA0mIKD9McTQ0F0HN4Rw8W8uMjZB1aJS9JN4G
tTzziRNRUT6zYxk+tTOotiknSejqI0UtDpqD24bGoxc=
`pragma protect end_protected
