// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 03:56:38 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
F+rUBpFIGQeD6ZP1+lFiPuxb1C+EPcXzy2eduvToti2uQAckVUk4p+pFumvywwQL
n3YbwvuG8ZUDtYmc2N+Oyyc8pJMJO+FXXdVzWYwoxOmhTYJ4d1kvbtdeQgJ30pyp
H87BlrYkvOdahWO64gVVrAh6r3TbPN3wpOCnH+kHSfw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 33696)
xFW49l9TfibP/CCE8I0a7LJ3BiImp0xve3+N10BY/Glrl1CCbPSBn6M4JZsvTGiA
aDfd7YtHi4UZ23+Q+IfUKjlkg/oQfnL14ijUfaGRm00ZBHlaqvyPSf3R5cHiUuSf
m41sJ1nbcZVBHSilBV3BFf56T5nKtW41363auDpiK3DDUNqREZElUB/ROUkqSeN5
FjoSJEZ3WJWI1DP3TdA4JuVM9Yqp2o1ol44+2odOF7TIxEYzJcRgs8e06FEK4cff
I5j2LT51eUhMjgGBF4m8FE4Mq9DxCDPL0sKQwgng1aFPq9ACDx/QvC1jvbbu0Qck
xJ5kooSxhTgStpIlSw9G7y9z6X47ncLuFGd3HSZ1HO+xBPVruYBNQo4w0DFXVMej
0DKmILU9UkR8oQk+N3EVLOXf2wHvnDhkY/K7OfVxQAO5/0Zv4NfmlhnE3c063Jbl
nWb8oFOyAdY2CD5JhjmZ1TrYTd7KektUICzgCZTg+M6wK8tx8shncJ7PqaiAJGkH
jV+gqwYLE3hOjowYW/QGwW5A+8opZb1KEY+5TnSk5yKmYu8GSA/OGVy8Jya4xdKt
MDQkJbTQX6FFPfAjgzLTFmSsoNOvdZd2AZ540ldZbLoLVWDkQXxvaUWZEsLBa3xw
2SqixIRNpWRdHidptefwpfxtsmRmG/2Dc9/03ZC7iTbmJ7Z92SZYAT6l/ZjTlvVu
UdIi5zozUzBGuMqkmqVl07DM5lK7iSNJuhxMGe+RJgQxrLBf4WzS0WCnT1yUPInx
e6A3lcVamJznGrWhLKAi2bgR6v3z4AC3cmPsxkgDuku+6WhP2Vv4qNHwAhm3xFTD
Y9Mkfcd6VPmvbU0b9DRLgTkfN6l9o0BO7BQkDXip//FshHNUdFoGKGCUmLWh5r1V
DCmexyyi9nCrrYk4/d9cj+UjLfS2L2ScQ+OlteUzaDAUrQnS/KzNcpt29aIl97b2
bStsZRE0LZoo08y5P4ndb6LV0dAdolzty7/fTkgiWiFdwcneoZWVtnIyQBTDnkAc
nkgZPPBQlJR31CRkNQ+pi3wPFq+l7x+UyzavGUx6NpVY9ss6R8sVWF7O+egvzHp8
eXFgoSLv+5fZULhjg+aWMGHaBJpHV5S4XUC5uyCVG1wVWcSZUQSxOGkiStTUy6K/
wGzhZ0aRQwS/B2igiEUzGzx7v9BD/8RTJwUd0iuWlJ1W+Jm9Gh3+pIy/NXkfFt3p
kzAv83thm2TVIGEHLh+2652Q18CFLosvKxHtJqXACHKB7QJpPiSr9Oscn8BPF22F
sSBhpp7n5Oo3ALseIO+Qy4aJ+RvVn6GXNaASLxslq57KCveOD4V5z9VJeSk3A/+p
laaThfxEsJJqaAqc8XBaRTfh9fN56/GEWm27sfhPMiHECm918xhJHhNgL5MyEEYL
oiWPXPp347eaoxyzvF2svXpMncQPDk9eVcxDkqire16UcxmJkYL4B9UXnSw5b4IR
o9upemITpda6Ht+2ywdt4UU4O6nZW2hcZy6dEyzlTGgipq85pfxVx87jIjoiUxYF
x10qzhgAQY3nkpPueiIZQUBv4VVS6tt0rYRifOe8lOQ6yrlbi3GMre4PjgUtHrF3
C+6+K/aKyq/4PDahDKJGGbjgRpyjwqmBx+tcwobOHdQjWvvyLY89eNYK/bRiYzwE
Ks9mWvDAVnDemfH1f7W+31kHET/v8B/8d7PUTuodIufOyeyLGYalZuBury0aKCoz
g/peWNOp+bEHJMxI1ZDooQ8acDi1k8joPSodSDgbM1uispr5+rO7i24eC7uAHpIx
JBEOyWveNwU3IZA+Ci6kYWlujnNae29i2YjGLPiSW9H9kCqpYZmEXof54KrnRQ9l
idv1Sn074PbQQveU7Lp9x3jTmOKeIuZ+b+6AinEEq+Xmq69+sNcbWBosyCbcGFyu
x77P3WlnhiBTeqeCTUns4LynyhZCvZi59ohSSoSDYgVQpGR7+WwthtRtjhnmPLoG
YMztkSsiLJVsfITXIOk5lKIlsln5oRhPQecJ6D2IdFYs4DE/dlyjb2VI8zSumF8g
fTZeE0a6fFQKZ9srkZ01pFy12I04YqwCriLd5PlTB0q6VL1Dc53sKBGX2dF/YWFR
kdBaF1cYclPLBIIHBW1SxWEu4n6nQvR2Hf3PTopk7G1uqGeLF3Q7QaSKgiHfpZzO
0GL5tNPpUVPMO3PV3dS19Act7opYJOHLBEWbSu3SjExvK5vNKbjyWRda4yAHzOj1
7dV2XjCTyE0//x/055W3U9kDJLxBnL+2pDZKtTQoy+7ezSfL/2wME0+8oVymn+GC
+bPvQbus56Da2J9HBgbBK1gNh3gxAmOyv8mL/1mohPLXwShUqMIsiGNgNSo7ButP
D+lVb5ndCwbuuvymQ/2QYroH7+zLacUZas+oz6GdvsUn8K6uNubLLj94gESL3+JK
6St9h5s8UsRlEGGuNAK60KqpAgFwvVhvsQgmpTteAgFhxtt24KCUiWNnS+MK3qls
BfutzGZQIT75R4U6YOjVU3nDPKDc4Nmd05xxrFAPy1tb1LWz1BWCL26K2vVGBbe5
rxijophdqIt85dZeOJN2NKrNqxjSlSs2fsoekHd/MHfRr50rAiEqkIS74Kf1siCz
acMW4/ACcI7/n5xMwQnHYa2vuufbRQNrpIZSC0xLayzYqsE5225+Pkq93rAf69gF
XPKVuLOxOREtMrMAXugKhXOidhVvxx4nLFRUejXPD8beNnc3K0Ay4y6QguqCZa0z
bvM41WpifXqz/4qoN1C6/rYUaWE8YnlWm0FqjIdCNR9h7kOgbS28+lopcSeE6cBT
+uyTvvGa7NCohvXiwRNcwglYhhh8uHpdVqwcmks1aG74rCAG2DJj8Fe7gdL4LRwA
Lxr++lzfronULpQ21/TtARLJVVLXJV4A542v78fZHEPfkol45Fd1iN3qHIqUOfHi
ZHgvrqkV/6LdWq502o2jOCYY0v9myRDa+uncBo8kBetPnHFFoKu50P/kkJFw6lNa
DJ4sfpLYzLHDXiLUM2PCKPkaNIrSiBs/cE3k7Hk3lwY1r5QH+SfK+T7lewyj4sVY
ZNWPB3mlvRNY09lxtiSBg+8Rvo7cHx8cxB8/qbGad8j9CGJmaGmIxtoX631jQmp+
TU02fyKiMxS7rw1gUfNbv4C1p3WDDuw4FE7uVHAEvvh0AV0itoezXVTcAC7dCRZP
e1oxlNThrxuZYxt0KgVQrEiSSsTo1q8Qu8F86MlVHYubAcJpN6mnX6LivUbPSXhr
LCIAbc/F9SwHgzrtc79ZnDiqSSYAzgKIVaDameZiTABSxT07XZdA43orbric8hnP
f23P09R0cGrAy0tMdIHs5pGK10QVKwO3x42iagE2+MxFG9+3zSl0SbbPx2Oog9Np
ZBRgU6npntXcYblrE9Ts1inQiSUZrLlDmtP7AILtxwLnbf0EbvRAdnGWJ+Psfbxy
9Zox0ZULn8NIDkejjidmq5dkVyjqqScgGMQjUm/+ZkCp8qH4gpGhkVopMCGKho4J
ToQoy9DmJ/aje+9ESBSQuPmzSM/fw4Cy+3usAR4NtTfOEmSUpVH0Z+wsaItXcxln
R368Ii4waf0jNgzerVYvnYQZvwATkCBFP9b07N0TOIQoSZTMOgH4VynH9rWZ4J5h
pKU8LzaqYFveNSIXHc07h0cUEoQQ37kPsKgZC6Dvgl35amdz0E+eiiYTIG+M5bwW
xhOa2Lox7PhlagPuTiiDKh/8IyzRpV3W8EtV9ebdjpXE+9ryx3VP/EtF6Z75aWyd
HRjyWl5oB8FR4UP0yTSLSx7zs6EH+pDxQe5EPyfyUFXTIlde+nZhUK84i5w5Yalp
V9X0A9gXzIuaW/9dnJwsPrvRPtscQ3v0572VXRflUo8ywEbieH/BIM17eeKdWHbR
NpXef2Ae0cStZxYbQZ/sPNrmiciSi5y8DfDkLU3AFoLVzaP67jwgNKyntnz3jDQe
w1sMzrKFHAB5haH9YOEypobBptn3kYmsjCCxWpjkkemV/rsd8gteK6QlP6l8wvmH
ry8mup/VrPoqBw9H0SjxLUh7yRGOII4r+CXA2zfnEtUMBHfTbpgV6XIgwksmXmF+
0nIB1+CjahnRlGX8X+fnAdAtVxmtieJ5BdI+IAfbYhNsmv1DFfIFbXfGqZ1wze56
aXyyglaONnWpt3P2gezTPUKI/w018Eq56dP402n/S9Wh1ILkNwhIRTEam7LJzFv9
1Wqg2/jReHTTNftBm4qNIWu6m4hbDYxgP4tBEfHKwKuGY/zj5leyq9SnDgJWM/an
rQTniaSUgJ99nJdk2At40CH4BjvAwCWZ+jnEt/52ls0zs0hIc1urrIS1DMtCt9yW
YslJM5UsFldWTuJCZyurd5V70zgVCHNA8WFhiekkD9uh9e/uilNyUZLti3QUln5n
rvRsmEv2a6GqH6ooA7ysKwU5h1z3CySKaXSA3mRbpRKxA/eouIShJ4L28v5IGOgY
3Uf+jQITtHTlUzQSwJAEK6+ewKv85ORhvt6aaXL3Z2WRgVUrVAGrLXXDtTs9/TM4
JPbhJDnYP9B3Nor7dap9a9nPd4DOmwUmFPDtmm3N+Ad73BT0HvlTG9As4fIdoyTy
jDWnyJKbovl8XkKZM3l6oYxEh4/SsEXbf3Yb3ZwrBu0SsKs7gU8Tnrdz2/hm58Wg
+J9QhsvZBgKkk3j2cP6KGACDdoyrRSaJuqQlUZUpe3Ty0lll2f+iCK1Nc7HZS9JS
HPrJmnSIQCaoahRD9gQGqzIVzdeUlVgn9mx/X+bNwA3k9YptVB4hVSCLaKc8JVzI
anNSuZ8p9AkvVPVWWROBbD0DGqq1ExbdOGizgmLCrOl/s18F1nDLyyXSYEgyD8AO
8Otfxp+5LKTPOll+S1Vh9LkPufAs+p6d9Az+BR+dcF7tXx9PFyVg3hn7Klnqt0L+
+rgbYAQc+yNF7dBgkS033BGDW5ARAHisXzPTu6dQh10NzyhS+CkZADVhAuzbNHWR
lC3Go7oHYCcQN8Pq+pUS/+/3K0cy1lAM/kMxjTvkU9LGxbdn3oFZxhSWWJZIA5tp
ReTXkDXFfaOigunuf2O+ZIGwgjLfpDtwS6crvEjcX7wsmEtepM90LX4XcKIxAkL/
eNy7Fu2SI2WBLXmc8+7XhQJzpi6Nz9P9UaK4s69n6CgCP+cD6Yjk82oD1eiI7f8p
6ucEF3wOdgK6Nh+di49SYSjnrxha+xrt5WL+8Pn6UTRP+7aVGCN8I5VOBYl5a0Db
HL74gzb/vp8s+xMHIRNHy3g0SFUn97ygljy44PV8sa1OX4jZOoC3mdApP1AqaYT9
qM8eenRuRVMrtLzoaMa0mF4nqMSvoc8n/5NDzAg9QbCGKbscdSXFHLaiViyiuPW4
NwbRhuf/1d0MFw2F0nFaQCbS90zTli2qfYRjIh/OT6F6N4AasSy4A1IC5rAKqRBX
HC8qNZ7ViGnM+SQzTa43TglLtfborlZ6Z3uxxXLlH6RwcddnG1claIHOitj6qpLX
ZAVigzYZcwTbo2VjdaY1dV01OH/QCfx2L7CE/F25dY78wsfoPNJpGarHvVxgLy+L
4ZseJBohMjOLi1Gt9JrmA5KkqotFSHE/SYa+Atwda8h4J7XDx28U+twJNIqEs4Jd
bYIXe3WHvjTJb1MS0uL/TxLM3DDi7xwVU/OKqhK3y+mnRzY4o7GrLUzTPqm+wtAo
XVVibgEvx+TlyTlfgazFd21fkXFZvFV8XUp9KjN/2Uinc5hFT0WCjHKd4aFZBBwv
K+vNk2BZjUEgSSzrpiHNC/jAFPxkEqX8qWIskXExhuX9Gg20pjkWzMWrA0aLQfY4
86Lzbs0koBVy8Yibim8NvvUVLT0EHwM8pGOZTXquqoDrDtZD8XLT5+svKXd+YIZO
OJmmfyQFjED8iDhcRdETB45kkwtMBs7YcVAUkmo+vr1QFdXcIF0ciCSuaMoTqSqn
7WplravQm0F2xBFNfjQFtCGpo+vdDwlz3Rj5qAHLo8OZvW4dsM7H+faw5/ji6Anp
5Yr0gzXUKtQwOOPqLEebt2VmkQPU9sb7+OpqdHgeyEPTdtigYhhu2fPY0wBIBaiM
yUI9Mc2i3ldaoQG9jHdGejawW1R7WxaM3V6Cxs82DLj2Nlgrrhwsjxmxv2blQoAD
na6qJV0tTdesbDOFvzrlh+3NDprEusGy4RLVHpurkyPt1jRLt7yCHy1ORnkT1uF5
e44KJcWe/BgCcdlvvl2FMjQ0S6nSQJ0G/rYCx/WCcwVoGGVIH9eWFK7pEMVxZKHv
pgHg9NRgD6xBS8UL9K1YM+OZiq7giTCbf8pS0ylwfA28WiPZv0R5axz4x6R6dH89
i3lrffHvQ66sgfZG4Qd2VPWbL+Cfv07roxSAT6z4QtHkpdstSJ22+jt5aRNvpy8e
1bHoRwZ52tOex8IwT5b3Y9woNFb70WRig/Xm4XYz34FZH9BodRBmga8RN79Md8Rr
+gxC9InPMv0dyg+Z1D5mWxSdAoNH0W8oZBYxvxYkAC13NQTY0mGPR4XDbfE67ckk
vqdepjjl3jDRBkqK5wMwJdDb0H9b4AoEj91mul5dhQemD4ELCPV6vmcdxaWVcVI/
WsgW/sfQx7u61O5xj/FZSfOfcCIBM9V5EFwClyIUJWWtTVH54PkyYIDtfw1XLgeG
3xI5PWrnS05zBtQFtXAmQcNzeRka90W6ad+vS4JajUMCBfehtRa6KCBKHtq/Gj3V
u8QBs0eBax7c+sL2D3GZt4WAOxCjtobZ0c7g1xoTnholTioLHHzZ1Ssy4ClbTF8b
2ba/ab0qIARaBV9azz6LNvfsTcIFi0GGRzGvyX7VsEW5PeanrWlKZbT9ZQAvI6nX
Yz8tRwV1hkQPj2am4priOJws9NtHvRstDZSwQeoIViL6uHgAqmmNDTJiFl46nL9g
C6OOC1Wh4h2DtM9fMkHA8/ApHMC6R6hXEd3VPDtmKre/ucdhodH2kjAzckphSV9A
SH8kDwKYjYDfo0MRHLmgI3t0lEsvvDBJThmF0vIrpkWul0MD6SpKf+L3AYHu60rA
90D7s1lq07FAQAHIdIHd/nY9KlJH7fsvhOKneZTTfa5m7cl9RtLNvwNpvGurnJ4U
t4ZDCm1A+q+gwhygSU3tFi/70kfIi5oBWyVfH32yYB90ePmAZSXvvydVCKDrH9ik
MdUPaxvGdZJD4GvY2AEQ9LoIldZL8/K6ldtz00pw7m+mAISYTg58KUWkCNkA+8ki
xx6XCjFra0L9oXwdf2yv0q/4r66FJFfUrLjJPp+bpWrytASi6IUbN1EJUpk7Iaul
yCjByaVIhrpoGkL4mGd+rlbvKrbku0vWAn/xjW66Xkrv2X6jTFOHutEScmUref5V
oKp9RV4/X6IOHk8BR7qzDFSpN+ogdJvjIk8dmQEv6FSEGJcriBkhEHRV6xYPQeIw
ZSjEU4H+S7QtPX9AeYzasyINMrhlgMVjYIGbQ1gWP6WvsN3dU/pCAITk/SILOHwl
+YberEdZ/MMqYzc4hc/iRKbKZLqHUM4NUov/q2ykrwE1mO7PThZy9cRzY3I76HRV
z0g7EauV7jME5EsMP8WTE0qHfe6otTqEVR1+/AyOTmhyryfBZISYCrTvZITfNzMS
sa3NxvbHVjF/AU9dXSOArFkuzuQtqNzV9J1+rwo05hKnCE8PoZpboAFaPsCoCv4u
0boA6LKGAckYLNKgemcn7/ILCKNnn2GLTXYYiDf/CCQznzeFJhdJPwEViMw+SBh0
0Lri+sFlfX+giJtOyb/ILNstp0T+A+klPDkiX3ff/7y1cfzZshRi9MvCc8pLuf+4
EcNUt6Kf6/WAWUMosHF+4FK5q05XRz8uuR+DtgLAh2FjEQWPm92zNuzfyxA4kMla
sMr59C5PeTOGqrTcKhiVddtsq0wuyRreS1g8+4Ut+z0IS780TJQpAYe29l90cnzo
fb/Fq62XyAE1c//2B4ar94/mjopGYEk17lB4M3oPuFkvZRMB61xwH1SFfjAY75P5
N8zrYTx/ucp+oLpLvrxAvgTPJ+nBXEv896u928R87bM9dyWiqwF9p8evyMK3eHcy
A2KK7+X07UMPOFRK3YBpUXEul67TveLHUqE6+J1591sECTbB2PiLCM8y8WqQR+PQ
fbAKxJeziNrSp8PwlIry7CulFGZGbBSCQ0XSmB48jqt3PMVAjL22/Zohk0HVLC1H
hv6jBzAb9F+Yo/Mc/x7aqXQIJUJGz1xYsxInpiayOpS7zm+Q+tHlhpwAWQphvRr9
lVGEv8/OTPHmPedJAzcLZ8HV9bRhut5ex8w0cjgzEmP69QLrOb4PL6Q/lEgPfrsw
XHrfKDw5biXsn4nyuwK0EdleACfSl+H/HK5YrFAK0aJXIUiK8ru4CJeHWVCKAJPY
l3sFATRyPNzAY9P+G9qbV7ZQkmMYQTIJu4UqzWLKnldOHIg7rB5kAuOdF23QxPa9
PFJ+zfurG/vZASgRHes9Rd5hS/02ORYx38vOg6Wo5NOla9rSziH94uSpblsoBqso
n7C7tDTxRhXzH+rVLXlhF4Mr6KxktnRErwrijP/7YrH3M+W7wY9OdhSspu8LaZ/Y
iJ2e90zjUxBQUSzCYFKNe1p275Rar4W+4Y9V1Lh9vwLLur233KtCHchZewwMke+C
js5+Y7yc4aSYDAKgypn1NIx8yVaEJCYR73cHHoaYSyEfhO5mEuBv9r8SQ2JgQGlI
u8KqjoiyuMnYbJ9bqU/pCFK4OrQ5QiWD9TwapOLWloqDg4KHNsS2v0Lm7JI7fjE3
EOZWuQLEBWAop1f96seKcFCiKCbkpYiwhyAAJrsj0wGRoF2VL/qLFVuFpqCr84q0
QCaiQHAwXCXH7QV3XKjWdTnYEq9fEW7uqFfA6FxJaDEHH9mrsZiKnwGNuHV8B8UH
nQrK/77B2BQQOyUFSqjr2T+Oqj3jBNWcCsS+vjY9/qI9eboj96IVctpTGWdhW/BS
ZX9W5x72z/9jpmPwThTPkXjThzfSSc2suPcKBFKa/qMH9/i4pMUC0OEJt/rOhExm
Kw7F5tKUb4Kab/2CEmzmmdMse/TxFKmOhxhG2fs/2uxEjOPjM0u2ZkhLBX1iEZT9
NoYjEbl+0NY3Sp2joFfUDWAIMm3RRXc3Oe2VjEszgqO0GxBq7oMq7wBPNm7ODJki
1TAV0xjZFSfyAHskr+zp6MS7afRCX3c/jDDPRw85rhYhghXndLunlp1jbqiSfsuX
FlOEIBT7fUNepMlCTC78tdiZ+LBQ8ViOP4Fev2cw2DpBrov08h2yx4Pn6vM/EL/6
QsEmZDZZFqlKphTJ+X/swa8paqxBMnO2BHLvOhPUcJDmJiczap8DPQyBdF2wumUe
s+pJpcvuXrAHG2okWyIsLf7WEQgw17eRXuQ+W6rrj4q25tUMUFueRk4CAHSl5OHZ
pLsp/DoQQKMuJHPySXmkiHsalrgW61g6jL3NFtJ4SONOL5D01W2L9k1QmF0Ge8+n
GNSgOUcOZSEgu8Qz/MpCx2qB4h3LZB49cQTJsucQ984KCROxP8lXizoW84V8wUE3
lf8c3fCjDhicgTp31EIydcRMo6xWO+94bqJcyVqBAbzfVI00IPQqHkfsC3J0+iUd
236h/4kO3qChTTQvv2rf45B/ub9ARFwuxJ6R9CazNh7P6pe9atGxhvC4YjNhZH0B
VtqtoYbOX3mojgQS4yVdv8o2TLKlhgWctANdZR3aGFVgTbl/W/bmdA8rutf+YRPY
btQN//ukCzBmStxmWObUGUSCLcB2CbbvTUyDHz+igxG9FTwbsx2DMTOMqUBdFB1T
4/g0hf5L/mDlAWx/h/XZXnTOybLCnf94JMXhxr8UdmoV4WXDf1GdXwA6nDKSZwEf
GT2XzSqf951etH/4MTZvxOk4w4oPC+ukfYxDxPMxYg1/61tkkYXkK/cWaLlwg80a
J9Jfz3QV1VSH7H85lndddlPg6PWZiX4HO8CFjOiZH+2v1SiLVRQZv1MGP5f9ig5N
3F86lbnEfvGk2HY2q9zx/8znqxW4q5RbLqsBvZGFv8IJcr5ojYpwOeApIrJLva5J
ECtC+4x5u3yjAXrueSrHb6IaQJ3wXg6zDEjG/XMB7igoj1XLyVZxWvPz1lY6a69t
vkxi5t2u0sxBX0p2X9UTKaEFvQWh+SGqPNM22cZ3k/cP3nIqxtOtuk2Zj/GLye/P
F4EG4xuUbqjER8xYCOiQxb284VKFmA4adb5aeQ5kk6oeof9ATjNIrRyJLI70fiGf
Q4BdPZestfo2NMmkGJNHx6J8KgIHgCcO2TCXXmauStaTN3/c17BNeKj5bz07MWvW
YQq4csTnsKuck+yB+ZOWPBVNMLvZ2P6gK9FFfPdnf4YNpxHwKUaWa6NRe7RssNN8
md4DEE/1CmVSyG5R4Bh8SYvr29qmvrKYWTHZu25QaB+buyTZikpUDZ3yWMTi9bRn
ThaQn3XeiY0gzD25Y8LBj1+uxrv8d5Ut5Qyo6BkdTGsv7VGuSOALdokPGo2XW8Cl
LmGp2kCY3ENRPWS1AqdHUI3O0Vcl5juDqMGywXHH+OIGZMHLO4/4MnPdNdPovWNF
NNIDltkwnVOePjSVmfUjeY79fFrFHpxXOGW4D85djIZiqzh03n4uJb2qMJN401B0
XCAH3Xnc3cWk6tY6xNa/1cKY5zBzs2gM1kso9uzvNt4I1R0jqJbXkiiSCEocBjfb
oDri53Q0i6p3pIXJlAWOOKEkIpso5SHg3XN1ZbCrd3fRYWOxkzPVvlvEx4BxcdA7
9YtcqLBHFrax0+D2+CwUwCvAHe9tv45YEan+vWqGqSN7GpHVA9rpWvGyzvjd2NLN
TkazgXX40/GuzU+lCZRdzhv+HF797mHadftoh7CnLTsMEMiLA+4F0/SAAj5xYuZK
DDSYdfzQ3SFouRTrtlimCgjVTHh8MA/9VtCg1a4XL28tAClMrdf++EtWbeZy/iYp
a2RAQv7VhgmqqJ4q2pJN+bfzi8ozST5cVZ3O2GarUQqWPR1QK9VfMeoKHFM7furv
tT6s1476AsUVN8l48oJKABTJwc+HD4j0LTlSBaffjTRNV9m/dHSAoPOJhkbA5RA7
UD1Z0gnhsVTZQvp2NfV/MBJdXfkd7euWI/1GGcCh90YMgJ8AR+/6s4jV+4krQfQU
+Ef1rVgUaEiBbY0HdbVaZaiaPmcoaOPxsmFG6ikETIQ34ld53azSLwVid25lURhO
YmavOvgA5z0IvhOUKiBriaG5zWP4cY8UzZGu5xYuHXRIGW23Gq3JG9HDgwRwWndE
KK4JAenKDmCZV5U4u5wn6E4XHhrbGoZQX9hEaWqvslhZE2vzSAn8cm1GcPNzdVqZ
A2eg5aHLiAd9QB48UBOjLhat7TXxRzfIbIDjoTOMwZMKId47NpAu9AI1Q7yGjLdg
EqIDvHhRjaMrOuA7ahE6MkhPknCtWAu6XbtkIuUPDPEnhsaXW+9j6Yzf952GwbIl
fbI3UknXDBj9deICwLROBJJss7qHzxYHO5CpajJ9rffeziYnbhJornptrlEPO1NK
aw4JTYcF9jIbrwW8HoKmNn+N17j9mxjW4OwxKsLhEq6gidYcZQm+VEzCyhGFmr0m
Xpm1uxfj+G/wDQWT/yPaKroxmOmW+d1C4WXzOMIxZ2Y97hIFo26IAVRF1WHqnJ60
qDdFdzlxRABi8yc893ZCIbtgQuOwZ31wTYfF3t7gRrILzDMTELce5RSmWD9HQa+m
DYYrBjqbWufElmEjXFULP3RYLOZgZJFtVPRPQEu1fKrPIpzFPr8gr6oUfs2LxXDk
djddVU8Z/vtOexvpobWf6dEHInRWz65giKW+svkqn7cCh2UzpGQdSBkcVLZC8uuN
y7w4oOQycGYrFCwybdmPqweaxilo5CI9kVtW4iOwAm1Cf6gLeffdUz4rPuCMkrSg
vIl9TNTSR/MrSpQKJtcypTrbcC9+Jg67aRvMSrn0dD+FpJ85fuXAjIXdPQaAXXpm
y1mKffsx/VUf5JZjv8gwrCyFFocI+n8d0PWRQkvot2RQMSRkqXn947QSqdmujE2G
9+RteYxD22oSn+jHEZ+B3M8TSNSNoKU4gJ42P+wWVdYPVFktCjaOy4Pb9ftMWnRE
QurRkt8b/Kv3kZXq7ODKssLcfcvBV2Og9ik57laYJtxZHX5wBmwb28CHr+20KtSZ
w9qI4n+l9hU5/W4mrjWHPtPidPamqb7S2I5JfOzPz7BvZUf+ih3gs3CFJvfZnV18
fo7IQcp9tyZ0/wM+ii4qo8vKE9YEJy2X8AfaawwsPJibConA4zRobgksZRy5PjTC
lP00/wLOi5/LCPpFQmhBorO3naaALL6WdzWzpDNFlDGDJxCX7hgIpYJhTeRtfR/e
Us4aKCLZonO2oct0/dhWzDQgKOli4oMwTGdKtVrU7rEs5OjWS0A1fy5YPAwewpmH
7zW1PCXQVxVu+OVixXjc5wGL2O791dW566umOn0G1oG9mb3jATncOH14VMRCt2dR
u2U65oVmtaJa+pi6hfqtlWtOWI9U1SdqZd+xyfQ+4V+nVxTuar8PplU2g6yIHpHG
+UoGLv7jhTBnM2ZDYcaYJnzVtvvaZT2erDhc/8rC0auflmbr2XvAcZfOA6ZfZySl
BmUb/anSy6HgbtS5kkTGsLDVH7OAdkfAcjQ2gqQpJuG1dYrIHlv/aew5pzGPTboo
mMheXMWPreH9jU2zCHs+AxXVvhovHnk/BaVEpDsCphNBUIe+WQGIeFjwxOmyDYvr
Dzy/2+O3aQsygMkzsiJk87aniWbShRS083BImRp1dG2YBcJTg1xEnKVQGjJUx0EL
prqHnyH3NwUR12G7hfqkQbYfAOqVF83feAIsibxs2UG2Jew8GqJV25mI7V3mFUEN
rnG5aeFf0tTRcOFmaVD78M+bTDxQZ5j9X1puAiNVHBl0XIAuW6/ibuuKLA6cpLiM
aLZFxBn/cjowoCi7AQqP9h5Wc1XbOcnvqA+5Uu20T2I/sfbIDs5H9rvCOD2NTKRC
s0ngP55QnDsyeKcybvYau/i2q0pt7xztdgUyB76oppkSknmcb1iYTo2TIalF3D5x
fe0dgSpeqMoWPFd/dEGGjZxX2ftcxVJU1Y1wAnAAnFT6x8LXkfloAEc+hhWNrMUS
SSMMlOduzYC/WY544TJPkNuhRUiDDe5jW1rQ8YwS5bhk1FG44gbvGDlPah7qJf+O
2qis5NTRmP98XbTBbMC9zwLXJW/jR/M8xqmNSvQ4OAOGZafqR8hzUBwVdzRhLhNJ
9HuIQT7jV73/BPlSlbIs0or7wF/nc7qGuYlLm65wIlpV54VrlXR7Bwm86sstr+Ky
H77T6nCKbXLJehmwdRZ7qECFpSHL2etWQj4PEOCnnG1vfBE6tok705GjF+xl6GCo
bjYiTZMCgvtAeiPqJSYV9rX3JSXOduboWMjR3ZDsrBJyM+pPYU6yx2AmJ9n/qJPc
DKPqRhG/vRp3hkSt344AXX0ogGMWJjWXBiVYNhoBYqW1gfNbBGW5o75tO48b5cv0
V0GIyJYVy07mIoQsc1VcNdjHTU5vOyVQDedJydS5QEaPk1clQTIq/flb26hyTo/F
xL5QKfZywLXKQM1ZPuT7Cv5z/wGUslYD9F64N1iStKezecv7CHIYl9c5uKIZWWoj
+lAHCnMH8xUsGfN/cGiVZ8KtiFmxcrtYkBv47+YpH4uo/YWF7dkkdhFScpMXWLRN
rHf/nCQrp+iR+vkKZcQNM0XAa6WcsBNvWXZAPzqfH3rkZutuoSEUN+2PGCf0GvIo
kHD0rJTU+Y16USelbTRIvxSBabSiqWuCbRdQDpx/m1CGpZhSeh2xOTRlRd6nveZl
HHdXdNL90hsih79Wd8kjmR1xMCce1lZtD3KvLTfTi9CaEOtZ7PgvTYp/jYXCL5jN
HalHluQfrzUCD5ruXqfYW2tfvBEI5dGtYK64QYYNCbj402ehDr/cgO1vc22F9SIS
hFIXR7h5Uw4404ODnTkleFKESAKPqxdR15PEqu53nKccljxFTLuMlVTUlKyHds0T
qnpZ0Xzmt3Bq+g7Msq91ugNaEFHsLLLbY1JLh8fDDFQLCZbjG2Q2DUUb3qIGTKu4
gy19ManfVpHE4T9QA8ZIcc2oxu0gerUfkyBuZCjU7ICmpQ5e6ivgY3DP+x0CoiMF
7pclTp4/sPWMi8Jx3jWfrmQQPIbcZAWu4C3EY9i7pZ+q9ghZEK+JwlAH9wwIbO4z
E+2by+yMtFJfCw9si3P1qpRjeq97yyG6W+IpNgtEUadz9ITbWSZZo62ephK1lKFy
0v7jJgSTp7CUr5oxPt6SA5KdB8MCVJ1GO0UR71aklC32BNhwAdNPkTMLjHTj2jpf
lT8Wz1XTaswXnRiF4QE+r8VW7fHC2cP1nHwxbyybZ75mM//ayhu8qzCXnaDMJa+d
1LaitooYZE2EzstAIpIkbLPAU3o2wMTDVv3b8Pp2jtdtXcquuQsYfjgPiM9ipzzR
a3lpH5k9wG8SBEJCJQzJnWjKzrBe+w9r4/5+QdXR39EJWV7fhQonjhJi42IdLNLv
Ua5eKZjTrYL4QT9pgeG+6asBEr2iDvMZNNSzULTydXOp6FEeFZ7UgJsWZMfQQOgl
sxU2GXO0YGHukm3meUOG18LPzg+31805aKIbU/ysguFR5zLnMb7Ns79CrCUib9/t
ykKjlcWxrSvo7erbr7grBQlEFCBHyypxdCCLOKwpguW/IKPnd4xBlJqD0jnWz8OS
qyyC5McvMGYSofS1ay26DfWTNF2rqVGwOjsWCDLNC7WufZf1jZ3D7B22bZ4Czi9I
Bo5iXBpFh0f3kpmx+7xUuyIHpeB6XsTRc1+7PxH48vlPhUg3zDTwwGhuF0PpEjXz
/FdkLQPq49wRgSKH70EPJKmJMq/KKUMzMtFWpdEV66h+jC7jVWiqvSk5CUStdMey
XESYXNcx+GGIREqAAp2rED8s3fAnodoM+a4oEgIZ1aLjXg6hZsimAhQiVF2TRUxm
UEIJOM1woknBSJiM3YEqAIZsxhLJEWUvi1D42vQydLgqqBDBwESGFvl+8LOfvi1R
lmoOSPrat5yBIrpFUAHG4w2Qxm63jPNVR9urdPT75oTJdUfnx3jCWbWElrcvmUnR
8d2OEFfQOZtBoFqksm1ytCD6pG751HEytMmIYWzLA0An1LvfYlrOuu62cXTGUWa4
zwChhiwQShcBI4bU8KlczSi8LuRWlq/ILnrpYQVtzT7RO2QD9iz3t8K0UJIN+zNs
XU1+HaNjd3YQD6H5XjviBx1i1cw3MJKdTvBHSGwvQRy5EKCplqJpt4EQKO+dI2Rf
wlWI8ONvFFxdxpLfYCeEMXiL5JY/bWDx0sVbLZ8N6Wt/imULgkSI0JcDFRDRoQuH
CffCN9C5b9CfdP8TlfubuAjls2cPK+BRdXLZDff14VbKM/asBgs8HGnuQQGmzVvM
5i/pCK77CSCAFN4Sjt24xLisJBHznD8VmHX3YoI0boXEw0nqMKGsq06bDzHvCvQ5
Q+NlRnpSNHDdf4LVucvyHyitG0MY2w573SrI4yAMAMQEbqdIV/J/14B8NKarjWC1
8sMS1mwkE0waUJzYJdKmHI66k672cIIM27z2V1zaUBJkuR86Eje6JcLP7xrNx3ts
m8D83mKmX6C2LI2QMi2tXJX9RMXuxRVw32m/aHg+x0BuVDzMCRUWdPxZJVLxzxy/
gf7cytManMFjpUfZp+KnZKvDFv31/2Sf1o4O8QEBXiNKQ2UUd5eoa9uuo7fUmWOa
pju+wbMK6RwJ/yQll+Y6DdDvy/JlbQrWr1ZjP/Wwme+sn63RVugkUayosZDQQrxW
W3lZk8kEpoPwa62Q/330jcT4kAxMAABo/G83Rdigt+897k/SSrXPQemhxIbjHDjn
aNZ2pzwrS6wLAIMa5+VpSGLTA3b7YS7TLXN/U1B3WoHQfalALr1sbrlj4SPNKWBF
Crd4rJNdmv+ZRFZMBzZZPLdSlQ/9kku1sJW2SFRRd1DDE6MLnuTmMbeHXfJaqZN5
xdjt0Lk81djzB/DX5iCJpcOf/FCTifBMgeV60Y+CYFtUrFZn6nPeMcHOPaNB6fig
Qrf/s1W8O+ce84DsgzGyKub5f+4DwkXuRDQ4rULMJgLk1sgT5yz0kmrWU9ZJ+Au2
242OF0HhxoObdFBQ2SAwdvpAGUzxa6kPTMhCwhtJ9Rt+2vFXV7NrZCnfkYEKlLnr
0WxS4a4909OVvBxEsXw1lAGSgNS9/NJ2kP4PJ0RTqyMId1QgQbTeJsmW98yHIxri
jwXewRavrMQhGON4U05TTSLIwudj01Whhbw+gHIqaPBDpwEFuIYz9HhEtSnVKoZr
y58N5CG5WaMBgPGBUAM2Io3J9/Flvj/KQKmP5WwIpYYry4LYVHXP9vgoZVGhAbDa
1TdOw0qYqlQG8fws1i1XGm94VgvLIlekBI3Qg68bt5FiNd9E4aFiwoNRppLGb/EW
4S0kHJJG9DSQ06oeeXJYARkZ8Nb9PGI9VGL439LMYlYGQqxUlnZN7tvoYbq06zgr
7zQlBbf/3R8CsCqEmuROL6x7Wcji1AT9r7mjT0bQy/GXFQ/6nL5usqnbBeAQxi7r
/Z2HoMWHh/HkKREzL4AE9h5Y1hQsfo2pLv5nv/R3NPXe7pr1C9YfAuUaAgF7w3Zh
WseW8gxcOkeOn7Gz1WvfKIQX8DRI65IVWuWXEKaMSpmWuzgOA0zU8ARAOg+2u80H
BZ/tG8y6OpqNarB+mG/4Xun7ufaEEKIs7HYK9X66AslEbeojcIaHu5mkoLOp09HR
1SLljTorBOiMm0ZeX4wJob4ZeLtxrE63ZI/Umxuqb20zErRpKgO2FX/lZOMYt5pe
hdE1HMnzTYkIx6ce4Nel5jC9WTmfu+5vngrV4YFgOFl+T56EI2Ck59tuaX8A3WNo
Ga3d77TKk/Ytnpr1dOu/vQmXOycKJpl663YX4jluntWyV6S1bfwNnCQpbUNKRT8y
q9PfNbG5ArHFOg1o1VP8g1IJ8MbO0zjJTQvMSuHTUz1A1toaSk9BeyXMXXL76zSI
H8NDbYeH4JqsMDyqZ5pnEG0qxdsIE0Mevo2C1ZPelyrjZN58rqGS1Y3KiHbcZP9y
D5TSTfI8OaLWk/h7+Nb88KdeQVfVYH/K98nWY821/Xomt3KZTKifR8g5Y+hOMO+6
oppOy/gS4IPM8dvq2z8g9ewcY3K5aNEnN/5fhh6NDy982BsPNjp95aZ0FPd3WlJz
leOjRvssytpleh8Z9bCrnbxaG4Yx6KSqTuPdMD4dYLUWF34RNF3vrmKGAe3FQlwO
Xuc26ySSWBY74m9sMxO262Pos8VJrQ8lxBh80LL+L2tZwNuCXkyZlSPWD6eqky0R
Pwq/a7nqYLBmtvrrdzC8G0tl7DUdYzub4bndUHbMq7nbmWUqJKqyudMpJOGYPVUs
qT02O3IIqXOGXDfHo3lQGCMG6cVGSRbvjuY9Z23A/4pRYPYK97UYTX7ZWIao2tfL
B0jgxBamrBj2AIzESU+0621uE18RdJb51I+J1kTK0H0p8lg2MIpL9oPOsOYQMtXa
wEeQS/siTkVPH1YuqmfoFewTgc1WXgC864j00mpb7MlRhS7jivGTANSsK+Q7APrK
IphBbftxUdKEm2vRU+asH2Dy1WJnxm+SQg9O0MJIlub+SR/F8mW25hjD2+i6e4J9
QvujfhkxzipIcJg68qM2OyQNjETIeyE+oRFISquloja06g6laErFbbuugtqlaral
kmb0BHtWZJNHQ2GesSZ1a25K0ZxhyI5FzSQtX5tWmAHoBTAjZ4De7kz19QnRtfY8
NJ1v1BhJqN/cdWA/8yxCpZf+DAmJ9NmCC5L2tklZmtflHUmqBNpMoBgtMhpkcsyA
uy0ub+WoDwxWewni4+V7aXAyLN1pWW8tSgUFMomCZYMyi48ejAXFckYGZlrApqKC
++NG9tBC64eD6sTEjZyFNqDmQ67mONhJZWba6jAsTVdana5RZsXMD7s0mw/TiU4m
5+rzabQG7iBxKH1sm5agBe67e0YepAgeg94xlpJYppXpRBLttesaVrj9OnWsU6Yy
qVZXQ7do/qFJeXPD+5DRRzEjhSl1WLW6exacT+BbZD895nOhPIzDZCF6yy51sIoe
SpTJihi64bxdSBiFWh5Dt7ihqzBgbNkoZcxQnK1BuG6b0oBo4RLukidjp8bwfh5J
RSXqUQ9ND8KbOHRfp1lGWOj7GfE6o6JYRm1ShUXoRL0PQyaI1iG3ASzC20eb5hgr
WexPoOSJK4UIMx9DOSl8nNdtVudgVSooH20zCiuJ5WzQKOgKA/NMpu25MYzMtm1C
PdW/7fUUJpb0AxBLdxf+eNMi0iZJzspm+WaeEjJF2lUo26MLVRxMwMhW2NZIs3Me
lubXCYoRfVjlJDsk/waiGpy5xrz6EwoYNXDzdUL76q72JOMkTDJx87SxvNd+hcOb
3p7igudi6Fhrr5MDq+zlxIoISIzWPNwPT71riEiHz2E3EFI9VO2YqM1gW7Fk7wer
K5Ake//ijYWaIIDKM82G4n0ii+Np5gjDaJ0CTiXwZFO6TM+PxlGI4dgV/Pxzd30Q
gRx9rOv5R2DmX98JYS6KcMTTVpgWGX2qK7hE5V2uWRjJNSzk6VBeb3ASxCQwhFyt
RUMD3KnMtltJoYlLcLlM6ACaGKjhs74IlmRlrp40PqAzCJn1LpCfSaaUCqBHUz4r
PaWNwdx7bbpgTB3zYwdKm2rrWlXVVH2yXAQ5idfPz1kSscT5GCVTTAz2+zDXJ6GU
0p0d+ZBzrW6H0/yQq8kyWGRIVnQPEouNjb6cE9+fNgymtBE2pxTMOBGrOdtP6q5L
kWCJiXWrs5owHcHdPrBy5k1XGKw1UCf33XuzL/Sx4LT8m9jk/6T5zJH0xvJQmLDZ
7T/Q14OnO7Nt5SB+2/nZzGA8iMJoOqQoRfKb+68zI/FLgjstNmLlRlprrkp2EwWL
vQCODHzgbOmQGMAtvhO9k/eVrcHxBETOnKwtU9upPzBDq22XmdYhkes2Y2HJldiK
fCtlIRYzBZvnhUJy/SfXDBXk0Gm8a09u/E+BJYAX9uzELZZiAysz7ugL/HOPtPpm
Bi8XUaXYb+3op25WJ0i3ir/Y3kISadu3/ht6n2chiHiQKBvkZfdgQ4+0H5ouxhVb
ymfUBqs4ssUisRlsvXJarBWkgHuCBvMDoPasnlcIXXkgYt0OLYMeJCneUuOmemPY
3buKBNLvZnxqqLmGUfHdGDvmc2yN9tZQVk6egHP7qjie6UHF+2KfhvJ1fvvGhJ9K
XjHEfWWqMrULf2Ap2CmVk/bskFU+iUhbVg31wYBU3d0YTx00WFnnPcd1CWCS/3m3
pSmLEtKDm9qEYmF+NGoBG+rvruPWXat+7zXr/T8tztEkgcfGfeuj1W1yA4E9Uz2H
IaaMS4W//lA2qqcbjf7CaQTOxb6HQ9F6cyDR2qYmIaFf8uXC1wICuwTu5xvPfxAQ
+qU8ycPWnlGaTV+DW2kkIoQnCSg/ve+EJ5JKA7AnzfipRQoKBAnN4/7sxTYcS9E+
h+ODxtZ5ufbpYRaYmRRycetLBMJVSNGzxO5vVRNltr5N3Id6QiFixAbRNKqLCKLY
BOsqsI+wkxh5JDeWLBitqcn81+9lYAA8EoOyEFSieC95KsUf1Vmk4XSwDjKX+EZx
Losz43aWa9gBCdnBvxhvsLPAPxc0jQGnfEdzgFs0FC+Z35tOCjxZ8QBWtICAF3PN
2LjZg3icKLEgxqGAFxE79CJGSR7kHW/8J+OSTnjh1w3vsAyiAFZc3p/y4UUVwW99
7iq8hBJoKmymsNnOTxdMVIb43I7tsGdbm8s7a6ZwMJlP1oPw39aGnH/iqPeZjZ0r
i9DRx5zJWGqNmDnEVdPKcQRMPlvoemH7n8ldhFLEzIyhkQgbXZi2lT38iWSECSkB
jU7TyeLznHKbOU2tBlMNu6sRc0ISIGFlcSWC5br8ReTb88BLV7hyEHTjBbBOZ8Rm
pJ7qjizxcdcS1flLYmJ4ax/jY2yHkKkw1ls9k4hgbIR3Tv4ga3hPEiFpmVYyH9oB
m7bra4oMp9Wcq2t3pPLCUSKeRDINIHIlVH8/kFhUecNHK155Onva+/FnE7djgwWa
bFocy/wT7h9t6B76Si+ILTsU160OYNddajrMTurS96UK2jMmsuLFgGGjSj2Lc45g
jMk7mDp/JFpko0IQJU3l6NqAM4Rvh82aQVNBXVEIoWTJiz6te2mMBjST/VLB85gF
D3bxf9JRZtdiXEGA8Pa/kZCw8qZc8G5UJ34e8UPRDc/Y+4OSezbwwEoejgXlXlaN
LkGLv9kMAwem1GoAB5OLsebl/+Iv1a6BZsAejp15NfuFdBeQyEt4YMwZd44R3CXg
IpWZ6Yjc++2ULBOcnbR7j0T1kHFD9jwfO1D7MLQj7w9w8JDcz7NvXJvCHwkoo3lp
NXZa2ssRL77zD6lLPk8L0c0LPSaNL7dsUtpTk6Mw6LDe2EFXZb99ppFUkEGQ08r8
pcIPgLHDzDgmIKkRnE0UjcK5AomDOHmaoAvmCBvwwr2GSoZNXjMYXT/3sufG8/pD
jecnGli7aFK+dKEyc2l90pdKyzeBpx7sGmEQEkWMxMUVKsSxLOaAHYeVaFI6Byaf
Q+9gJIN09F3D4gFRKWqa5hUMLFv2fmMQUdthP5NOU/DqGJKgwdNPN7wIsIKzkUe7
jZkh2ZezGxRWACUIIhi8fKIK5mhJlfA8H1Ov0LjGP0WnsqepJUWc5b7sLnPDdvxs
3qFjYyQrBZU1Gjz+8AM54gWWBXHrt9qEB8jwaAK7VTe1t8KHlNacib2dyKRaYfWs
/ivbH6rIn0Cr4Una3Rz36SYzJnLNXxPXJq7coFt+rm4YcswJNHNIceCjcx3tZZfZ
0FR/BwXFbb0gITT/LI5qULJaU4azHTcOpC2tV8TSoALGaczxzV3/BbN17w2OlBnC
sD7TvvRQxsQAqRLcEr+GguB2EWnCpmGK5vmFi9vLD3zTFukpAvIk6jdupxmVDM+q
Y+4EYYzAeyqPLcvEkzoyPH+kTo8zT9WQI3c7fIVUQwL/9FJk29+HzNYD2WGUwlAE
aT1lQBJ9kuZAEt4U6AoBoLtQNTvJ6wLw7yoDgUlmdc082ZDdvWD2kCpfIzh6mKm9
EHkJk/LkFC/1Gv6R1d9LMliCy/n6PLAl4XJeC7aHJ1TO8tyzdb+87AjT9xw9LtGX
iQ5PEMiVkKOWwprStgdY7gduBClEESDy7HAwtghe2ihzaxoL0ucatHz+mVDXIt+A
qFRBb2Hx3aYI09I4YnU7e/wkwoQUYiiBcj2GpZOyGaf71ZB/qen9Q34ctf8uj4+w
uo7pqb+9KMgutY9CAk3NktPgXHhrjQsoNQAMxzCfq0sUVJfBrBDVa2vFoLF4IBVl
9ZbGkFpGcU4oMYFRqwcA5iQdMBsNr8Mzg0+kYo/QKmeogZqH2J1nYHvVs+pQKwLy
XYG/BWuzGwbE14uuXR/INeAwnMs6YWTLfrg4lwRCjYgqEEt6A3M5Bew2Kd6AAutr
ePfqtnCtThDtciIrN3zIyU05JjLF1R8tGj/IskxpgMbhTkvo6Clf5uy63oOkCtJy
wprf6Dt/4+fr3i47Mu3ZgP47M1xwAdoU4dZzX3/4KU4XRx0wny6e5wTfjmGIxV9A
7Kb0O3+Qa7sh3q74NniqdSTURCDzLLptwJKA361e2k73dBCk3VA41ZBgiYP/PaPx
5Ro5js/X/TICUd4z0aK5L08mV56Q7vsGzd6Zjgr+OEhA6CMkV5mMGoZCWC8zAWSP
zDjxdpHgxACAeg7t5vKOmFDLR+7j4tAQ+2HFw9umkwF51UFshFdhtsHDtNmLSpki
FnyBXF6bfuetXCTDuCTJPbpJOmPSbPbWD/jTR/Et+ExI7lP31zOGpD/SbLJn57qT
Dp02LUOGVLwl6vqsAj958pEmrDR38DwPET4Yj4P6An+XeWPwCm7jZ2HnTOKcgIcj
ZXXMbYcgWpMdbY4ZIRp9BCfHzr1ErEGm/KLdCZ7wuBOFR8yWh7NEjM4Ln84ui1ID
LaFqbzxn+gHFknsIrOUH4Iozs0wZdG0ZN/bEbBJQeses9SvE3d5HKFx8ZVuaDs9n
V7lOszHmVsgUXb1+p2cYfG7NY1zxUoMHqJFnIp0/38RSViKPUmTyhcAzfWDhcUnL
mLlIjwTAU/OswcDcilCP760sLM3ThZSrmOUAhm6Zbtq825UJLKNKWGI+gTRcqy6f
zZtxcDuCISnPKR+Fc3sMG1NMW9PlTZ+uqF5L4Svz18arTzemCDFg93/DAURly9Iv
zJu5SZ8mL1HlI43l5V123D/NRbVHTxBKa3uNh6iIp3OBeX8qk22wfsaBg1Fjy1U4
j7pgMqxcGPTj5YSfBevkE3aMj06YS+5pEJNeDG3Z+jBVamfIPWWo865hmYAH6R4Q
gOWfxqAAG+2Z2GQzjXXVc8AlDI8cDGNDQpFTtCt+VaAqgBsI9/TBaUtUXNtpvFQM
5fqUH0iqh4ADIShsgE388CCGOUSAm6NtSTauefV0CiyeDvTKXoh8UH9xVIg3yEhN
cWU4CptqsyhdF1fkIZsk20B1qsLH7MNXWe6FNiAkegiihJQVMlXLscM6ubnoloez
PAYyN9qmN5e9U8j7QuyZUVW62rYEpRni/D1gg1SG99ezJXZdmjA7z985RpnuFW6/
r0jao8cz/LqPToqaDhVl1HO3Hef3lRPAuH31/EM+BxARvC0BXfkZg+QzEVAMIubz
Otps+ftJgFHcAmm3ZYMjEzxOaoEZFqbzmCAHfx97gPt8RNmyhoztwzRCA27uSdwq
DP14B+zx9EQYLLfTQGH71R4iZ0wxPCrBdlL9WRanmbXR5EkjHxdfWkpTsPVe8YMY
jB6Qh1dPootPVskO8TY0oGhLTYdA1dBx4bmkPlfo07ODaj9p73mnikcWRbriqiQX
2/YSqX9U+DvXLgLzrNHddUpaUgZc5A3uR6Jbjc/F0G+sl/15TNzIxdX8MwMlC0u5
gTOPOTu+xbOZcNJrTO6kotDXq3LkBGlC2k2ETOsWMEd1qEuX7IlrKWZG/SEVo3IJ
hZaOvkm+ArZxihIWwNvFIJqOGegojVO05dUQzLG0+cEojSrV+GafheLsZYQdXXFu
uB7pIqHRyLm85dpC775ZLsXRF9kARWmaaYZETCxcLBvv0m+x5AQs79wQtE54kc01
Th+6Ct4cKs5tkOjyPmKrr+3vm8RS/uNBqtCB/f0vX2NTJFs4zerimddw+2qMOXOV
K8fYO/+Yi8BLk2S6jcwROEXd0ON6FrgDL9KA07NeplySeQZ8ygC05LxZCpDVUdOk
GkqoeHGnCsXJDw+C0XhGZOESPDePE1P8QAXEesQOVUWuDP4kTlyLMwQacpjjAw9U
8Qk8w/dqWABFiud+trivMFr5kksDMSQ6VpHOZ61s0zI4NdyFgSqOcJTXaEggVLb5
WHD8oNeI1KUjQz99A5iKshGkfIupyUoVMz8iRkMcRpGMgPJrxq2BwhOtoSqwEjVp
EWg4ZTT3F8+ElQVFDsT27A3G9JiNIu9LBOmx3CXWodi+cEPQ09J4H/x9bArcdqT/
eV9/ler46v9wuxC92zUyGNMN7C8jFNYHnuOVu+q508pqQ7ULIF+vu4bJAHCXcuTv
Z5ZOcOZk7RqiQ8aD8Yo59dCaodlbfQj/S+6M7nlpJu+pJUANBC5bkdYD3eYHvi+K
Dz67oNTq6n/a1lSLgCMqYNq9MPpin4pjdFqUafXMswxIP3dtcELrTxdmKAMOePKT
/REDRt0UD9Vl5m7qtMtIHFbu2M9PgubYaiMPUnlH7NxZMOjVqkgAfzOqkMS479MJ
XW7CGXNC9cOeYWhFzqXSYNzuzWxZmyOZG1HeAlL+GRcIpKgXAeQkTohA54rihzrR
MJ2cAwr4w3koUTjl3Dg+Ty6uxmREXcseaiF4YAkFXLdA7I4r7PcyZErDpQr/zF6W
fw8K8tAl/87C+H0OpnggSjaJLwlg35ioIqI9gJG3c5eQiDuj1gwlWoUz/g4ALP+C
XPWsMF9Q6x6qvxTJLIkhBoaI+/A6+aUlJrQF849yl4CuRvtJGo3BvDua+G5GWyYm
OEklWCnZIwTZXk8xUw1e01xzc3f1UNDCWJqZ/IHw5Hhxsik22idlPVjWZkPrIEsC
K8nrx+FO6dnl978cxCmutTp6oLxUgWWApfsSc2jrwbQg507HFLA7uv1nRajPWVpd
Mujj7Zp8qZlCtQsSc20yZDiTm+KnZ3vPvA7IAqpgwciTFbsSlarKoDEVbKqANwG7
VPYLFVOFDUR/Rnr6pyvrYGKNgQBp4LGHwYM73kx5yx5JD8XDU1hZZTXnTV/EWRSo
b/7w4+k+sqqI52rwFWYySpf6QvO9C2mXQTFXr4XZLm9rltStM7VyNbQornr1btEy
O+n3uyyNYIVwTE6i+yAxWw8PdCIrEm5x+4qD5mKs+0b6tjaFgiXIScfMRJBp7J8G
vZNBN0bG3SKYbjf+/zq29K4H+yWvClnZukgdwkJqnCCT8QXl1iCg8obLk0D/ctPx
HSC+0G0M+2Q0XPKPeDfZm4NjVOReB3JPkdwuEBCnghG+GRWSTzFLSSx7Ey1mc6eQ
/dfeXjPEHz9GazQiD5bSR3zPrpf+CRJW5hRcRNvbVn9bU5D9DNHllGrsFcGSc5Vp
BSIL/QdLKUolY/9jQqvzWF3c7hlKQUg+NuK0so6iJcQoHqq8ZdEHYafYY4vCztaT
uohtn3s6wrnGb7sHxDLXj1CcYpFNIiupO5jEadI7I8ubQ36OanIAS7mOG4d6LhwH
ZHrnyt9qKaXqhdeEts6GGB8j1p8GcGHpFao/tbdQJvJinm2mQHdtKOjWe9Pc78dG
P0uEQk5Pk+9oO6wggDZlmq+gCvPk8IzEAd/utvOK3BVNSMohYn9NmLC6rPTOxHfR
11O+Id9APTUzAPe+ZHKAHAQcnzcSH3SFSJ4LY7t2FjtxOfmc9ByLlgcyIH9OWM2d
lMtfFrAkMpYnf3jeulfUR2RDgYSst6rhtb0pba9tOL52z5FUBZoGb1MMwb5qiUof
24P2JBJlM7/B/cyVCvLl0LMguvZgSeTg9bx+H/ppeUHWHXixehqUIs9a24o+SgJy
hHpaiqI88lCVetTWtv63A+Zctx03BCVzP43+Rhxlh2jqyg+VuxPXIZFFSnZ7Zbkc
xuK81JX4eTfAzCnwEA4oph/0w84hb3/gdpxJrQ1Z08HPxuBIm6BGapnhQITiKMCZ
lWIaMCXF6TKDj+bSsX0z9/b+0qqM32ERfaZV6XVtifBz/JVAKDg4P5sYQNxJ/wYs
JfD3GaEOXHK7ioypcX3cYNAqDtPCd2c+kC44o2+XA29OdiYH8zEV/X0guobftFUw
Shjm+X6EfxYT9RpSFDeiFslqP3uskBNjzYKdU6rJCBpbaStrmacYgMalk/IP89S6
aBk5BG2eSekpJ9O6sTB2ccBPKfG/1MKCyG2/9IloliplddggAe9sDsGtMCavKAXF
RAuSGpRQd+qMtBqeHfdlViUVLnl3fKxPIi1Gwj4Cirsu2P2+25oIXymgLuEz4/Jo
FY3GJ0yAL1gshiU9jZleSrrAKJByayZGmIzlPA7eYqz2shLsvLIoSusDjM4P7NF4
edcIFcaDIBwgp9efkLMhUlGNlcOt/0fCj+RE8wXmo9Q2RZcRRPLSJ4ZAjt8VwamD
549yAzMbTMeFdXEI5GcP6f3/gXtPzzYCzHXCbFM9ebr/TXE0ZzQ1JYrH7PcnKXz9
4SHsMnzrxTbphTbZSIj0pbffgRz+RDcaooyBE+yVyFri7ulrluYTPW/fOJ8mjYNF
zVVbwC7V+ZplTKQ1eo/rf/luRwEsseceMP6gkoRkXQRAcZ94oHwJIzY7MCuGvkx1
kvxX11T+2zZYIlx3ET6k+OcTy4iKkPjQbyyRr/cRTGVllzC4TjzG4ZkLWi4KuYH5
8+KuvBFI4o1cfFV/ye3cj49e/xkUJsUfnB509l3EcEesBP3S5+G9kQuWzzW9bvKO
GUn8RJwsiNzSbnPhvPqathPIPXnzoOFkYRTKeJwZztHocdZDT+BirSxTR2NAgelN
JftBjc51MFw2EVvmlyhz0pLQbSRUJPFRUXv99lnm7IdgYbOQoz+RReYwsm29YqfS
uHjBXoQNw+dmqBJPFuM20sYur6i7K9jykHP/ilkdHMEMSEjOjOHvA0O8Auf1azbg
t+GDnBGwl9Btl+/djHD72u05Bl1cOvfm28J6ArRse7ERwzZgZaf2EBA7dK0gXxbc
Oz2oQj+ZJPbJILT/6sqES9dQR3o+W1tpObaYUAu7StkvM8jjSJCPOFTyETowFkuy
U/I1ptWYJdZDhCAphDML4JvWnTTGwUvziDIGd/3GpYC46oTE7J5ZxK4Nq8T1mNrP
9OIYt6dMWqrYhv5KqWFgHwR6zfoOCsni44+C0RSPpFvGI6AS9rqrWTinoWYwuDn4
uz08npjMmOJe/+90n2PPrOEdPuMngnQCb0OG/89lsXG2CzZMzjvbLl+jWJKdrewO
mx574o8ZbaMCvqJwelmdeZ6fp3pOwCCl1Ol6DYGL8J8hpYHN9PhrPvshUlJ4nM6x
QSe8cQdM0O91s7jDlRp+qaworR6Dv2zDMoooOEKr+uyRM1oqIm59eGsI4dD8Diil
Wub2TP8G26zvZmioTS79yytjccO8AylfYGfWZjGollMXhwc2z8V1//EcFYwMj2vE
kqprtvRhsbSdA/9WjOvBEs6I3UnMPBc82JyiTz+gY+5tUvOgWB4QvxtE57OYopA7
ryMZb7buDtOfdvcU65jEOAkfJXPngWySpCoOQcBdKvz88/32tg5LvkbN90dwPoBd
itDu6bc7GQ5uKUJTpL7JE9PsCcckSeV3Bxr1JtHkyFjczc4MZfZC1vX60LyRp8mP
oZBXr/hgMOqdiF4B2DLXufHV4ddnwGVOnxbV+U+Wp6dMeF+BLdHCtCQ3hLIgqPPr
4/exFqh+ibap5VcLNnD+YpYP3Woxamk3I7WhSe4RGoU9T1bchvya22krUgSN+1k2
miXshYqxW+usIxhLoikomnuP5bX5cHhoJbFlAqetBDfKcKyQlLo93Kx36P/CpSug
z+WfV3H04iFyCK4N5VpD4yX2n4z4uev+on92tD6kB8XZ8PbR6Xk2BDqPRLERVMwP
z9EleHBm0xaCVS/+VpDbKRHLm5B2Pnj+68LHAWq9927ZF53rO54gsA4KsreIJKLy
UT5JUOJAvmzRWBjX8MNKmEfUbxMj8nuU8Up9cEoYHkX+j7Vh3djGgAjEiWKs3VMa
WHjJByVXNGKJyw1IXD9IkrZPqCk1PHe31a8ZqSzshSmIzQZFwBJX5le1+BAnZH5L
pfYvfeseTHlGl95k/3xa73QJtkq/NDU33zfe88VpJwwlqb/t/q6EFN0r4rVPF0IZ
kFnQ+3X9Fwv3FK4ZKWcKWHBUn4aa09nSb2IJ+G4KXWs5JmbOm/ibxE+8uL4I7Kwl
hmBK1iL7/2VunQFqkYv971McHhDOae/JAKuCceXMtuKgyVGtr8m6re+sTZSKlNCX
076I4c7JfYy721DoYt9h+yb+ABep+Ma+PhKQVWHdBQiZsobMVKkvrAgbHIB8cNoW
1x+7+jg0a9khB2xD7hdP/VvFr7+BHxT2Hg2xsR3+pGZ5ogtX+uXrvXrD8rp03I4v
DFtt34StLnM/xb/LJF/gxeGfJ4WITSnqEInPaLyL10pBjiDiXgnGSYt35A73w1zb
pRP/pXwygH0EeSli+O45PIbip11ZKBjBTVaEQ0FBmnSP+LfVZOxmbR3W1kUpl3Db
+lF7IyC4lNvHweL/nZ9cecvTzjI5U/gcLaDgnkJ3cTiqYM3XG3z91ykOS5dczYFD
rJEur6f/LbVUOKwpjGNFMqVIjiBq8TpdLZC4PM54f3KvClTkggA+Pnqeam/CWxGy
+6bMIsEhhmkIxD61xD3fVYV+LQ+nfXJ6FPPPnJRncyaZA2aPQ8KWJuRQNX77u5Fd
eo1JMaVas+xZoXFxl04YoTwxn2d2JdeBqW1RrpdaDvn2MWEMGinZFgenKyYnpx+l
2NAMr9ASeoi8kV6m4QVDD0c2yWwPFx74AtfCa5Tv+U599XL2WJdGzPkWr2McbV9N
fJAKnJsuyEyRlpjWKTpfi1rcpWBRm4TjaL4gwgav15LiItSgr0AyjzN9U2ZRRGg1
kpSjDuoR5HWyQBFja95VcIscYprMpUcS85EF/BBP0zVD2CxMgsax5ZjL3qv79ZK9
UQa4+OUk34ctEkPlVogsva+cqFub2IamyX/n/u2cOs8bboY8oSXX6S+bR1wkO3N6
cR5zWMLZ6CCCyl3DOhBfGjUj7ItM2gClORvRlu5k7n1YNulnFW/eJ/WvBat6VIUP
EhyF8mhKPRi9cz91+nvI4Il/6eEd81wmnlS59j0mePU4a0MuGAdca6bPTtvfhcpF
cIiQtCeli4bOzfUCa5zMGd1mB/5oe6Kbn+znicoMei5Hz7dhFuRiVMZOuLbF5lv/
RV/ex1Lb81Y54nUcY7In2QGfjz2k1MNSdV7ZFnKDffo13MjaIdXwotJdEW+Gj9zv
Kpr0JtiGajDwfoncALAMxNz6nGlga+8y6Ftj7M4BhUgFcuffIofKwxePzxPG6grz
qtNRKOaqpjjbK9ATmRE90etIxzBUqjart9eTOV1OKjGmjuAuWSw0lWa1C+W/EtK3
5CfudHkb3bNcWdaA56FAAwZpJBemDFuV7l5for7qlUndnRdKk/Aw4IjaESKclL67
JEy9g2PYsFBhFGx4WKmSTDx9ajMzKe1/DPuIEtzia4CghGwldUGxsjt6Y1eOfDXi
5/Iscw4e8OQmH+S7KgGh+vqzr/OVriUuHeJ6C4Af0MrUia2AT3dr3tg7K+K7ZTZQ
E0n2El1wKIlJNlhJ6U1k2Lxoz4tI8uFPlRJGIo3+1xsUDiGglt3XkpjVD1C2AwPe
g7sHXU0nMpjJoKTepSWwYm0s/r3Pzq0VZ6Hjr7znmYHO3UtrfeZIw8AG+3LD4S/f
p/WmKv73JZ9swrUK4UykBrYix1RnXNhjCg2eFolvsEjqakUaRxSGjigJYKMDYQVN
ng64S21WGl3yV51EYQJ9ggF31kW4MeovTUwIiuA75iT09VcygmncjN9tbfnafI4z
X9kR2mj/GRCP/DWXlPzYMqbz4BtggTJbREio6pPxbbBBHOKP0nywfaSuSnCHkTCd
HIZkPy9EQXVjNPZqeDLewceNQ93JtSXLiAE8FpqaAvqIQqZsOQ6zm1Aa810DK3N+
fQeUUTvygMrfH828zhdslgAxDBYVAnyVlS7z+GCTQF/yK9X/xiq5+Dwau92QL5Zb
26lcUvHMRtMUF+tYRbe+NtEUqhYxRu9AqIW/qhmZyc3Zg8RPBxDVoafF/r448r+E
Upzi5Zep+3n9mRemsIVWTUVYTGCjacFDGSL85edvz6o6lNC5iSjGWFXj5ZbNhPoX
VPz1e5i5gj85yjy9w1Jh4+Q9PBTloMVcQdYQRxswrVtzex0Inut27jFLOGYyUzHX
Y5A/LDj9zS4W7SFqypw1qrHsV1c3IdtWPqjIRmEa9sWnNcr1AX1fFggQldCCV/4Z
Y2HcGTKDgzShNhUpjIuO+OeuA8nFMXu4vtnyWXbdNVrFRtfeHA22dkz/P76wCKtJ
gMcdzRC5VQigAusTGgqsiadiVk/H3dASD/p0K7jzETinzvGTnYRj6ImxePaNqDCz
iPfLaOX9zgnJ3RsUCAK7oQkRytaydkCZ2PUdhzwj6nt577C1FE0KO83ZghijQGe3
WJX48MeIwB7OZMB5tv6+xb7D/7LhjSgC6stCtBA63lhjmpuVemHZK/mYveKJY3mT
Gb9t4n9J7lkMnmOg3QL9Q2PIYuDuXBmxL5jSeZIRoI4R+i46wtCsZTXb3LGY/VE3
K6mIYLvHWVUhYb9us3ASxULtRq5KNZ8HPHR7o4xg/Xbos2HQ1huttb0jFeDt5wpi
5s89LHD5GSgw1C8g7Gw6wRf1LQAgtM0MInZPxVGPD3U6iiQIcL9elk5mY8H3X2Gk
63YRxaK1YYdG5F6ronGnb5S46hzjJ7eHlTSOq8Z6dm7WDa/93t4GdHGoSEBqwyBp
/XUDIf4onl5ygCUSxJWeyedm5/6CrCGfOh2dUqemBPqVdBrKop4VGpcweSU1UVQd
VukBJ+tXMI9M0R9QU4MLfNJirl/X4pTTmmUN898SgtYNf6MB4/i6kugYEY297fDy
MX3abjT4JfPA2YuY3f1OWtwWpW1yiEc/GUhTqaL23BKwCXQlMKfzFndXJptnNJUP
GtfFw/xGCgzQz85YyEz+8z63L/fMtRe830YT55xjVUlHSSo333r/L1fJPl6pXRpC
0HNyGxaJsoHn9g3pNPBXmI7h1E2ltJ4TyzBjRDvYIlawXcaNvNQ5NojA/WMEnWdh
h8Y0uy7eOg2bmXjB4QG4BVe2SEUpuv9l1Ej95WEPenS0EsSyi/I4acwNipGfn/Sx
KzDcijQtY4p08+GhMr/MfKSdP3zMNdwdJ1NPi6+Uj7GFyqDkPb4eyjQ0K7aL0Fld
D4o5ADqPUvAnJwE1KyftzOtnPfLpyBCz0P51RIpZWgVH1g96/vM4u6asdg7RXvNi
uaqck7+cF8dm6+PUOTRjLntPwxH+ERjyl7T3ObwmrqGyakj+djMSc811c9iCi/dL
Xxhb6Ba5Y/1ExPUGvkUIyZ+hvggye9lzVaOHZyC37FBwbGAjl7NCflCHyrOnsUMp
1uzjbKpOR+yFgLkKWK83x3W9D6yEValEJ7ToWJm4WE0wzmQ8Ypi3sQFJe84Yc0Rs
Ju3vhAUnYGHo8hJXEsD+97QOq/AQ6SZjRmgFT1KpVvItkxyVf9CFzzjs327vFX6N
XzNDQOO1oVQIkcLKw8ZJUpomhvaMNW7dz2wzMCL4J36s9+lHh0+VzhnxSFBqZ7a+
oKGWOxeocf9RfeBqOY0fD8rp2Tz6tgqhVFntt2jz95ZXAgrHnGddTVL8vjmdbmDB
4d8D6C1Q2MlBbE8wRcZZGtYStL+xc162Ucjp7wUfCp1kkBKnA98LTs12K3zp2zUH
65a8pNDs7TuGV/KtJxquiGN9p/a+mr7d8Zr0mRCmsQLLqw7Tv55iBndOnzpkQroZ
ylZ8H6PJipdeSgqrp21e2JK22ns2+5X65M2csNO332xGqp4KLCbVwKSQ4Wy1Yo72
/p9HxENZahEWOJFvZp+cKKCz1h9wCIP1UUOynzbOZUJOSgnTjXhXjFjrBXhBnJmN
IXWy8gDTvwtqWdSyH0GRREesfuGaUE3JbkZ7xv/JY6CLn0mLYz0aIJW9yFprFYuF
qzCFV7ZpoXFOZg6IolUdWuEPHWetNmwJas+VUee5WyLEyR03iP94la+VxXuWvU1G
Z72qol78NsH0ESiLWDaj1V+Nl9igYFseHwWftPsGOPJtY2mK61+T3cw4xQpYmwAE
+N6ROQg0aQS4KjxEuLaw6aZmixdsJVEmT+SUVDueW0U+NmlrJkUKKF84WWcqUz2P
pVG4Hvbf0tfYLPjd4R70uwUoDIXHVowpjEpNFDJJrM7AuF14OPAFLuSRDAb6Kxjn
rJNxDTDTIra13j68aesofbr+rWBERGZUhitxw5+PMapfKpqNLaAS2h3kfim6Lxcl
/7L/mLtyubo4yqrZPeYxnE+PV47lCuvid9plQLsNmLi9JchY9jf0VDidhoDS0U2b
qanllXxiEOAOQTLCwmA1kw6n9BQ/xhPVNMrBwJBKNt5PkN/ONvkM7Coi6cDenHgZ
L6MGvYxWsjyYp/G0MO7ixonxhTh94exMwWVSlEx0bKakjC5iBMw5KrRH6Fg/JCZO
ufqrVitAJ3myJNaTwbxlsk4eccVGboedqdgQaSG8DY5y+8ykZOBq9PDAscgu18NC
aPiOBWJse26HQpX5BYNdHaNY/OZGtuh83FxEFXzPn0Ie8YCveY420g77zLb3gNke
s8y/Leax+3cUS0g71fw3w+J85uwU6hHGnFUCxYpgwBbuNbWD5/P8FN7511I/wRgG
PZPEEtiAe33tlo+bcnkVnEfyHMvtn06d4GNdOBloLvAIbSvQxTIYnkES5NMmPJWb
Vfwvy/XcP1k95wi/f3M8HIAlQxKFthyqqfn7/8awJZvOPNH4sZ6wrSONgXrDZw7w
86eZbFdjIoqtlINgn63wCjuvRB/FQDgw+LANzDIi28N3T5GhGcl60MOFvtX6aS0z
pRHKxBpfIG9nwrYIpwZ5L664TGjjskFtp5Oo579s9gXPxtkHwJZqe9tVIf4OplWY
pRGxpdJTjrpU1EF426FpvwzbL1PZjgmSEBzCTOpBd9xJa7mYX4fX2rYRWcLlPzA+
l9kR1a2fy3vHRRpdPi6/IzIPyf8COg/l1RjjTQC1qDdwIlwrmWqZ1fFNsD+iMPZe
KCAAFl/Tv2pzR2++utFZGWSpbfuL9WiDM6f/xIxnPkYa50/ebapsb5RT968qkXrj
nVOLLXorL9EAkbfki4vuS0e9Mc0golsrZPJ3pAfmmEO98g5l2t4saWa42Z0w16Cv
o7osAkUwVfEUPP/yfjV/GpzDwqqXFHklf/d1oBSte5MR5m0OQ+5gYYUbZZs/pJK8
bgTLp2qUZP3wSHG8PzB3eBB3vr5sY2fP1pHQuIXnYmzuAbn/W7gw0NckANFrP7Gw
q0qCWdoEPYCgrEWHEVScxdfJgs0N9Yx/eZ/p1ug4shBUo2OIJc4ZLsxbCVl25ocy
P8BiG7XWq9aKnNNZ+iTbkK6oFIwGk7juCTTBZ94a+L/AlEVqYIc2He1CpGhj3jEH
yBOSMMpr3+Ra6OMyuS3Gxe4mnAFfkSZaL7EsACifs9DdcHL/Ll5q+J6fvjKP+zAt
JE5hwJjMBYG3xkTTQhcW8eSvyrpzGkfeF/h/SOuol3zfJ4drUNFrIFKtJxWVdoZT
dVSlthEsbOL4qJWwuK81kzYOSVbuw2oziMpkTH/lKFEsCqB6QVftZawqhJWl1mCg
Q65W+vqWxh3CfWcFPcfEsi7uNUyBxlmIlkCUyy1ze/Mbd3Ki1i3wO/xaWTTNpf8K
+CtiiDPZFXAX70tiiTPFTriDAyf2Utenx3V8EAyW9ybBAF86x70ZQGdKW9wDK5BH
dGOjH6z4Acxhq+g4hI0oENhyG+wN08e29plo2u4TK5L4pe2JfvDUXfn6rgcFmIJz
UTzl+gzHOTo+mKBRpL8eQmiyE/nLkpL3VeXzbGLb+Es8700dJengeN8xTTDVu0nz
UEbVq6oFVZ34BrfyrwIK0HuCf+lFbSvNfAWnoiLIGc9vJPI3iTwsHS/qUQadRNiU
mzEpDG/qErz601Gt9I3fJVENfyrmAZcc+i1eTNAY0pcX2rlXHTKK+FajipXDBlfs
IPg7MkGjET6Nu/c0DrFgmVzfCIQUJ+kVzkAZoPTPMYdm7IuflfMg5v1cIQ1UJnRE
8NYHuQYdWw+K1kFgk6fCHgpIDP0Biy+IG5fJglgzsCFVfpHFM5XAEl8tUCsqygnd
API+y/0IVYrqY6Yt+QHq/ShG8WXmp7bDbtnz4YoCDBgDvKgAtDi3AiFiFgW4bMZm
ZOYTEWFxYLCnOi1M/P8ix5MPt9CmC77EslpKSjaoiJvnLEdZKDTmzS/pZJUMhYHu
cY0w9UzaGKKf9KNImS8bTSPhpiSzy09BZRfwTlJyG3dCDpLdM6RLc5W/xMuoNng1
rsw6pLqxIjtRcer5gH3N9AcW9+MD4wysh09+2PdApuWW66BWikHtDcroPtmj7You
J6+2vv4ov3yVjgDwi1k6IzoWBQkNVDZoLCaQhMFASJRvtk5fTrSMXUpLJZlGJjQA
UWz9jmAPBaqauSDPPUedHtUiklLC+ZgD5chFUF71g8wJvAFfZfC62aMJ9zjCq8z2
hvMr8+6O9gJQloER9zCZciqIPwIlyoqMRoow8EdYRnW+LUBqn0b9BUgr8YAXaP1z
0hobAj+Y3b9iNn3o+23dx5arxVDoiuYpUpO8qfbWE3FILSbrX34U3Evt6rpSon40
cmbQFTn6Xb5g8+rTyNf2tXpJSektCxySAxALZzX5IDvuuqFqwRkmiMVuKYeMdN+8
IjRVAzACFcGQdhMl4XHy3ln8KsAjZ0L3gpiogFMGT8ddSsDOfGxXE3sjKlmdLLk9
nwOVKp/vFoMtnmveTB6lzW9Vfietrijr3NBHjXwCxzZzf2y0cKBi8E1hJ4rZldYD
zUIFtyFEOXtuGDUZUAWDWVPxjTFUZkNHSf0sdTPENah9M8wD5TinCdlYepKayUol
Rt/TR3OC19HpVuWHeFuIZA3ggnyma1yQsexgxRlb2qCKthpTMXiYuiwXQu1STyAt
u67Olm8emC4Zxc7GffouGpQ+VwBDLMxiMu6cS1NAiHYf8nxGTAfNrMVXtCKn0D5+
ZNRBmDU12Zs51Q6cm/HWMR9A6REf7KDlqFTPrp8ZOhHf0l3fzMkDAYL2thSz7sgb
yR2qkKx0rLUzm4krpdnF9llS5T0sbhwLmcm8sQLpynyntqaAxIVULtwIuwCRF4Of
RvBGTImTIFDqd4Ff0CvecNErR9KxSGyxgd/HOUV0FtKTA82xUMZemWsaC7qfw/Ep
R9GLaxuyIKJVSZAxotqigWc82FAWWAahpMuyutcWwJkj5IA5z8/PIFYAmCaDygYv
QBFI5p8zAQ93AygcT/Pg6vGLuPXd5/T0d7BvGGFfTL1hUmWVfA0/c9Z5U7jeBssD
iymgIg+8kbg35o0ehQ0kXxkVYOetx8cVlrCpEDlfWMx5PPAjxjjaD4X0xCrWxgFT
8WaT+ApAmCU5j+2sZQiI7m0U4t+p1SizxlFx0tpClXwg2/++ndN6ZSvR5UnmcuGI
7Awk+cfEYC5yBnqjIwwdDyUtX10J+5yg6mDYlAj8k7M0nNJQUbUGtttd5xBfQpZT
dbmegTcSp9g4uLx4cIEysuDB+wkHTQfqiGbZYd5zkbRTb2QYS+VyxiMqp2Q+ioW5
KJjKsP/MeBPGvR1lGR/8t/wGkYIRA+N20jLBB51NWFpl05UReY23KznnlWdDZJdQ
jdeaxEVF6GWbhHaWGsgAF1aYwCoDlmUIlbUx+jXrRaTjG+FMEnmZUWSIFiYJC3Bx
gWpA0VrQRgOEvBrKtkxSmNVV7iw008jJee/Dc7aojA3q1i14e7yFWPCedW3EgzlO
n2UU6DtPf6OQ2YPu5AaA/8XY+Scfy+YaH946CBb9mhT29SyeKxoQepmYp8b5kjxl
GscPWWaCPU2Dxi/OlFSJD6QwqhN57EYY0PtDiAs3p7igXZMsAcA1lqlpXi6yRgh6
lrZXD0BW6F3A0juvvLi6ripyw056NJ0a6qgDHBcEbuHEOdkb9d3jlN3/KmFTiQum
1TwFdy1VmYpl8rsJZeWHov/R8NhOowa2qXaQR+0hyTJll7nF84dJNijb56nksLGf
RInza7+D4BEZhx5xrvZwzScd0gX/BV6RM5y7LJKgnd7xoqUGvVJZ7+sD0moaEqxA
qToFmhRLlOO+M9D/jzNnps73xQntKDzzDCAOI+wKeKnt6DCgCq4fjr/HkOs78nP9
yFGClhkxy3V+f9f/hJRA3wcpabA21nNuTZ3GrQI3B4JKCQDN1rBfNOwtY8NKPt2v
4D1eOCccQ6aeaOR4+sB9ROWYMA21Q193YLT2Xb2eHCvoa+ztAGamTdxCskRssMXS
iKs1oyPZKcRvGzZ4CTXFEvi2u6fb0GAAE7+P0XfDZcuwTkZwNT1omZS05vaYPyDZ
M/1+VxgshzbeR+7et7GPXwzvHEj18rb170NLHiIGcaeB9s7R5LAs9gGVD2TNZ1pv
qRjN3S+4QRjscNZp2VGk1Y9C6CqjM330uAbyZbq62IZPWkBrQ//V8Beu2uEZSSAl
tYJEiq2Yn1tWf7DTgUFkkVBr91yLrqmJbgXgq5aUacwo7p2kbC5PtWtMWTV1Ay+f
aL8V4QPiFEWKmw6vriT5tvFgAWUP+Lo5tmeyxXTjQAXWOQFaU1LWq0wgTp6v3YYr
xmSxdubYp+OOgx4m/20WEC+/y1U/v3TQgxdQgVKNiwZtaSP9LYyKs9V/sHlYT+O4
1ZOR2+P2kfWJ3ySG33Pxw8YHZyOvKRxKh7azeXlW5oIxa4y0oxc1Jlr85iemVskf
SOu2Ar6DUK+U11rNV5nSuGZN3jvjuSxFJAxDW8xuH5xmVt2CFD/AoELD0jdnJxtt
GX/ciR0Jj1E+fLD2VYJQUybUDmGefdp+Vp4NfzyyBZAv537RE1cocXvNL9EL8X6z
Iza/d6cz/STCty0bZIvHdXFCtv0M7iR815NV7ox/ATIat9AZugKvs+JnZkBuW11H
Q+DEzBF2tcdfeliBc1KfunOyXwyNyUOne2IO/2QsDykJk1IIM62CJDuh4W9Ny8A5
h23i07q6nqpSs6tnLaCSwT9oBU9iFDXIPKhKC0vcfrlBr/wBLvELuZVo9zapuPHZ
2KaGBpwXQQwDb+dfCZxfIzoS2W+DKCDrvrWNCbDcDuH3CHX3xvEIj7eGJUJ0UHjs
i7EHfbhkun3I3ZOVgAbzmaMr9Uw8Yqri4yHpyj7Hcyte/4bJ3juXIG4MfCVyk6pJ
npF7ohaaOBuoelNUmP0U83EvG/d86Hs1zq4+NSXdVKfSKgd7qlc+S+PgvkErAtCg
N9lSpnNOkXjTb6ApwZFQd3j/TURhxqrANR31D4ni0BLOYEe3h3YSgqgJsTvK5hAg
cxircHekpz7ZAuIWxWz+xNDF6OCWiTAsSnSu2LcYDBdaipETIs1g6LeY0VKBfUq3
2JCM+rCK6qFtm4X5iiq6q+DxUhhP/zbZ7Nr7hG/PMQX3lxbxMWWCOqq7Ke05dgJ1
tINzF0bMWOwl+LUiFgXXp/6JfZHa0yXwls8EhZJ8qvZZmktZWi/G2gYaGTrJkcYw
iq6QWgu+/B3zk8EreNYZsr+4jnMHXaCh7G8A7OCKUHo7tJkF3SKil0m7pinTvJQ1
TUbcPI2Ichm3gZsGdcm5KhI5SjaaXXbEhJLA3gMGeXreveG0GFuhyluFMTusG89G
2GhJna3x0V+A+cbMBugyUb/fDs9cPWY/QriHGZmisNoCaJ7g/PHpukvX8+JjQ+BR
MABoPsB8F9H7QTyi1KJVgSQOnz29zJth6QpXyiu9y0fBmEiPW8SzeQJdv0kR9uPO
TI0MQh9UqKrAbUDxVl0oscWP1k4+lc1Ce4ho5PqmjnH4/rQ65TfufT6GpFjE4nlD
SEsimun4Xs/HY7J9oFHtH4nH1LgcbeN2L55YPbeez9VGaNqLGbndbxLInk9vbBBG
924hGa1+8pvC6zerGsADUPvEhMgyEqhUmMshnaT8nn+GbPXclocqaggZ0p977K/F
/dr/c3micllZIXMX/QYI2WADEf6kkj81mWa4PRS8nU6mnQWO5GNPp6sqG/JgZAKe
skWdXCWfc9QHwUzOWS0ZfUxHRVBNu/dvEy7wN9IWaFGWm9DB3Qevdl1Zd1wewAjh
YgtWEn1D3nCl8XiqSp4Adx0Rys82UfC/th5K2lwINnQX/jwZSTKJ/ARV3PXRDgV/
tNAq8E3PtOkCDoKRX8tTG6Et9xa9ZEFekgfJqMdmyi1vt0VeaghUOD5l8m+jLqN3
S0Ext+tIZZm4MP8qG3cBpBRp8eKvaHPepks3vHpLrJodf3MC+Ajb7dwt/9NnSbiY
h2HeQf1BI6HSCVadgAODIGoUX3SJ6tU82tSejPmUg7gKR9gCUaL7nH9MXainBjH+
hpR/QRWVPqbxB5wcK4NZ3pzexp9tVd7DyhdCh/iHEnjF1kf0CjAygpnrXhRnLDV9
6OPIQVXWX3gHa3UabRV7z3YOdVQnxS0bnBQSTxzOxedkCqEkdSPlS0ql6pMed9jK
IOpoKl/maHECI/PDXkh1UV6fCsrlP8k+E3kP10+zNuZXsaKsPux59d58ohKE9lqf
OwAGmqGtPkilZdVEQWZlKl3XTN5QSkXHrGro1Ffs8hjqi2fErdTAySmxBX0T+172
TtBfM7vS+RGom1HtT1auD+IQ5U478yQNaF6Am1CoYnyAsgEnEx0eJtyVX20t1v4B
FFxWJUVzemxsK4Co6/L6V0Z8rFcgyOpLMzdX4rfzXhsxI/Y0FXZnPkQ8Lk5VH8TI
VJbzlJX7DjhStUEZeMP25HYG8anSSMF9huvVwGR0gQZ8sRmLxf5Kbb0qO2EM5QGr
STmZiYbzbvhENsnBGQgPXGtK22+xLhW/x87cQd8fM0lKs+Deu4VImgUvt2oYx6Ob
n4+ecg6qms8uSqWmFD7ttJqB69rBNI7D552d2n2yrVrCsfqLuaT6Zbm/oSHrmn7T
whVchUa2aYFfiSymGN5LBwHMacRUIqqvcP9mshiaih/nwwSuiLtCv0JXPhxfEI4v
eCsZEi8Cbbxx9gdXIiMx+qyghvr/PmzhUeUjve0NxCttU66oTFI4DCGGWOCgb1t1
N5LrIlgbd/20hNmSArSPd69wYoBLdcCnvnAM/lx1UTvFZQtLj8t2wMozM6R84Ggg
z0hrr6huUy65zes2nq1w80VZ+2z0AiKOugwTNljgim6Hxp2R088lTdFJHkxpKIw+
IC+e5cQfIMvrZadNbKwW99Qv534WYhGiMXyaHVfq+sblaEBf0jtqlIIgBYVOSc5G
c4dMW9smapbj9LMGQ6jOGCVHDsv/npTugS0Cg6z/nO8Q5lEM3qia/GIEqo+e7Cg7
YYE5xfrAwRtZ3l4jysTjZS2HepdYiMYHnlrXzwnlXohPbT1nsqLbta+Qq1fvZrpg
LvoUwxrgHGY/gz10lc5SCHBzjCNPMCbHjvXgQ4XeZytg+b8mUR+D4o+kJqHsCr0m
VwISffzV892O2vas70XwbTO7iTpwbWfL2hN95FX9mJXOQeXFUsqL/nLj+Zfn9P2C
rRcpSQWLXp8kNzpq3Z9lxFMAYTLuBS4pm9i43bXV8aJFFHNJ7cb6udo1tv9n+r5A
nY3PnGAv7X3CJuR8hDth+ikqqhDBEQn+mqm/nMOve5wR4qXHwie4WEnLPjYFB9Pk
X/kf0d8GtUFg9iLHvIdpPpzSLXZWlkNMYemIJ53RJh8RHG+ju1z8s9AuV/mJfyzZ
oRufY3UYR7d3xT4+TOYlUh2oM6voyIKK9Wqi4zWPAVRXcnNFSljEF/Hc1zF1dv7t
8d9xScrPXOMd2ZTfgt+fbnKAS3gpcH8Q7UdDwEiaTVRda/KhkHLXBvDk/Pm8YqkI
aTYCUkC+fJhl85V/hoiIBSGjeIN4FYzi8II2nS9PvZJAGK30926bfnI8B88Xsh5F
sPTNEAKSoXMAm3Sh102ebGCEcD1u7kKm/O179vsQ0VbJAT49WF9G/8EhbGrfD9H8
WfXb2QFQj/uuJXJCerhaFDklLjNEstbyzuhLSA8l0SZXCRYilaNQ7NiIj+qG/Cxm
YF/d1+9YHDu1hS13s1r2Yn5P1XqMHUNdeHjIgtr7kUpKlw0SHoQ1yafj6/JPoL3K
Hb3kIGgXCzfUV9EYmGXB3ZPYXAiEq0vzOYmXqtCFsqq5hLfVIyU7EGfTLKQt5/mX
CuMO8BPV+/o+SUJg7GsncgjztNmwH5rmklfjgXCleaJnDe2PFxLa4tgjkdjlQojQ
dgnS8ES9Vgb+e/NqbR7CF0p7+VxRb04BqLhFmscDyw6W9hY0nymj5921VhHcrHXh
xwBnWdL3nILVXn/los4I9NUg9HUBdBZuJedwyRQcNLvvioHaN8XKCuJkrqAE3SRi
Pu4yzeO+d7c0Bb5JGu2TLu0qGsMUwMFXoRoSKRpDRjPxjaE2+OJD4SfYnw+14D/p
8ZL0RBSSDpsHMB4MsGkoBAzN/gakVuUV+X8l7r53jkMcoLdNjz7e7pL9QaCnkh8A
PhOZNtHKRwLTl9cD0H9YkEa317uEotq3ff/xK7kXuRVBIuSPnf+q6DVLFCkqJkJN
Q5nO8kxZPtVyvxwzIS2uPcaqYdlTklHOv26b7emoA4sG0mto2fQkwhvtaLtDL6KW
KpiuBJ/nr6JlHV8akU9D0TDhoMXixwsewJyWDQ80MTQg7rjqYtpJWeqlN/r2oj4f
A93CEb5wtLjwb/TU654doAR8BzMCs9MF7RcipVlAweAXTGYz5NDXIFNz1vTZz4G8
/MI1xQxBuLuJazpNAOrpTA5gVcWIXn5gr1wth+AalVup7ETCYsUHnFT5fIPjY2k8
2EJADBaRZA9jgFmdk+CVuSrSV38Exu+PxvmrBrSm6/HkPEQmkmfPlCgNGddic1wm
m9C8nqXNbGZS8Hx/q3gjmWWFjDMxJxHM6qaCbrymepstqg0ucmBU2z3XCrNBmj6y
A4nZG+5OPOjLF12nH34/hRC6ZgRHXo76HaLZlt/D9ikDXMGCU5Ey+e0UznhxcqZF
ovDScrVHgTi7+n2sl45eoZI+IsqqGAcdOHvHMmCwvv2ai0tSu2a9B860v13JVo5A
6gFFqIJpSnRHJqgDbtE/COj+/LgI3cnQLSOcNpkhzlK5d15K3ZVfX8fo7386b19i
6EZxOOnex84wXym7ASdM0h3eQTFmZqRglIYjSmoS2AyOYI9aN3WkfgIpr0vDtmZc
Mue0xzVt39J1T5e491/00CExD3vXGUTuhpZ5f+IBYJtjU6Fs/AzsQaOvkMP1kk0a
i9mjGxsfMiahlwyCjKlmdODGoqrxI0AG82yLKdxmzocZ4EcHlBqiMSO2ZZRLJtDC
uNvsgaTSiC+iMG8e5T3PGZqImk64DziHYcjetcmqX6C/k6iW1t+xpXFwRs/X/PQw
SmUNKUSBlvj6c3isuSQkiHyXWEtafIg5TTE/ZGBww6nlF4WHOatD+yrxkpNod2DC
9dop558bFufBiGNeSbHRyGJByhHCOXRewJ2bNJV/dzTN9XiU7c31SVUqKia9STYV
V0uMhKd2AWbhxZdrfWzKFiQ0aPfVtWOoPqgVlrUHlBhBpgKqWJUIxEHdPgdCBsbi
LzRpaCPNnx0bF3YFexJsBWSOY7V5jNhfme1xorwge6G53L2tKsYtv5dFUvmZ4+H8
Az5l0gM/4cbPJIe3yb+rIMaBI9EoqoLItzXqq6xfEirHYOXjwpEcHwzlomhqYqif
CNiq6bMY4C4V0LHssqlWBjzvBr6s3Nco0jFirmKd6OLN4IuWrFNd5ztzzdBAN071
zj+fy6SIinOIOhu0ZTlmcOz6KS7oZSu1g+YTu4QqZmrcfe36SKdOU3hqtZ6qjaov
cc/C4F6NzxeqXBEwwKcrUUg2/nMr18Wm18J7NwdpRvhwBMaEzMFRDXiz4zdt57sM
fDj1SVryYzyCr1G9yYi9outgF1ppp9xrziFghOdDFBZtR/Kv+7BpQWSh0TGtrcna
r3nR1In9yUf5JX1JtgIKfOIGHouevgDxpSnkastTzC4SIJaNszwBvNpnNJiCIPKE
WHSkf0Wn650i8RUmYwNCloJepecPpGAhOhNguCH57uvXZvExMi4z2EkI+RHcgCM6
nhypz5vDDfpjH+UfAdxKJ6dV0YvQcEWUre0F899t81Ak8sJ8dVd0DtWU93je9Lm9
HQTMPCTB6l0fSfSfOQWzoIVVg/hc2pZHiZrMLQfwRNynUzKBB0I2RcSxnay5DBoq
rZRSoANuOx/0kCVVXPp/Z8xgrP6AUNIhft7/1buJBiXAewOEEKueJRvfjv3NcmUV
83u3Rq1TAoHkouBvx8aYOxeOqbhs2vozkRFBc2E1KSJMOmXpnZxrD9XfA6kN8Jw6
4CYQC3xufBie0il+6AudbpfuanEfxgpMjUkIgldTttheQJ6jNX04jZxUY4A67pto
ipQNVt9RZugWWPwli/BX93Dir2qzDGw5rN/0JAqJ0A9mwCyHPnyuj+/huV++AJej
y9WZCfHM4AJMoqauuVt8EUCpx/CLHS67+A3wiE2IG9rfo3y7yLvSCL9eRz04D+yh
oeHutXRxCKnAyq01yQGfC3u8ooy5WUPF9ki3xy5C8Z1VNCs1h7s4eu1MObs/f8B2
UuyW9IZcS/1VezEXkgXMm3v7p2NhNu7d52D67suJCx/2OFW1GjtSVhIwdLN9LjS+
CeSNYJhiCA//AmBOFWPxxjiE0Ma5zwq/s9BF6CsMo1FSgzZKdUCHv23hpqMr0nFE
VYXB4yDZwizRwEADKR1bBPCVpD9+A8m+n5lAY++wlxgzDjZvi13bJkB0crq5zXXG
CdASX1wO4FnLlbuD+VQzrBPSDB8MMWp23NeurjuVQt9IHj121CFJsjK/m+zTuhvB
+ZkIJX9rFg9dyw5nelKnkaRTaia0oaY+g4kN/XO+xrMwQMn0hd+HE+h20/nnmWak
DEnAxa8S6k2Z5aM2pZqHzlNxD8IrIzvNXDvEb4URCKYuO5pxGBhyBagPXWFIG+x7
7aMpfYe/xqNWkRR3gXTtnOi8SyCyPhYVGOvuhZpqVQ4groD6LnAL5bROq2YUH9ZN
w2he5lWeiLDhzfI+cigBoiDbM4uR4LpFvMpx91YJ0vOA05u89kRWYgm9oStOhOdS
h0GyhbfbfCxuOTYvYyRrt+U1mCaoGI64Cy+NTDRSDh5kDRoYYbh+F7evBPaqXZAW
IyQyJfqLeIgW3F6ao7bMZz5vABjMI17ZGIeu5Q4aF+VhW4L9LFZxydXgShGt+f1z
uvRng0M55GBN9pnlPJqaDaO0HBAcYXx7cTkBprul7X6cnORUOgbVo8KBB12Ka3gH
QSN/By6cZjRdTYUbX2rWTtA8cGF34C6SJg9hdUbNbD+aaJpCA+Bbd+Sw8v85u/vn
lfFigDzW6WW5IPg4HmRP39W1CeataG4HIVGh5ffFHK2j315ozMvLhS4QuclhB4vt
wrgMeWIkHd/xWDFvCDqo4QmLnsRgt4lKU4ipK16ELOHtWh9v1EwRuIYSfvIez50/
eQ7EmyNMoKv27eK7NFfKOjh54Em1jeknQZIjQ9AhuqOkWvu7HS30xJ4EIKidRW1l
EYufq3cqivEQqEkXQrrVxU2mn3KjqQisB21BAisV5ttK+RMXyYUlvqsVvC0vncSt
i750y0oYYK9cG2H7/OUnzgzj35FNG7rEE3oGnASA+9kF30R8qqqawj1ErZOccaSF
Qk8ByBhqTSEuoaQTkXwaCsrjY/qoP0Hc1xk7ynybm5z4ZLYhLsIIaQlcfc/P3f2B
Scw1aKE4b6PnVhA448eYodHWM+waUrlBUyankmjOczjrj6rmjFiXr1w9WxOsHZQZ
ont25ckAe5Q5WlUm1l6MCzemS69/6wdnwmmNNSxRALnOPnMBH7s90VBqih/eWsQa
Fc0lmXnGhEXY6vRvOvmC3MVn6W9k+PiFoy6T3u8+uqa5e6GPftgRGwB3kji+/8JY
QOzrmsgfkBjo48t/YMN8cYAD4LZ8NCwtHtByXqshh+cKAuNStAx3IIbXtUwC745M
HWfAtkf13Zu6r3Qumnm1OFpjjRc34TF6UW6xfDssnLA9thz9aWBZ3GII7AgVUxuq
M5kx7uIVhhzOZnGWxPjsAPB+M/S7YNvzdnJdSrW6GEc4iaj/KLRwXZuaE6snuQLw
UgpJgX1QhQbx8h8HtNp6akU36hkV/kaedzizXXRBZ965G3U76iGNNVqGGm5tJQKZ
qwZyQeR1BfeqYpZURhk3dFc6HrL9/OHjyrQ6Dytuknl44LEJW0cyd6h9Y43WjvEv
1As93YqHND9sE/wbyj8txMVpLJMojvjSefT3mp0CBBCVE5qnogC0Kn50MbQxgStb
R8yFD9NeFNapJgQSzfRXrvbxol3sa/kgfCsAGmMaJJbwRgyqUHyp1C5RUdKnN9p7
vL5AhUgyIaBCfOqit45ObnVJQGVaYgNfzFeb2cQS/KUvUq64je1lgA7U+AEoFo8f
6ZwGc1B0pCugODvqit6dCeuF5orhxWCtPnwEnCXUeKeeXtYIdGYYz3gah73cdQTT
Tzw40papJBMpn1r0uHYe9xru8uBM9iL83d1BlEFpO+zwAthOrPUOZCzWLZR1Muu2
rwOPZWUjsk7s2jbbrxkUd/RbrU4MzluB2WjqFjI85AThtedEfd449WwuCpALx/Qt
SuP20TyCMTf82Tg0L1fpRupjWBsyddjf8a6HywMrVmvdsCEc4m/Hj9kobyZxTskc
u+nEVrryC3NgBV8ZEXjo2HqOK8oQX92+jNDx7/pNUqICECwMMszhBb3CjV9I0qF+
73VClWZwjiPFdsvWkj224TKKxdl+z0ZELLch5z0lF22IufqgssDNAnTwDP9aX9Lo
elHuUks17TLREJwH7UblZAxyb7kMGy/SYjdV+FXbuq/AWkH8TQBcv3J2Il9AV3VT
lDw11THORH8h+IxTLbBl1f8uIXDHcozjeJCXtgPmm8JAHnH/ACIJA8VtFQTgOzrA
MLCJQtodG1DPgfXajWD6f//4QtLkC7BHo3D6aUS4oXHQCfU4YaUnOFqJqPSsuDHh
6pM6nYjfmEAiz95S/VaRWY/Zt4YEiIJUYasbDpdaeDEu2wjisi1DPc5FIfg0/DOF
9uJif7EVNnGDs+BMa3yjT+3FNnr0SAOGFjmBR1EKnDPCS/LKNkjMf34svWy5JWwJ
7HoDlvY1JtF2q9tAMKAF7yC2Xu81QcrTg3CRUSJjvLA4aVIPwLy/jZT0cL7HRvJ6
l+/EDSTZ2PuDNgtzF/0+nmIwoyQN2vgIqLU7S58MBXHSt5Ff9JQNmzDnWa6AhY4R
2PTA7dc0NdkJgHg0M+veKeeTG6qaZDM5hXmLoPw6A8Bdyx4IemvHnHR2pSDVDe0H
hzf2+XQYTOhn+LGaLT80n5UUI+BfkIZPcmMx3+u889p3hRIRz5zfB6DVA5g7hkvo
NG5C/gXgv8v2e1Krq930t50MiT/zbmd908JcTrX7JeMDvkcP56ME/24HK3d6xfwJ
SpBKeFqE3gEdz9wWUuiSkpcy68+fIz2HFHfi4hXSSoqYgtUoKslfExmeD/TrT0x9
BVpUiXWntV383bPamcJOKpDe7uCcQh7ayOpUCCkMkOhM+gB9aKaDc8+sGw5gTQry
`pragma protect end_protected
