// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 03:56:36 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kzlrKylbrdp0Mkq0V+DQ+/xXUbNrX5rMkh8WHcSHVTuOKgTcR+qdV4kfSP3S/kSA
cJ9gJORB4lv2OTAbCvs2aaDukVv/fAWoUWs7IBVH1Nb/kAZTxnX7KqbDekduvZnn
dAwlIQFLIxuPtalnuCdUAdAXUnC2f0ZAgqD36UBkqm0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22080)
gO2EUFjTCkEokNO5LLghXfxVt3gzZoBkZu3EKd/aHbivCuuNanAQ8V1RouJR/oIP
CICStjtIsKFKXnGghgKgP7cc6aj22/N9PvRJXhzBS4bnL1L1Xlu7kBGrI9w+bNHN
mt48vR1GWy3FTClWMCIO0qkjE/EyfbfmxSCJDXE2vAVdSaAI6KilIiW1E1dAlXa1
cikdiprtQOwfdAWs8QfK0SotOg8Sfsgz599xxiwpmUN+Y0I+q9Ghr2Sk/TmyWgc8
1rhOp0E9m8TCgbcnSzmeY2pyZcqJc2xpCaTtexIfHg9PxcwD+sx20nlQBBv6AVjH
RxeiKEKDHmv0thdr2x9JFTXgeItV3qPFOMQnrhT2eTRh1gFpHvobAaDydS2sPP5Z
V8TFb/w5Bimkr1zh2gsS8I8Yj9VLAgMEUsLresGeUwlAq+yAMTR71odWUuua9oOB
QkyPw3uNFuByZJnkLfd6BALSSaSah2U38t80Czq9QBKxMk41lMSD8uJhrkt2sOQq
lHtSHL6zSt6RnKEDB7n84HEPGXSet9GKqKRa3Q4H6biUl9Ht9B5PTrZp79sxSxnE
ovNCM+Ea67fyVgF0JUDTKJTk9iuP0WbEpqffydGk7XFyyz2a5rcIfRwotwxm+tWH
5j5PbiTrzJ8dYm3Lhlllm0Xax96nzLJBUnL10gGplBEzCTu4o8gEpCh7RbvWtoHF
973tej7Cojyzqnc5w2qx3LdRJMMs4a2yn4pu79bVNFLzCLSA3UzybauSgZPRkPru
AhNYBWuVHSUjRZzlU1krmHa74Swljs/6GH3+ruZTs20Dp/eIqdOHjRKeOGScVc/z
QIiDfFBlwllZ3mtVpQ5WG3aoV1uX60gN78+iRNdFzbNc0wR2USzhfJxtyPbgMuNO
emQBIhvAw0gJxaGMr/wZzjPs00ttrKmVnFzGg/yELTFgSz96oDjeZnrhXSHlV9Hf
TC4fnKeBYy6KGIe4UJxnfaOPOOWkhzlsogOGxjVNbCgq/1cKLA4RDpf1rNRLcGRV
j5Y5nnig0VJZEp/Jjsj34jbocTvzU1zPlniGFMwPacrvFh+OzkNUlSBlnvZJmWGI
xvqOzz62nyvTst5Bdvmc9N65HX0QbIMWb075Bg43iQXHtYeMU9cY3H1NoaupwWse
evd48N9Y6O6/MK+6l4F52mNAie9yYqtzA/Re9D0eXkXvTIiw6gD/kBRGEmIgXF5C
jqCcDHal2lk4suHiED/QXY0OT8Vb9JqasPQSObj61efFFgV+ztxioI72Cxwkz7jF
gOPfP1U8duZQjc8lvxH0tu6NB/y8jiX9zZH9tNnnSuq4ooabzV4m8WDFlqPc40e9
UpPX9Xw7i+KFYyJ8tKsd+QxYKV1IJaGjWpYSuCo9mhQZE27ED2mCMtfdo6Sb94lr
0Ux3qB1fGozR7z6XQa/k9K8emyPixEchv0qZp3EKvueakQ3VKGyUBr/GEOPa5sk9
ZAPfPEQraNhJ6RYK0/8rhzjLyHzbAhgzc6cEbpILum9VC0GPjX1JI5xrBpjjfWN0
24BXVrPJ7QuhbcVzlvF2Eexxi3PxemNANnpMdVhDInqGCgqKeawfnuta+d7eS6KT
VUWjNZSLCZjLSh+UB/jAhdmHKdYzyTtVjWVx1mnnAT+MtYmuHwM9e3TND/uqYZUt
ICF62p3w/18/hoSaqltP9Wz076K1KlGj2kSzqZaejWA4mdcEz6C65vBOu2MekoiU
ZDiuf8P83lt0ZQHlmHQoBrT0M1DaOYMS73raeKxu5kwnyA9VbDG/E2gf8pk1tr7u
CRmNk4w4DR0Ooo/Ltw1Xn5KkIrpg9x5WAt6SxV0g34iJfxuC8I9VerC+Fh1uSgoc
Gppurb3brbRbT9IAvF20qE2z32mEhphGCYHYEPkRRa8Y8wpCcxr+zLQhP97b4PmT
fbj/jqfxaByjBPd2f06Vx06Rf+iDIYtVeKOm3jb4sFFsJmMVHU898aUyCOysL/pC
IivQTI+lIhZ298AyC9zdsZiUwTfVYtl08pGFZe2uj9qeiyYtOvSz1sa1pReM8nZN
EmalQiHABNRHlgCfYjlPefvOzfebSmaFE9V42phiFgrWRUUmSmKMYXq2h8aVVcdT
l1+U5l1eIYmnk1mgC6wUnDqtBR2figFre59SZgF8fDSzQEexnkbpoZ6A3rWQ69lA
IhYctxXKXigPy738hJTbdDPFktNh65jUkesMxgQ4SCaqZ/0J7F+OKVS2meINcib/
q4Ok+M3fUSz1zqaVRcAcTVl1EayLky7UTVTxnN0pCYayCRBAbkAP7tccgIYRMrWC
tpJ3292jjrnn41LgP9Ug23Q4rqiikme7L7nrR4Btzvm2ihNH+SgE03RWM1bYrEQB
OGmddRyKOWfO+bxD7XbCUH0KotyXMpjZqMza9FrRXMW0hgFLmWaExWOpHd6jCku8
we60X7vyNZksfIbUr8mFqcPbWF6vcexjy/9+1kTAz0nxNikB0At1mJNXNEgfKAJT
AFq2gXiyKRxAMM7TSTUVamWEfJCxS2YwOTv8IKjv/AY8ELtZgKnUbDReT98K+BNy
MWsqfuMPSbTvFVah7JSrEz0SfmwqLMP/Yml20EoLxO88T5JI3shdBYOsvNYlzCGw
Wo2PAX605kv6uYys/TeqjWbVT5ZknIoT5HwLgw014sM4aZDd6oF0PHgY8FmVVHpk
os+mhsmvIlSDp7ZwzttD+UEP5uBuAWpm73QqWcUASYccqQ6yIQMY7HFr4gddgvxF
TCiaV9P26EDLYTWlSfxUaj1GrBADIlHlQYKp32HAYEJquhn7iiQG33SlpH9DWiXX
HLfi9sOIfH/NRVFuH8ftAAvqmaT/5Y+AWoNY6SHmluqZR90lZC3hER3CBUWkyznp
sJ7dvTK/cvyMB3/HjqhVsIaF8tctotKDBOfEd2yhYPpx2vkVyUPnZpSAnzZ1Rrfb
rATj79kT64RTk85QE1qNfN3Tgx8U10feH2+9ScBFl74hZEa2/J8epylvadC2apwP
L+ABF1uD/W9sWfcbzk/guVdQjJVtn8pAcgIImW2EuxsKjlyWtgyMLy8fLSjU+ZVl
T1h+NQjxqtj2WSaMDTgWiX0Cg/yOu4KgyxjdGnikqEhgkU9XeNhlNCIc8x7prf/w
vkcw/hwbkyIR21Qu0u9oBSd31RVcBpxG8wlJl9zv8Yxz/Qh4cOTO5mgpw6hMFrCj
HiagJ0dwkNPSnvIRNEAp1cU88sjjBr5g9UfuDct99i9G7c9OgXLtW12Dy4cjW9AM
Bw0Sdamkd6paAR0pHIjiQMDRe+Szhnr/9FdGMepZpDKnoc64eHs96hJe7nNoSPZE
3Qu+86AjdIFDDaqAC3R5Skwr5vGzYKyR1toqryOp6sKTlbf4ZLWQKvlmF9TtSpGI
VT2ABA/UttQXONHcFthF0+c48I59bMeQMZ/8DN15zyUf0THnlHjvhetxDjmYK+Yt
ItGQbfAfPEwnWKAznPtQn5x45W3nGeMfNxukX49m2SFlafMcDlYHIcyWl5eSWQ9f
jM78vCiduEL709/WGyvZKWihRN5PVEiiYZmlSceEO2+vEosDrhwJ7iZvp24cizSB
i/NnYJzUhGj8PdLeBEcWa84FmoVbLt/06cQO5609JzKB8G8FZ9zSBNaD63Fhj8nH
dzPefAAKV6r/0Yl0i0zl0MbPKel6D//zHb3vmhlS2ONXsZ67VzPX96YYU6/h1X0W
t2Wcf/y6RNpwv75eo6d6N4v7qXbjIE9KrZiexZBx9KvIo4dl3wkL/DR16AFd3xHV
4vlG0hEaDMvkejWy17r+0REaPVhj7MU1fKcbYI12IzQ6hrraATxbpWOF9mvEDGfk
p313B6C8T+YWRcDywqvAyb4FHp19mViRtvQ7Bpf7eK4cC4PN5lYEyVWrScBoa4JP
r0uKdnlC/a/i87+rxV6DuOQrOjaLGfzBsHZtFflqCC+BGZZOKfp4dypBJIpvLunA
Q+eYvXQuZoNNFlV2wm/sPwiMNIZjg5db1CNLh6nSwzGjKLga+tWhhzZ3DuoRPgwM
CyFA8Y2Q3f2UbYnic7E1xxIuAo5AxMUuWo6ZgQ6470rHUS4yFMgtBN6yOsXcs+cz
jy88UtRPDhkXUj9VqT9fjvqTJwiaQih9pzKrnMAZFDpHuf9DJwdfXDqlVDWHhS4j
ovICSerA7ITCQRforWCrOAJ41xkZkvyHQmQJQhYH7pV2Mr+0G84nHFZooX66iWQX
6RS7ATu9XAQCSzB82KNmDsW/e5OJIweBL9UOnj6tJheSOHad8YlLHuwk/Blt1Sb4
zF7mEfJQRPldq9cWbpFwmOmt1Z7FgB2aQZQnhllk1Gk1cWmsE8Nkqgu5tBS3AS8l
F1f9e9XjylbjINW3zjFe5YSTlK0usgES4L35kzmg9nhqhBSsz98vbJKBgzOSuX6D
JANoG+5gP3gDDPT1wNplUp8MQUCI4XlzhCUkumFKd8uFwKbeXW1maCnQpTKGr+Io
1TZZFWh6LeEO9M7CL53ipKasu0ix1Dh1NFnUbPmpQfTXg6wN0Nwm/3kfFNEvtXGI
IccqgNPrbQlCOK69cEcveptuKl3CGf8mEGtay3o6uwzPEKbveX/2TnaFVQn5nxKT
bGHT9vdDXahgf7s+Zh5TaBxAfaeBGHwyaxT3uvPnI5C72hbtJLG8Sidy42fwuVfB
j7vOlCSjCFddnBeMI8Kwyi34LBMYfBnq0OoC/I2zoHS/fUWHU5PRlUISOW3mIgGa
BgqBuMZsC6/d3zwheGhErlwOj0Fgo0nYaVxsy6E9WF2jQplojFqTN5JzcW60MQD7
oKZC0JotSHWnybu+C6ud+qd1t6525tmAJ3+xc2Q8QkbbcCn2ner9klgInzjMCECd
zOsL5odeE4HWY9tHfr+mbts1hYye+siGGLro9XK8tNhff1JdewT/D9xzGkZtCqNI
8JnOLAVN8Vo6KnjsSEvR6JTw09BvP+Ix0rxL9S5wSN2RT+eOneSWUkxcj5S/62Q1
gZ5vUB6iMqEK/tykoYJ8NShrNfsIgtMANlSFjWkhAFD8ZoqQyGJekIlAterQ5Vod
D+6N+81kNYosId4uHFHch+KIWygrBEGYuDEmC/77GCmHYWMul33N2YJAEOkHEbCg
WTtJvDUPvU2bPCF2OaTN8z88MzeoMNea0Acqan90q/Cln3XxEXsr9ho/b1SM/G+A
hPXHcWy7LnXNf3eJTvDffXZSWZcufK2MSaHgipL4OnWIjrypsKOCWaVWiDB0HKmd
01d0blQne+0LvABQNXG6s6ibdDLh7RKCFXK0Q3V9703hn8Lg0nB/vZfJuqZmsQMl
MX7Trt2e3ML7pZGgqChD3gvIExh9Qutn+UKO2kYpdG2bD6MZBRrQdJJnM9+2lnJV
8IYuroaUPmu1uB/F7kjw+cHBRXhcFOXjHrpnwn9HtX/a/b1eNozIF+R49Od/44QP
Roj4FOGvnXl07JCYnU6+uDKMl+PN3TJxVVf8lqy4MPGCm7NiGPfQ1Stam+Wu5yrc
4eRioanJKk3XoEQ9vW1DqkvjNYLQP2eBFHdl8c4QnjiNivG0DaCa5q4vOZt6zn16
OHOp0Vgt5wP66pCPpbUbNtBoVlHL+TaZjO9gJ3lPZwp2qniVJDdn7xxDTdi9TQ6n
wfb+qwib+WeKFUI922i16sLMelSX8ycEacgFg30ccOcUlmzzaoMRsfeMEqo7D/iH
H0Ir5l/D7GeS+f14UaSdP6uUjc91ruWJQzTeBrvjZECuyG5xbdPDtQjS7kSV1GPg
asT8nK/PeN93Sn1cvuUVWRzuuRYjPOynpJeYhR0OSHtiTnQKKTTF0oqGUO97jpH8
oBa/+tNoTtgRragJguZtfanjsatjwdjkqwIDPRD+a77AsHa4dAjYBFc9hbRHQb3b
T6jl6r/5t5X23if+PNYPKpg0dGM+jASU9Qmaj2+havLkvtaiSKdTHwpsIRwGi1DA
1W47b0gkeeH7o9mRaGIffj1MBETLva8KsIym1lhcA3SPYfbegnGqhMfKy4jREM3h
mtKjINM9j4W6G2BnEuYZpXWPW/533470exoIiLmCP/d8lIIYwP8LvnoIln5CgvP7
0EjBQoQXwtJ2pgyOLY5rHLi3Wz6tj2zfO4MwnMs3D7PIVu9WIhFtlYW2NyA+qW4/
BtQHnPWjv9i62Im8r8pCtIhFtvaiRCbL7c6Zub1hQuzSA8pXqx/yI1JBQnxPwExN
s3Nimkjoqu4uxIPkd1x+xV2NdHGPlGilBr8Ll/W1D0pQi/GgQ7Hgdn0B9vKkJPFw
CFsmugXmILj+fZCGbZNTXedjWLQuM82jXilEbNBwuECuIv7PUfET35mwOkxS7SPX
i12Wjrx4okVuKkaFjvVnu9EQQNIhvQ5rj7mgUeiXnz1WiwSHl8vISj+SWLFVxY26
AuHynV/1lFek2RaRL/Nh3lEDQGKTWXD5IRhel5453TJ2KEm1qycEVYLEtPd6ObyY
u/qJlVmJqaCbnER/SMXHfdkdunkt+up/c4UdHiSDUpGTIA/RNA1j/W5+nLGuFtmi
sCqY+RiwY6LmuI4Z6C/EdrVgP9oFvIa/WIa1pUPfmzr3c2Jg+kZYeGnIeGMLo/zB
irWMkDkNthOoM85fMycS1LBnds2APOyO3TyG+YU45o/uIQY5ZoDe/c3b7se6YiIl
ZhouOsnKS2aDTOA9EVeGQ9ye3z9xYQBjnwjq9iC2URgeF1BKEV77W/a5ResBK29h
YVX29dqrtSaty0zYX1EbK1EVxBAviEuhU08IhI+h2HQ/cIsiN/rgR5GVOa2KdAKn
Amu/j04vGUcFzyvU2NGTDk5QVIIJILvA4gF9DFXcBgjS9IGoasRRj4HpFJThF3G2
nH63qWIJqHp8VURdUBej3PoMelGwUnNEtilEO8xOFnbkuNX0Mepa6/0fQ6KybDqt
NhX3vjY51qhrMPBuvGx78uD2/tlw99qWBa2HEbLRTWFSFJ3UBuVJyDxV8uir/ddI
3oJq7gA5EEl+6CdZu3f0HgzxOitf7zd0CAY9NueQ0gJVw1uFIV7mjWygwU1xnnFJ
QOnxdhFFj7a/6ap+a/LeXQslTsPH08D3P04tGalmpExc0vUIJrIxzUcPOv0LdnIz
C7OVnPsjDgW7HIj/8VoK2GcEDfFwR1uFsskSbxFs4/GqkhwmQ1AVll8ttIBLTUGH
OmZbuNDLgCFq2QnY62FPQOJha6ruU+a+qw0KF1HImdj6EQ6P2jpyAipGjFnROBRm
xtF9ek3XYRvGxMVZP8noMesDyLP+gwJ/AKY6px3IH/orZ7wF+9s6SJaNAK4MdyzT
EDoyem/rcwm0ExVboL9tizvCW5FGDmKXjWI/sEIdqhKnXjlAWMo1pRCP5lDC48G8
H9UuCnTOt7YvqA81trJEzbHNkj1MT9E/L0j/1GkZqZ6gtW1RK68xnBcDfXow1rWg
f+uhEz2JyzbAfcrV5StHyBlAl/fudcSqwqYFuYGwOpeAbV0hLD1Ua2PMQSieCoxn
qnZT2nwjizMu0+/E2sMPUSgoPI9JX+z2i8W/1o6bTmoqIgMV5EVzrChyIz1zXE8W
oGifYA0uYX9k69WozVU9kGT8b1/USrREuNHAi1doJ58ip67qtyI/edTyAi1BaDs2
Ehwip2DLtjx0gJvXgtFdqU2+0W42YZMoSHyj4ZILdO9JQFcT+rHVZYssQrZzGcu7
VbPjONkW/nnBZkn0TpcIYGZQMDO5pavdM0H9nUSrBN7iyL57rL4GFLYW/U2PRo50
a5reM0jLshVHkIhP1akskDPEhFZO89QykrXnzINzitxa+PG2jGw3S0flCxyMUw65
t7dymB7gTVIwsjB3W/ul+QEdnA+qR/n8lCapy78tI0/q2DzPjyhSX2oNQH53QQkq
w06Fheog0lahbBNasntfFRuoONVuKrVumrhmpDHbT1BbNci3QSLgrXVuSa3R7W3y
Z9zcU5VFNfeltmuqJW6D/MlrWyIfUOfBP3Ljv3gqaJO2/AcKvJFzQCfYbVi+4uzl
qv9Lu+mDtn6Jj0YH63RCvTUH7+v1jzemf+52DPP21uH8rZFhGMStAr9EVIFSMtMY
QxHpJ1q3KupALiEQuXmq5Gm/TU/9eDFsrw/FTDjLske4vso9uRW3OLCVnpBVmPgV
wo+hSR4lq+kcwUORW7V/sErwCU+UB2W/wQ48wPyHwBD/D5reeTXxBx5MaviVbKpF
aERZVHYifXbcHgvhny7JMSW+eKVFvcwSyf5a2jx5O7212yTmK0VP2pHvrxjn6I3w
Od+Kr2CcbQGLOONjmgZtXqmPQetsV5/MK1tT+6oYJT9kJUDOfsMbK6aCoWNFYgo5
/AcqXet/jL3AtutCnhdBBlwQtyoKbQHB7OMY8QNRpWvEzUTG8WWzFESZ9OloforY
Cz1sng0U65lLwYgZMsSc3vE+Lf4vTaCBGJ4VimQ5TZQSyK8p9lN+iQlcq8d0VEXT
6j0Hijs4jIk1xfYN9CML8gj5HGljRxFZNzXkVh/srOT68JuND1NQW9SFh3ywGMaK
vBy3vLqQ6yVCOcLHZFQ6uUjv2RxAeTzSWtIsDO/vIXGba/YlUNkbaEPrK8qDHj/J
H+GGbq7t9kfo3iYWf2v7xeVy+Yz7ZckpwQ7ARRcyYf2+4KIa1miTFFJOndy+11Ep
fcNoGvwU3K624Aa1KV1LkmkvC7xi+z95JHzezEpKRXn3e+oBshLABUF31jDNTS27
fnNSxwKx69Y2iozpJ9lq3SIty4XRCVryrgqWK9g+xbLl+AReeKzouSMWAchD/xGY
Si+UDEx59hktbhWMi0iwv3Ug6mgau7mcZTWwFCxBJ3QDq+/3y2t+Dx1t/rB0Ds+r
Tm8pMcC8iTQCl5Rg3CMjyYYjtdPVT1VczP+GarKq9vpz+He6AMXJGXvE/mHYeyI+
l1b74fKc5JDQKNzRRvws4+bPO+SRpX3wKERu5hlUGQbdnro4vK07mMBiosJIyWWL
3yu8Gprs5GENhdrxKXytkl6wiyOzubT8qdT3DTy3VTDeKmyRe3zTjTZuagzd07kB
ADwbjd32oQQ/Q6CgFy5Jxba5Zq6sKhwmZT2V/cSgLryoIx6DeB62jvVfTa1dc8SN
TUOjDEwbL4y8A3oQiKevLWK6WugYrejMDn9qFjeZ/KZz3NLiYFZ1Iwck9CULSa3D
8JAH2vODmq1sIGAqyzv/h3bihJ02FoPZjT5QId18n3L/87bQO8OCjcUfZMZemRAu
hQfNIMMWvBYgdvow0Lnbbkg9DRoiZYbcCm1q0aLc9WG+/c+ZHYq3m9lXuHI7lorW
A7Yk8BOnfVqUnRd5gDkCdfc8cweTwfOgDWo672i9/RFjsB9BlPnSHy7x3rmFbPsg
/VhUResVdXo1SIyfDly4SvwBbD9RRDfnDrjSf5pFjZeNGk9sbcM5ojC3aYNhmb54
O1u8SVHzlpRsZnzFi9UZ7cUiT8fD+ba6VS+avDBHOpUBbPurWXVW7R5KEST3J+BY
SorTZmOeowLaBFMqrfC+yWO2gcJHOJZ+YcBA6VGuDbHWKyeg4Spt/ACYG4Dt6P9c
wJJ09+Mw8Eb5tNJfhmTa3+y8kyDwlmPDvHfV0l9551B+97tBiEzwxSGWepk84+CQ
Y7lDFNvKSEciIsqc3mU8g2xKNAreM7kOSC9oYJxt2gqKFku6Ak5n3lmC1YjLE4KY
JIHaekgLYsJ2AvYf1QTyQinDk6TPTpyd7r3TWioh/cb4QKAAV7NH1Q85ujdr6ahB
mi5f78DN98AsolblL4liG92tjUOXJ0hJZ/1ZlUEHid+xm8rUggFyTvCuLu7vFCaI
KMvmgsZr9eHJ5upY9hhOiOSErnZNQ/kiEt31WM7BbU6yp3sLGfu9WAFyF+IIWQHH
cGZKrPDrX1Bzr5fGiRAbKUsgmSZ8KZtAie5Y3Dvkzu1l84gnjNUPO1cq6a/moYWm
xv6r7CF4c4jiDjbxaM9EELYr6phfE4nJOmUtW8ZCnr3fllPBowsF/52ukQ8cdWh8
B4FqPyYoQfKvytTACa6y7+JTMn0z/LaGNjqu+Z3AYeSs4by8OxXtERywNw5a64wA
jqf9B08LertDD1xFm4KU7lgT0Qw7597UWkOrcG2YR7qAnIiKnR3J3jNH+Pa7jFr7
8/E4qCBxVxaDyN4RfzOZv1cWwbaAfhndQC/wiAZ0OIAqRBcOUuN8l0y/iYActQrR
8hFXUlm0xwu6beLlOft9PFKNn8qlsbnZUyFVGIO7/ovL2/qYw2ad1BfA09nYqpdJ
2g5pSZVJrBKCWTz3Y0Ykaoyup3nog46k1JqDcg8aQchEYBeuakrbz1FfqJjN1iQZ
AoqtAORi8gu/nWT/C1AB+Kxrlguda3FrV7XYb5iO/dCn89DM0JtIlra3BljUmfGi
n3N+6BCXUl3+g4uVj7B+yeASRdyNMiBUy2EvMBaapHxdtGULIND6EvbzxsmkAvcD
TbQmjoJxKey2OsRjnQfeY1nGc1HGrwM7gM3wbtGnZ9iR0QmjeazvflsZ9Ow8yLij
nL363j6VEyHJONvqNDNcEcytPW02amkZV3dbmCC+InDkCbI1YX8RVKa1R0cnpjgB
7f476z4Dg+hxacMUjH9lpNF73fVC1HOeOfrMJrB8k82hq6fCJkaNHxw15eAg0KeU
bYGrJNjzzqu0v6MmvOmHOH/wvpmX7MfpgcxgKSB1UYKlV7ECYVhxoIZfqGhOplYY
x35PZRSNajiDQ+l0hPnqHZFk74JsqwRqskIQe4UaLbaF1my72RmEpfXwC7o1qmfj
kqNQyrIEGWXg1fqOQ90oPBoR/rXeueuwieriJfM9E/Ky8kQ2/WeoBJjiVCW/cthG
dCjX0v141H5V/tvI3OWN8zC+mABiGYfWxh4g3SNwyN4IoOf41gOGQncFvyFfE8pD
+9BkiWKFc1vyFK9qh0EKeH5rNzB0JX+8WXTQqbEdPHKSaa4xeltZkASZVDxRdfFI
8+u9D8//R1ZKHbd6K/cc3diFjS/fhSTya3TO0tdZzZHLbHWRcRMp5yk4XBVM/nT1
HJqYX2DmVYCchr5nyj67n3jjE4cy/gBpE/3aAZ6EbEFGRPdaV0gY1mbSQi/B7JKr
DdYw8rt9/H62E81IgwVlxy7upUQ6zuBEzZyl70xfOz5FcJ/0aojRLD7w2jtcxHFw
1xOMmT7FnVRvYZ5uSJ9ZDiboabhT+vzAvUwnDoS1YnBHCDM9yduKfDRhcPa7bo1N
eJSp927PcM96XGK04z5iY3kvlHCnTKxP3RiMVYdzOZ4lk2U/HuWrci6xU+PSF+1B
fXNHWAK7rxGcpDyX65dvybUYP7k77wWsfrDsejUh3h3drRIWRZLLQy0FaeLsxlWL
TZUhomNV/qwax6LHzhzMI+Q9IsOFsFLk5/6hZ7jGShGJKdxAi5Hy0qsrup0K7FfD
q08SJJJ3JA7PNCi3lXIo7TOa/BRcyfJJeIkJ91k4wwvxN468cgccN32/k6DvfyEm
CTh2jDEkn5RDMrHDT0vU80THhf2NeWcwKR9VzPMZwLc4XGzxXtk97u+mxpGWuUCf
cBbQrvqg4Xjnhjc1j6zxgjr5S5vE+7b5StMouroxsP9iJkTSikNgrJCq+jJzwNfi
v/ZmQpf52TuNzl2jiJrNLhQ/MUFKvGpP38V+CmAFNuE4gKzoabaUy+959KQAzZ6+
4sI+dpEdnMefbhbaAYSOeeHl5H9WPJTxuWAGMOrdds8fj79Dns4UedxLXVZeFguh
n7tWXoigL4DZZ+lIcp7orepORh4kOKYbopF+pAHuOAYSo/2vq5d/PTaUIgqhkoRS
eTX/f2JWwAyZzJFBEGyk4jwKE6MFwHUWJ+0O63/y+AjFkAbkrAILjJS7uQQiwj8K
dWzDtRekVneeLSCUKiMc+cPfC2PkSTCAu5Z9EoTB8+4S5IkMte+l32H1sKbsECV4
/Ac6MxDsc362azFTHRBgN8PyVy2YtLSAzIy0a/j84DfIdgDdLZvT7En+eW2d1F1+
qkTE7ARJvwtkdbQ/R2n6zBsEj7fYaXKNPAQotAqRkYwCfg4+4mzfzoulcZY0oyiX
dOdIqG2iwXfp5SSVSkU2XL3xhxzeSTkcpfizNLRuriKD1WDBZx5I/4jdgtDDbLrt
pKDHPMmASEGdX752sjBc/g+v1FUTpUZpT2eKh8TfDI0mPe4/il+nCkoXxKjT+VXv
VFksu07tNeA+mG98vVgatagfFjb5vplgh+NNnMYIsFjzcbgm0C/o5t7VxuHy9mrC
NSRdhXxIhGqrLNCkpOZejYb1RRTKFUiGyNmLAzTfv79Bo9+Nzhq31Ek/VSCUCyqq
PhT7rb842wy6qXH/5KG81fStng/FYCqSbT/k+ycIkdTiOQRdlDeZZmHo5xd8e2oz
AqQ/pyzkMXTNLIrQxqMZmnwpSXkeid3TcjhbdaCKl6kNDacc4oohLfP82WGqzEcQ
ZMKeE6KXGtMx9hL29Jx1YR5ig+XCtBcu9D42g+9w6NCE/HCtNgeBsq8KldYEDVZt
Fz4/roeN27VjSU/d1Ma7sYOXb8x39tHAPet5jebPxWa8QjKYE/SMiUOngAfOE2DT
6huki8Uz45GdQv5veBhtk46Gy26yVArDnALbGeu3AuYxq3rP+9jIsf+SYutEo5+F
kGMn8+4Yh13C7ZVFD+SmqUGgydR296ev3zWYLQn8j81y2ZwdrV9n9ngs0uCf0yBT
yWjxWcE+OX/CY6Scp8lH+OaR71wSXucPzeZwSqLH54jhrdcqfk3S6ARHrhD9MB+8
T7yxcBecVsK0yBraH4y3rbgq/DrEIpVI+ZMJLB2iRINj7MrG6aLdBwGEHqZX0Il2
lxE42oLdqLrrj5H/6js9JJVP9oJI3ujOb7VtuENxu1HKNNDE05lw8GqdhFk6HagI
y6dM/QAfq0U5hS/Q4iHJlNfZAElRvJk7d+Ji3f6WItG5NbJWYRH0Bwcf197vMS5E
5YCP+v8wX3iPYxS4eLA+cvoOcvJz8XuQKbtz4GCTRvope1552ELGGNONfBdXF8zn
UpijRKQVMzHsbQow2ewNmS+w2jfKCNTqMo1ys9JkikFotHjbDXUbxK8HuB+E/dFx
r79zlMgmdASi4gG7saiThAoFHHPK/NvJygi81D2D1u0ot+E/Wh5CnMx/1Q8uUde0
+WWw3hl9RdUIMq+61ydUVludlQHHmh43jDoeAn53YwZQC9ebfCK5NOpGSA5NelHP
srjUhYPV4C8dKaGiXSXIYsYyV4iF+LXg0QjXGeq8cgIeeIlfmmFX1PEIHizXJHFe
Ida9NwkbhGSXnbsCGbzpc8TLB7h4in3NAttVTa97uehimVFy8lEwWkQPW7H/ebfR
99kz9pE0EYD3xa/mahXV5O441TlUzCRN1fRT0C9VnZpG8gWJhh/zlpkwxLTEUrRo
v7yHQzqBqGEeJy9ET3E1lFZylL11PEhoyIl4kcc6JL5JryIEBD6hU+HkV/NdhcYy
F9BmciPbuVRwYxOA/ZRNOdcEbnD3uV55qZ8IMpgc6I5+C1VtAU0eZ/sroKIH+Ub3
MYqn5qaf55PGILQUOyRwHQ/YqA9TDEixZHHImN0r2V7d1M6IYmyIfalwU8aELcOU
b/KAoBEMbcJgxWVMF5ANRxExETbTy6NOBIm0wZNp46Sda6kwZNOJgV0b96ec7L4K
yttraTosfejU9gYIQlGghw1aeBK8aGtEOmdMDWRjQxcDBDkiwL4MO/N5KPxQvKvg
CT201lmfNmECbA3ObYw0527SqTIxFID3qdoeTZYUA9HcLf8gYkXGVPvw0uffbqcf
LzLeQPAf030+66XQ4WqNbXvdZU5M3lf9/nERqnJP9jPjAOOgVtVfRXH4rLQAs81O
nfrwKZ0JnVvVH7FrH9Yu3IvAFNrNbWOJPmjyrWqtbZUvbARH1S2ilTdmr5JoeE+k
CeHExMbQzm63TqdORfHynYWjAVp6FWgpIxeTzO7ytzWw1zs6gg4ZMfmnY2nFCOlT
U01UAdB0j5sXQncXbdJ7mP8sziQAwozlEE/tPoE9HQ5/JE9RaC8JS0u+3aGKBRBN
DmzKEGUG0L3w9dycRbfwmmu6+FAZO7xPnqcHgQqmJZBlRKFDZ7/k/R7xJCjsK6rh
/tyeyzfX1UtfJ8s7NosReU2X/2UYNI7+/bspEGyTPzH60QDPGCemCuatdE/GE3OB
L4iY2VK+fV0IckKbbml9sGbpoUazoliL8eEyWIb94oZB+vOP+zThpT8NzP3S67tb
t75Q82GlLSUYB1WWg8+EPztsBdr8cckrkP/3gm/TO35PM6KqD9KQg34fkwUSMFhx
hTik6SStHL4mgQx/VqYOvyFZo/2lhBZTKddnFl3DA/oDLH8whzzLiuJQlBXE5HBT
JNmWtEkAyBImWYBG0Jq2z/A6Ma2NH27+JNdUoH0OeK2QEV4/qE2tndNGpt0e/pgC
s0LIUdfFVsWyS3VHIWGqH00b3d2524Y7t2vnRcT4fYvgZjVLkRQ7C0rn/yW0r4pa
e6xir1x3/5M4ejq524tfjNcwZR85/5zezPvrMras12FU7QswBH670Q/NiYuaqYbx
7pyN44zcFpL2WEqabaqZkEDCIQemkm3bXWkVzjnMrPDKcYEAghi7+196dJLGItZO
uBwx0Mf1+g6FqBqNKd5ZJZZHFTEzQHKVA8PzBXXhPBS4oFdk4PUj2dQLaMz/KfVC
Y/IXU5vR54CJfQt/SSeMjHoV3V3tMA2HI+HnNyOePQmWZMS7/3Ksaq3ThdmXGBgr
eFSY0W+sEDPgrJGemWZWXEFn4hZvOVqGc0hFaF7KoeqbCYBx4e5T1Oem/2Rm2KjO
HNEW3WaVfw8u/8LoEmETpTgIB/NA5/YxvcvC74OCkk+b4WpqTqbozhTl9cKH9Eio
32S62WPxefKST1MiLoZ5T/fQS8Ngh94SzsfHanZh/WatNKbDbDVgvIxZNqc7QR4L
CkWQcI9JUn61IvXIEewWerwDlwbLESEAq8hAMcmULD/NL9mEf68BIh+PCayKyzQd
k26YBgWEGt6DusSEXsReliab69fW5z1ISgmLeMVk9vm3QxzpLjULQ5tzdQ0Q0522
djQAjXTJW7iD1EeSICWIgNsya2reW/MdncYbp4lD+pNLrF4opZRJlPg26VYjJF8O
YyKFQB3/D0x2aQizKRUBHYw5ghFbAndYHvz5o7pqyKo8xZ0NQkecNH6Y5sRk2YsZ
ujP1V6sOPe8vKS+JGpSrSQxx37DhbAdgUKAHheh0gkHwF4MtAAZ2W8sj972RH7iv
Z6cBDZJPumeSG5ers+NvgreLE23YTbf7egqvPKKe7r7mytTmacEPP2i3re3PENlX
r94yS07DwDr1em/ysoyrp+qOruY2xPkteCndkDWDll93njl+GFSodTE1kXtX6XWe
OnRzWavHIWJdjkZ7yiu6M75I6meChtLMgg74ihqwUvJiIrxToAplcDiWlQdDHkTJ
vxNYHUr0gJ20oFZvFLue7UyLPue/5fOw/dD0BpsWdS5k+Zb6qB0RliRtMviOZzcG
05Q5KQgU4K2ywYJJQU0LyIaRvA8oTngeDEPt7y5nbTnEAQ9rNjKlR/TDiWDNdlqE
fi4HteHIfVUQhWkFHd+Nvi9AQgTRNn5IZusuwhDvzRWCVWg2nvvgD9ZuhG/LdX/A
kUGS7mfd9iIevXosWR/zz7w2nqw2DPoXDVO6jHf/LbWkAR4TuC85HmfN7oI6b3c+
FJqNmWGk1m+8IdggWozGf740C3/MJYcn+xLtLmHzanoeuMgxCN5BCGs2rs4ZVETI
qKSNHYOktex+8zuJUzKPrEXij7aeaWpeT1DqA3IDjkktVuchnCfs+xMuy4yJHJVb
0sJTJH7uAcPFlNm1KHfquvVp1XKCTtAyTP4P9LcMuCIiLgHVlUL4CWmuzJ2AV+nk
gSPc8TaS6vm2bzEfX1Px82goVN+6EI5qLgy1G+EdyAo4A+lWaFvedcFpYLHDNzp9
vHcnsPrZh1vVOLbTLcd1Cpw7oJLFdGD3WdMZVIaYwst36vk93/Bv3DRYd9H1JFRW
/O4vSFkqutkLb+ufzEpcpddFVazgKI28PG24TKT2LGs8eDjlXsyWgtnrNtQaTkHU
C4iqkjWw0XgK17uJQLT1ftNrl7Oc1siEpW/2tlDdH950OnvmqhfLWJcYXb4bDh9s
oMFew35v4CHSU1yXm49Yo+SXAe9ehJLNLEB4c23EHCHoSWDxIlMJQxQemSSvUg2w
mGUINmNVlshJk0gsfg7DRz8DmfbdrHtne/c/6tdAnaO7xMN+AI6DdomO3RCtguoB
hddz+ciB4QJCPJVEu6xf/H6XZQMs33zT8aoXKpJm+rvI1m2pz3REKiKEji6aiOZ9
NbHdEwFvKfRWab83PyvkKd+ClvQqlB/27SMKkrTQ3kmIubBFF+JQBlTmDhjq1r7D
AQrAbCRx6lJrqKDwIbGpNvXgZiDBYR1rl/hSf3RKsViCtRSJjJza8hPm/I3UFQBH
OopLknbmARBwqPZ1ab6o9nI++5A6K1Zj93W+JS115s6v1NQK1e8zeNK6OIKQmXeL
HJXehEqwd7u1cwlreWalhquA9Nof4soegMGmOVmbcYJKTSaeMg4CMaT5sglozb/J
n2sAJoD1n+J5qIHa4PaQ3BNINl/4O3Q1GbpXhF5D7z6GHcWW5j8IUVRG87GyhaPX
l28XIiK8YsNtT+cjkQ8+Ljg3202y87aZp591br/dBKl2GdO1wehvvhb+dwUXkG0w
D+YUm+a3GuOmYNTV6ewPYdY8N3JAfqwVE1yk4jWyrU5ASJNjhTn96ZWF1zP7oDci
wKGswO5tYO/+vpL7UpgZkrtt/5sWD2bKhCKe7ay4WUxpZ2uYjtX5IW1JQ9ufRwLx
30gCiI5ODRpJVt7SE8/uLa2bt4nSXeoqCPypehn3ZbPTHbzekY0nRh6qfdECRKLC
5oeXSApRFYlaogixY9awUwx3p/f92LYlrWSDQlwNicIdvccD9jOnyl3Cc9plNSDF
oIK4F1A/kh6WGDqH5/nTLfTrhlvXXaIS63WAf3T543DT6Am/rzq437aHLgV84TNS
pZD/AEZkqNQ89s+C8OoT4vUl31t93QnzKBa8Rsu0THjW0L5xj7l3lYkreo4rRYk9
8tNJnajJLgt0CRPFo62wpqD9Ot5Yx8mZljH62yb9cytq9M4+90G+RCa8XPSABHcf
jo1AYUWG5oxdHdodcycNwPOF0az9deTwweI+CPzdg9fX838gMfw+oI0chqklts9o
On45k+BYhrCeO2qrlJEshiwMyJvKQ3p4XeFTdNE1ZAvLbyKnnI45fj9Ub9RJ9rmI
eaEmRxUBMaSROAKh4jj3CbafiCnwnOO+RFqnYIIUTrwMPtXrtmr1Z3wSM+JfsmB8
LbKOdGO9frrsRvroqHqnHMYzxmzIf6UPfj5lo2v0V7wZ38NqNNhxZnZfUBqcsKkx
/Q5djUwx18don2Mm4POOL+6gP2ci0K03HE3v7i5GpTZZpLGRMjT2Tbji0WqE9+o7
JRfMFu/7E+vQOjBh/LJZukYWG5hjDAKZyKHhVjIygm4KauxQyzvXOQVH6/0PMXPK
3+6BCUTILHUYlZeCduuGZ6Mod+jP1CD8vOsK9nhlYL2a/fPchgpefTOJVBUm8HBW
IaIT70LvJQHeHzoXgi4dmCBvS64EGmEI3M6FNo5pm9xYITwIfOTrhotV+g/swrEh
X+Xp8Yzu3ki2bI7enW5Po/9GZ3as6NOkvprxQHMIrlBHHEOlzVrsMLB9Wytf2BZK
XkOWlxWeJ44mxocPo+hlZuP2k6VJxG5GAB9leF4UjTMtROmVGZ28v7qx/Po6Xq1z
c5ClDtdigRkq3LWNUvyvxw6t0AXw9JeDsIAsbETPb1hMBmRrM9ravoBNgAt581d8
mFS0VqAFREFsEwLSwKkz1SjRZWV2Mq0fKrXGaHwLuVBx0XCOwNH77bxL5597V054
cqjBi3IIrnUsWNfNuCdihOtsceZOMdPN2cI49/206DbC+75sIXjgQc9bkdGtHpwT
xWkBTabdn/sU6PiomBspEZIQtNEyd1u9f6ZDB7NPU9O4B6Er0YAcImPm/mhuwtoS
F88saYIwj0JgvPy8788HYk60AOy7CfHZHYf4x5Hsmx/ifaLxbf/zk35fJV2xe0uw
5jQur2asUZwOgw4p2ceipqaiAPifATZ5ojVoIbrOaVJ/Z76F0YhTXB+gFV0H1dTu
HeQNDWSiroyvB4AEMq1PUVTKaYiLvwudi3SajQ5O9UQee4o5yTlWUe9CuKzd5ayk
OFlsLa2PLAOFVLG+qFsJhIQZEI64YFBzEFjD2CIVyO9syAtAqMWFQnvwZU+K8VE6
NxhRXqnGpK1T+cPrWxMBMlkw3S6xmnmKqVMcpRIfwxPYUUWSwe4SfyxRJ+DsKWyS
bdlMGPRTgaq7sJCxFcFPXDhaf0olf327mD1nqShmDVOA8kMFBIB8RMScbeHHoAku
B1vY2Aet71gwOmxJz6AhTfoVp5lRk8JcQBQNgHLOmfkY8VUxT9DxSoTT7Kxau5Qk
pUSsMbZ7OpUzbqhKf6CtummbOvUfsJFgm1qzo9pTLbIuD7xB6fdOpujE9B83ZQLN
7kxdgt0dT+jEtYy7Si0ec81oWHdrBgYoBiG5KJdiqd84fuFfP3fr1c5LlI6PKu1W
H11kcwEXlBScJ7GsU3kWs1n3C8bVoQ4T7ge0YNy9/XCdUK+Y/peQZ+AL4KLq2556
Lhi06J1OElSveCMSsy2mDy7w94n80F+lnZOiQk2sr3DrIxqBuCo0UJ7D/HYsKY+Y
ms7D1DkpzZODS8psZGqWde0vQ445fZ06mPrPMDc2wCk3TFa+16Htmp8Uo0rTpiQ4
GrRQyuPPzw6Y5+Hs0zITNEkUT6FeB1nfcp2Pgy2GLSv00BBVryXUjYWWUmrJmBv2
HcHXUrt89WFKz9Tk0uR8lgRwytgZAgna7Jne22pmLuNn5Um7U2pYn0vIxkuZbHMd
WQaJ8bagoLoefa3Y1uWFJ6Lc49DaiBPR3J3fcoYnMk1p5fpPH3dXx6U0Q4pc2wlr
fwhTi84Pn+iTGgNprwodYBk66vsS1hOeW/9LPBDVk/yKoP6z6Ou3FtJNAPHZAjb6
dIl4mFQvd9sbPcQWbVtTjJeSc0mtszu54So6snhOLm0WIln4/6wwASANnhwj9XsS
Y9gUvGZmaSU2n7vA0oA9NMTci2yZ5itxyyOYc4sFa5qT7EFCis3OUVrXXI2PGI57
5v0AMZu4cL2pDcg5GX7AOjXAsebq1bnWNgx3vm8vWD0K+9j75eIRKh1kV/lmQm6T
/t4Tx/YE4LHBtDA0y+skqkDrGW1Y5MHNpojym3FmZSJ2hRMk2B/YKQN3cXE0nkgr
yn8Vbm4zGu7bnTf6YwHiFQe3F2KvmiQWQbQXftOKBHA9SEu1VXZS5P2DFyoMPIye
VaHVfF0u2m66fLKg0U/AFq02X2pfPDSObgW3/5Un+Dx64VPWyj3HrKFNT8AVAcwX
prGEi482mftzF4UMfc4U+KAMc/0ZmFVDznOQJEMnVScl5As7a4vPB+lMxV9iftMf
CEbALdT1mT4iTeV4LjSetJw1l20/cJcsQWlaEWW/w6vC5yNYmpo/eYLgleFqBkxS
sjQ5Ysyyfh1vgNPYzsmBFxEHY0uetPJVFBanufQpw6tm1CPpO3TanihyCezvUxlu
hGVXF6JPNjKob+m+1m6KNtnKszBdXK5nPfTnmDh63ro9+iNdg9+I/blaNpTbuy2s
qCqK5RCQWCVYFcLLXFlYOSvvGL+898+8fttzI0s5EH11tkta/Rv2V7wF+PK1qrYK
RVaB453KHssbfffs071DhBp0VYGLSCZiA0umWr2ZGyTgSJItbcwacWzcxa7/mWXn
DAcgTrfFcnKcXroIVgkAxhN5YAA46YLYh8hFd53uGhuAdaYFjqkZyYHttq9yuogb
P39yXARZy3k6B1rxnimqL6YYC61v/c0Y42Yq6dVSgLLSyjxBI2fSfGLq+x9rj5pc
fldJ9rVy93n2QDk2TihhC7K/SzOOm+leQs+02zUHXVzegIrt+DOH7VUuyyc64FJW
LqEjvJRJI+zcxqcODXXsBEGhrGi+3e2fo7QDp7yzzgNPnp0SbItWOH76T+imqUCl
QRO90Y7VEgGR1ceW3m1xMFIzX/xki5DmAtnuItcGp/G3FGGqxzOjidTHzmvhTYYy
l/ePzIN9/PGh0VOsxL1ofSd581fJsxTirw2biMnid71IXtaHUX+fs+oAfdYbVCoz
xn690Ru7/0qu8USWVg01Hc9wszp35Rixm7FwqgwGc1hx8DYElh/QIQzrU/iKqnmB
GUyXZScXNvFlP1E5FoOPE7X1y4u3Llra8jqzeQOxFvoj52sHmI4cndIzodVA33L/
NstVRlyqdcTaX3fWk3G4b8ooCUtLI80A7o9YmMCijDdmO0cPZlVwxjTizkeWFXdq
pgNXnNK3yR+J8UFcGGoLrOj01ZLz48AGzuVBXesbd+u0XKqEbds57yqsmYipcAFl
7MM85g5SIzwUbDGeGNw1IMDuyh/803ssLaPdwkpSbByvUmdErT/jRro6cof063gU
b9J6aFDud9XwGRYr4kmdqbtFF8fMwX/fYcU0Iy55pV/579jKjEzDwhFXPvHoVYqi
Ld9hh2dBMzRgR2AF8coBAzBRY6edZT0qDa6t15k3ZuhS0LJrJq1e/vAIV3dzIj/K
YYc7mSH1+/0RbmpNy/wCag6CjlLUnlxcAgNMqVW2evsHPOmPh0AWayvwCAoKAsKy
GXi8Zs78qALvVUf9WB9KnGE0wbkfqssOMRSe0AM2KmL3pvieYkVTBST4OkfRbeGV
7YVmHARFcZcRSvWIiE6v0A5sSKvCUjskSW/lKLXiB/Tq4jCmsZF/ZemfL1dFkpz4
sBCYuQ8652dDKq7zWCg9nm5FapzLVDN4wj5Dz6zijFE70yEeNXcU6ZNzjA2oE4vH
SgKk6CMyZCixnuU1SaN5QR94G3Yp8WSQs2Q4hZaAgbfEae3Krnq4WjVI4cJvEh1I
S7lWK5XlO13ZDCgHF3gcJyVGMwL2NYLsBbm8unZ9O/lFIafsr3Td9c/8KiOee2m5
3FZKeAG7hZBqYpQaZ3yK7vaC3YVcuyIuhm9NtJnM7Oni4T18vJaebDtV6qJHCJQr
aZnxxgl/5SLi99OjWoXNhvv+S1fLQDYzV625r7NdISDLtJ8s5Vap/260idPjuzq1
zw+y9TT3KKeqagGNZM4ONT7jJzlahLAF04rEgm1rv0Y0q9Orj5Nm0OxMsO0UWSlO
nj6n6Q5vZ7H+bS//Xd0LbvSlweEHH4g2jjl6cSMQQYEfG7woEgxr9tluXq/eZNnZ
+IEpZe6/Vo6O2K4+ePPLHAqczc47cPTiGQKtIBNa8HjAv11lRSJL+iV0sAgs+bPr
S/iqKjrimYFt+kM8cyI19neED3u0ISofjCrqXx8p5/Ukp3WvBwrz/LHfEgqfS5LU
U/tg9C0Aqr7zZEF5Cel8Kt50NEPj7kLkQQi+dtgZjAyPAhCq4UKOq5O+ob2ePvBn
05QxSlAezYvl53sy31faU7dxio16uxriR/DVlNLySiIDiPpcnLVGhr7hRMc9pkuK
SP4CReWTwhVXwTYsh58Ekh9hCW2PCZoMOHSVYE54l/tv+Bi25fM3ZKuTXo59KLLb
6xOEcQweylJ0zZUIDDGsTAcw+mBNwpKOwNp8UgJMyp5+C0n9FpE2bGgt6sbqwYWI
t7HqGb5YpAEdobA4nFAqmf76ewt6kvWiAQgfvhb8lLfrOIhTxY/OeZvr0tPpLR0P
JAAQWpB3X+DDkvgBMBOvwBKo3I5+HRLyAOLm5rlH3et9FUdpvtLoqTMIk3jYWALt
ofwg/p+Qy5muye187SwCFjshu/EcniM2ri+vFwPrDRhMdV4c+KlauUGJqpGKE567
0+VgFlxdPD0ls1p5wOzvEZJv1VcgM3X5qdQJjWdTiyFOUCZgNLNoOOq8FW8haTcT
dFcLZIO3r2J8vsTpOTvLjQ/9Q4bMksRGGQ2+XECjrxT1Dfp5unq8J7Blpxf1YY6K
Cc2JBCL0vrz96T1kzIZW7aWOFGerD7h1zICfVofyqEOJj1GLTQ22Iy9ZLZtbLG0T
n/385d1XH4az8nKOOg6Xy/eBEx25q9EpJsk4yNRa/dNrFts2XgiYgPiN/BKG2EUl
Tdx5aXxE4VS/4Bm2UPLMN0xTNv67wJck0BxcVxCBvSHanUywC47ixz2n8KyWWiyf
9T0IavH8XzGyMFLvxZOpbrHqoTvCZsFNqKL2tG6f/jCFmjjkBULz0ezq7sPJ7tZH
B6T2IIqX7EmP9ViOOktdrtLphiGkR1LPjl9VOeqDspvvSpu4FwJ9nHqj/CUMvmYs
JJWztunL//VFt9a/X1Uj/qokLrql8x2iSibMnfI6G4WpTeg8lCDdkbpqW8Oyu7MD
/0tgpN6E/ewCZs46XQelvCPckz8IhXiysxmXBSMdAoME2MRdwUfh6BpMVk7OSrnj
Ygf/203tf1fr48RlUHS11oC77Qx+oaN65VHFfN+NB8/8O3AkxJygWqLr39oa040P
KHrOU8Q0vUZkiqsEQR6O+kbgu3DT51cNnLOV3gXiGf8ys4LHut0Pqhan+o/JGUgx
AfP5/PE5m40VM5xGU99wn8yzjIxKTxCX2hGuLbDiePS9z3H9dL8n9ak9aexLnMkT
Z29UaMU5afbB4BSzqRSQjXa64oNYjv+JfPz0kfTUCIYd1ptfNWrcmORT9YU8MSsD
/U8wqs1w32nvJ9RAhKIGfcWoB7RgZURk7dDB/XOKs0UOqSatCI0f7tu6L0k4Fisu
8LZP20criYsIJC++emWcYqOhWtwBNawrnfVK55OR6MxjeREjcvpfdTsDBgd/7y0W
Vsm2ekXBi/xcULVg89rs03SNYJTgkm0sfbgK6lo0d5MczdLtZPJjAt/jqjQ07V+/
/0olb4Lby4H5heAWpm7f+HI61cI7qjJNagiuW0UHG7Raw7cRCu8tr4l8bz0Pj47n
LskuaEqu7jgMmx8Rfq0HBK8NftHmyZOC5Le/3oqw9eGQePGe7mhJenD61gGsb7Fc
Ys02bDY4A2Nwoxq5KF1DjUxyGHYz5iGdXcSV2HTkEAs7b5YS/aMoY+6tcDBA/qbi
e5mKvS9fOkpC0RcQ1bPH0n49uyUd/JvvjczQQhSMDFeCZOH1ddiqHKycltLKvJD3
vRhawP3B3SSbQknjSi1Bk7bGmbKkg892tJynILyUFraaRkouxYRxlB3fc/V4YU5s
eC2jtqsrEQLAPN/3jDkFAL9xJUtUKnCxCQMj+tNZlfszHjVfDQ06Tsui2Nkzk/95
yz4bG98xlufWnPPJJo8nJbBajqEUNlAkd4yd58Y2clNAXmModh24DIfs9T7zMqLL
Lqv3SFm3Hqr4l6IyivGUKVDl7ywVARHiqq/1WvmQo9wAMPqFb9FN/gR99lZbkH39
uMMYRjcAz5kgkbDzvHGXBZ175qsmSY5JUdjS+Y4OniLZdCde6RB9WrA4eDSzwtdp
FjEDlF0GHPoVF0aPm9EnwMx1lxDDd2bEPQUwfRAW9wDYgx+Zgmawshls7hy25nKP
c60LdR0wYzkdBN+YLf2C1+TWj3PJdmaYE0ASbP6CF8kCNIfFmqbA1Oa7o6qLqWrx
50m0vCELN8JePhmvzHrlbFr8nelW2yaPQdfIQ3VEm8tr86MPOz8+tq1cNWFIgvt8
GcILMc9enZWBqd+ATZ5sRvt2mUSj6xznJhIThuU8apEvRkZwnjoEa8seHz6HYQi1
Yo6TbW82TQeCYvEEGvFGExHsdp/RYEYb7mSXxlS7dQjMN2icfrw+I8rK4xizYSW9
OBuuRD1PtSvC9Dfc9nQyLROznhvUktzuqzcNz1mC6Cggkuk3kUJw+MfTp8vt5yWi
cywiszfA0VulnQPiEBAKgrSX1E7aag+DMwUzFDNZ0jg03X3Qv6zlMaF4n9aE3aYO
MOCdkP01O8xQn0zDLCFjUfwagDCbEsOnILnS5XyKqY1pul+RE4nIjpuHgXgFamQ/
po/QLcSkEFeD15ld0RhOxlBbraw8HSYlNBKdXDa9uI7DrXQgX6YRShIFMdopCjYW
mms1uB11hZ0oXQlNorZ9eFWC1gU0lTYp+3ASebVu+AUR1kVBTZKvvJEyTG/Tyemw
im5QwrvkVTyH3f63pbV7FNfXJSZjl+EbfdZDYhE9D/pAFmnQxK4kjFWkBiQHoA+1
ZEHNca6mhu/ylIwtmw9nVZ2cOzXEYL/qY0L0sQ60i+1ZJLcJy6eqR7zeXsAotok4
e8X8ozfNoFfr5bkqMagnRhx77FUKmwTxhqpxxYOwT5L1h8FESIQk3a3j5CAR19GK
XWZ3b9MDx8Qblf+f6X5lMBrnJVhdxi6fsJXj1TxPl6yrmrEzBstmnhTXLnGaJUI3
fqGkZWOiQpwNydV1ztdWJaIE/g93OFggq/XeepSscej1pHUuF3pz447zKfKHC0Vb
R1hvFhdolDlbBXj2KQDYi2kp4FIaqkreMKCJQ7kqT2adZaaWrYNA4MV5jduEiSEY
iFS3NOH6bMxDlmxnrY9qPVU5cV87CkFhLtWnwmvjEc39IXU8HlSCpvW72mghG5XE
3Cky8ApbloyJDAD7+yT/TlCBOPq2jJLIL2MxJXJxGsgK0Aa1nTbXUWurcrjA/AcM
efhatmeoh2541wQSKmFVZGevnAKZdn61u7HJCgp1jHupYArzG31dxpR3Zj1yQ3rN
hPAYRdgSzAhdBOLn5a1Y0oE+zkB8lxOdhRXT4sWErswu0DNVm/8lUZfazPUpelXj
pKP7ZubnQG+HSxUwtlzNkHAKU5/B7HszJ7k5hgsObnZN9EDMgIJpvXtCEI8XJg3T
h4dIoPw9P2JCV8Zude771tASNeOSd4kxdODXYWw/gSr39Tv7D8OBcIzxWd90tQr4
f/FgmnUEUQl3R4MfXv4jIPfQMZxc75yPNvtNqqQw9S6P/JB/bqAz3f+LIUKrrzLs
W74rs3qJaefDAcfhFXs0jofY9N3/97LRp1TLMGzI9hh22of9OYkn9Gtv00H/6gan
8bcCO7sK3+eEyOReQsz0thY4UVM2bJYSASKgsHmLt+pINt0nSo+eRzo4osL0ag9l
h96ptJRicjj7HJ17fWKVIvy5eseeew4Dya11STtBT6OGnpv/vEfaLkyQSRCml2Wl
VPLOruXv9ntwdfKJtmtXW7QCkOMLBQnp15ukaXXaedk885krpWXygBP8cyMvIJLb
PRusi/NsHG5Ip11sHjMMhgAovT8ARPeA8rRT2FAyj/5sAzVoI0oVZlY/tYvOP3GJ
fBRXjqaODFFy+QFZVDnkcxTTWSWFBItnT4Q1ktkVToklohBdBCTK3r8ub2/9vjwg
hQLNm2RhWxtd4QzKtlin2UYOydDF06YxsowJP8LhvUWWQirUH9M9MnmnfVX4Y0ff
H5Vf3qFCiXIY708vZnQjeWdCv2sjgXLvJhOYElx7+CbhGxuJsnxAVXiNzH+mzUVA
zZM0DaMx0YUY11mWA6/LmQpXnwGl5gwY+93Fw2V8rscHDabZzEFDuMFXxaElhO1i
iAbN5MPir75QVEUNeVn3G63+RuSJ/NY3AUeU327SzamXxomzhcBipzDwrj9Z2OFi
vNV5E6d6dvfF/0mB8Oplv0CkSQ6NcGovn/Lqah1JDOcXsY9e3o2c9HUKrkiMvuES
3aKH2pVrXsa96ig3leZ9NgjWKzjGX30PTXROkO/Ba8IBdEiu3fed/kQzjnHecBb6
fTE/yS5y72gdkxBQmv1aZKd+1tSOYuCUfeT5vpoHLEvBmFf+U2KqUlmVhRdNLeSC
Ygk7djKCsFgrIcfa/DRe29Wl51Dd3OukemeIVGfEHXi84tjUPFneyIRXSCepi5F4
p9qFcYcohfuKUGXfPv7VnQpHSEaN8P66rviKa/IW3w2CB/SeVx0UPBhd014BPZUB
bZQV+tQs6ycKAhOTdIpwLWrcT6i2VBhiz6zG1ag0PQ1whZITH32yMZ0D57PpkGUk
ccLpR5dY1+Ym+wHzbN+Dx9jFA4dkk5hg2ZuSLNpexidvwVfe27mfI2Wz6vjIAgwP
+RCFSZCBSXJa4POkiF1mxEm76DeURjWSYTZyYgaCG2ALJEsUJhwHbqODXoygpkPx
51GSH7SLds3FZQ19Buotd6ojiQgiqieu1x5YW9EPGJEHB4JffQoQUMkgoVJDHmt5
4RtkA9lzZ7HHPodST/4ktrr2nFxr2kQ3YoOcaDNRFx2ZXmnI1CbyW8oYtEUcKl4x
BXGo4jV+ZAtluuJ9lxmCj2zPrZNge1zXh/lV8L/pVtdFt8Uu949ZpbaZ8AFcmKzh
ewsEHs3FRewtXoSNWqitReKwdVekW6olEAxMVqyE1JIoIgBW9NVEBTCrP3/p30i8
q24WY2BKQCXVv1KvXagaPp3FiU84j99paUjuU9kgkVjLwD8Cla79VtozQqzOgYU8
eM0cBLCUJSz2vI0wZ04o0aIEr7FE3aIzesiTyvUJyTuWKL4y4xjBtvj5N08u/LJZ
GTVeMlfVWubUb75Ez5GITEPctw4KdvPwrI6tiBb1w1tg1tlCAFvA8AZJjnSGj1nb
KEZOtGQwmtPMxL7YL2FNfl4tFLSbji0ECan908unSFmiY97twaY3X8sqlucnjnMM
tpydaLSylN5YUV6R/GIOXz81R5P7hiBfiCRr6UYNEji6zC+RKRt3GSQfzwCyiLRN
rkiW/P6ilkQ9UmhtJ1c6PMDlLMlT42Ak5k7e4EsnXAfFeDraxMU/Bv22GQyB85Pp
m9xHCMoXWGLBUU/WOKOxcQhzkAhotLrwmSsl3720asru7++NO6eQPPGPe4OugeJI
v2DSvdEgl174kf4bS/Lv7hUrA/OCvZ0C7xIAUOVtipVekzPN9/U/IPvvroLIUlhg
yzIG3vo6dO74ah/igpdr4eylRg2TpVuJ6/cb03VArG46FKnrYgAeZx4ZLY4YFkrG
1B/ID4GE8xR+4kf2TouUAMDyB0gHkDu4RF4fMJY3H5c6mPcqmRcVP0UIH3nTpJYl
UI20Td412rRaJEAs3GpIyg6nzhHaROuyZ3b3cj3P+asGf+/TuQsNJMtuu9U6Jw8R
hxQIaVgGecTvl1LnE0GEYCRBAmm9jTSbtapQqoXahZ7JMJCsKRBCEtZ0S3kyf07o
cPf03MutKVUhdg9DHrBBfVaJO+Zu7hMk3+UYPybMbeS7s+DMYfNnb883hzkQV8Zh
BE5/lDrsXMhts6TqL9yFVT8NCpdj+8HPmr8lqEKgk4U26dAzVYlYKeDXOi34hOPm
nWXdz3oors3c9Vc7qUsp+61wMxgmtHjieutvnaUzt1PeuwEQekrft2ggY+3hFkaW
01CuKspD6nSLuQ8hujrBIcyIvW7LMUHMhmp6aFVc7eE3sh/WJ2SNRvZLDYwfY9zv
Dm0K6GR6SVPsi1K502lYUhRKflTGBEcXSHnZj37+lvowy8QgTdLX6KmlseOZTFVO
Ksu8crT30MVOixOZJzFMWxLz3hvLEouExk9C57kSZOHcG48v4CZIjvUy+zrrVHE+
CTwohnRsZD5busf7QmEwE7bK4/uHHJcAETBR0SUkWjs/cwJZ0rjPyFqS90tSqC6G
NvM6z7CP1GbBJUyRBKTsvb22Lwr73wK6lFml5gJUSXKtLx0+lZQRIcMheNhAmsBT
NvLp4YhlihVquchvY3OxECm3iJjwJ5djtTAhZN9nGGh6ckLDCkFyk2l8m96kIbUL
2CmEClkFyNCbevB1vRRLJYMwCHizmtaNXPH/h+wFHoxgbBO0K+duuX40HAKsm4IG
O2HGgwfKdkz+l0S9gWJDmw6t4Ys7MsDL0akO9hB1T6MTsG/gSYmFM30lQs3zBdYf
3TBL9iyQ9II73TKGbbfISNQXDomCtqkEtcpXMWIa9cC5HlHxO5bPIUAn61PHaMsE
i0epGno7QkKuBpdRUoQ1kp7dBMjIDNXh9UnK5Yf6G3xL2rN2415h5lIVoR/hBP7q
96JidpyGuvFoULGbVl5NSAn0j7+UqbD4GtXY5TvCuv5p0bMvSO9b6kgZeyDk3/iz
QZOhRyXlaYWJdEXpZ2NIJ9TBjq9f0xYgeiR490iUdo1L0U/2VrKqdQ+cuJdunF3e
U551Nir1DTQpXV0QL8sD0MgK8YS5PAWnYQqe7v9R3RuUpjD3TOz8UPEAiWBw9BHG
jjeBr+8CeFKTg0Of/eYh78rqvDX2QRURvK1whtaiBmuncaJ+AxJkNPD7a080gZ44
qGYGBd8NrVuXYbSnI8rRB6Xmp46Qxt5rvMcXLR5NOdnnLcsXWtcIat07wq6xxcDU
toUv/ccwUt2UG7VmgmXiG+3E405Kz7etjSHkU/CYL/DujcIgG/GW4htL42cw7mVW
A2PwBeJt9XMpWaTOXcFLgUQatDbVj8CsO6PFZJ35nB7nIt2XNF4hF9DdlX23V9I4
B+859waaKeEsiKnnsscGXeuEZeROKdbDu3l+IQ9bf3WHIEp9bJO0vqV/D5s+FgmQ
PlJCjB7iTjqxkda7CoWXPCIhFbFxOHRNQMIIwlZWXkCSqugnZ+cQFbnQPGHmZAea
uHLXjSfNOiJ8d12vg9vZb6kPjBmmQgd+3pcLe3+ntQUqt9ybWB8h8OxlqfktIJ7c
oeXhlniaG2Hfbq7dhJM93eUHq8nBkVqics3CSIbSu74IiBGSnVe/jMx8QhpQKC8F
WcIyHo254Ann+18N1lLKgz5J0sIHTFkXDmlqPDEiJHqCszqbNccVKR+0bDmrlLe7
DA4/WTLc4Ibrrul6nhfyhtHlcrjsH7G/eUvxNlZuje5uLOmZT2mlatie9LO0dB+p
KfK6ls15GQzUMoJPIrPkjc/85VENTd7CsF6MSRKblLTi4d/nufPJukxBbIyKrhEE
gkH4IcmstJcUj24HsgtKBOQtdDk1yw6XwTrl9PTiJusGJ5/wGsj2Yi8NkncWiEP4
86l5EEKz2lusjuHYL6FnNQVeEsNEG+0zB27OaIWXrQE78/lMEq3P8S499q9TyMh4
4QbLQaFGaXCtqelBeOpKzkKNhd2bLjmemWK6nsAZdbKBR4BvbEWM0pvWT78qAXGj
sNP7172KjhemV1r+8ff5zZ2JcA95iUPvbtifP6zV/wvbxgb9F78mXT0M7CQokmDP
QdHiaZLrHocNw6BKWk7nacclPkUFM0kibJcAagU03pCSGQaaDwLWytgCjdna5tx/
Et49puc7xDIRhu+x4VITLXxodLmtE85yHd+h1M1+SWSrUfhJp1By4x0pPRRFYMWl
51sPQ+dDiK8yxK2eFnISchzZCi8eo2bItjiFpuOoI6TbaxScsbt8bQocmQL0o3l0
ddW7/FViqPkVnSoiFtCLWCmbRGIyNmIoLAKNv0bVIkjPrzIsFrOY7hXaGp+/BJqc
BOFvcl4OCc4WOUBSaqpKuPYh31kWSQ+1+5Lgxs76smMTVCHG5Oxj5UAzIGQJMk1A
`pragma protect end_protected
