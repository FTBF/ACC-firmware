
module clkctrltrest (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
