// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 03:56:44 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SdkPinroSHWonkraj2rWfWjsMGjuLy1UXVFG1C6KPY8v5FsTCtdeEvZUiM64ndRc
4x1pgrPQDug9KvDD01S2u3EvFxMftQHEGnAv5tJ4iHr8UzqSdVMAmEcuDf8BN6jH
PRDyz8nCNiRO3FNDdnavGHIqyEkoEaAO+BaieH7Taw8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 1760)
RgjA5+H3xGioO6GbH4Fy9wUlFOLWEy4aF/TOkJwthWdX7DaPbWePfDAn8Q2STpfv
SP4Zm8usT7JoN91T9I+wqBXCn2MLB0PizfyHS2XaueZCx++FnLj7tNx7zQ0RWvoO
Io3fk7ngjkWabZnBBCqM3qi9faFuhz5cWW8fKvyZzukWCxN81UYws/qpDwJpNrIX
JkoXFuCH6ypeb2WSBXp8MiWonmhUAFSgqNGbBpJXWzuSJDq+JTw/i1cnRURvwwnZ
nL8tOmFGJSlnWTzMwDH2V0xMWamDdCc5uY4DathBNFb3lgA1Jjxv70zPTMd8+Qgm
fo2isnilIXU2o1LzeA4BhSuNEwI6oCXwGDqZ1WThYWddCj4V4TX0gT/zRcsc85ie
9ZSSJ5jw9XPMonzayZhFyjEJ66sy3CLW7UNMa2mfIu2ehTLYF9H4pZJw8DVFKjUf
kjOQ05fICFM7WXYr1+2spddglcBWJN0Fof8LThlGGMmIrqhRHuLEkTstz8rv+0rE
Ld/XSVtu0ebfj/WBl/I73l/2mvTCnjF04CsdYPVfUXBdWIXyRdsU/i+2069frhrb
3ZUQ/+2g3LKNijwFKszh05jxTcOAaKAlkAwVZLCCyKCelRm6hifXGy0SXoWsKYdx
NunU3sJ0wQ4P1w5C/KqyYpEfVQgs2RtFToKMw6sMMViocYp8gp4j55yHnsH6OAEt
aG7cYWdMX3h8uTh79mAVKozIN5HKyvjbIbR2n223FJDwBSGIEGW8auAQGA8Y0jFG
XNOwv3KqIp1vlm0Zujtx12ZL6QQw9jiXLjNnvG9MlIUDuet9YFQklpAD1BWHSQmq
TyiP0vMoOdxDQrATeZMf5pfpLop/+h/rVPWEM2DbktHe3nRPLqaLXR7MmXvq3VeJ
Evi4YgB5701Tmj/mO3LehTh/wdWEw999nI4h+n2O+BQUMt3p2tXrlktxykBT5+H9
zEcgril+zMXL3eiCU8eFVdn70ngoor6o/+j6TfPN2PczDU+q2Tf3KFFXDdfZxIw7
T5qJmv0sK5i6v+AMYy1gkRDlS3dp1jK/6qQ2Jo+t6sGH9EReELZkrID6CFmSsPgy
Hdt8ueqle4VZLsPFfKHzHpBGTUaqHeoEDVZXNUgzQz85QFpsvXxSaU+AzOnEZtJT
8SFw1S03FgS/Wa2l0vyE/uOTcq3Ak44mMjdjKa1DU6zyVX5rQ6Nd5CHcuPso/gZl
5HefSFxQEo8e2szP006VzJ00hrAhH2fpjxHZB0lkrdD10ia79Llkz+zWwQWp+4Im
ezCIo9cbhpv+ozgN7gJCbp4JDBLx8tFBBNCDV5BfZaRf6bBH9kaKXbWSw+OeDPxc
X4OWnej4VUO+qebUmpgRcDDzL69sTs2Uu0Iw09PStef5ttc23HJ4yJewvxNvAwxX
6I00++XmTTojS8/Vvl1+JxprDWYU5eVyHdXeDEzvwFOaVR0EguIK2XOCbHrks3z8
dvdCT2XIs4nfoOX9azGgLq2ZEuWeJAkZmcx+HWWDtypwu7DI+unQwKBbP7RXW6qn
TO3CtfkCJwyRJrAdHB+q8KecyIPi1TrHglByou8UhO0b5f31jFQLJKDl/1VxRoJ+
gI4iWvLSpNAVNWn9ChJ1jjcsJigDTBYBoXhPJmwilG9J8QSCwfWTGj4//jq3hIuE
M1KSi0oz/VlLiKnpDU6ASzqZjITuKhK78V2qmIWBIIDUUnCHaGT05ELc5nhu46oK
bdnt/1ldzOC5Zw6THWqTjPWf0GowEUW9fhWk3RyXuR0tXbj6Ru9IVzMnrFBnyEQp
1+BjPlzCT9kWRuNLQiPaH3DRRs2JiT5pFFGgb8v17QfTJ/dewnt968R174z0L47z
gTkopls+QICMqX1uOAt8p4EVOQJDWODO5k87Xp7beSbikMN3LA2/f/nCLrRCkoEh
H1gvQlS6KOhzBF9sBkLzhFm0EeTxW0eLUJihzVDdEvv5wnoFaoj7jcl6CpgWUe8H
7SFIqV7za4TGyfTHM228TzjM4QvDr0LPvofoRKykliAXJfTB4kbAgP/4+b6yl3Sw
v0ftQBcB9s6j9BxsMY/It/APkm9NGw0O8w5Ndgtat84EQR6a55FSiU3/ukvLl3RH
YGQNuFKYCZXTX/hwdQ15vX9TCY9AJf45GTXXhJb8EosIlIdXmjroOwj1qQYs2HeM
NHhaEpYePEyNEYzrmgWQl1krM8n6DtapQIyejZHwEf1pmuYi4WNQa99vvZ9mYAL9
QGgDS/nYUREML+Dbm5CUBjILvaJNYACXe9QAMOJxXBTj1dRlRe0v7gGdoKamc8kM
qNHL8/FGJVaeKRfN9K/kEBHhy9bJirHAhia3UuYLXHY=
`pragma protect end_protected
