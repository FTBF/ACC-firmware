// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 03:56:32 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SI6bnSWe0jGIzixqeOo/UOuKFHQ9+vsaFil2flgUqYKWRCmoFH1DHXoI/EfWzKe6
vFEFI6+4/5WS1LnFYatWwV/lWJ5UGY7XgF9q3FQJ3ZNFwW+Dnod5SO+AFvaRtpEe
xrN0kijBRk6pycc4/VGk9+Yqj9XgYq+cEpuGH1euatw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13568)
95u/Bq/Hp4EqyLwh4qBtjiVsIQ4IAyoaVak3xyIyqJrlFD59sDUZsdN2jSsl5624
HBMKDmp2CTecze55wiAG+rmm+qn3dah0sGUhOPvwXgXVpziRXBFp/GZHqMTLyMgZ
SpGpuGj70jLXF/oRk+BEAn6AQM6XB+QWtMphrQV4Ojm2S7D/NvYqP60gHLjMA7A+
PPxTjamzCfl3kVjU5hp/V0Px15zg1+VTSlDekc7xCVXFOuxra2vnSEpCUayx+Eia
b/TByldAEiLldGethztVjG5ZS/5oeLfED4R21OQxcRN1K9xjbfQkkRLFTBQx2sqp
u+Q9uaneuDiIrTpx7ueuXnmTxOXLa/7xXqkqjQEX5JpMiqQjcCSDMV9lV4w04mT4
E5yJ0Rb1Ihz3eCknjgzJ98Z+Pa+7Pw0aW7FglKIizpYT/lI7uHsGP5kLV155AV1C
Jjut7N/LyidTQbJ6Qn0Hp2v9H68MnEgMfaVdx8Owj4mIBAQpkY4vQjtrjXOUg2fO
kCzxI3nmHkGPYbxOE/F+eAVnP3SHpBPoGVFsd/9O0eGrNAN9RPTo3mGsH+FJf4Zq
JmBErXQP5bdkVjvw+KKulf1f1P9dUQfjJgmyCx/veUXedDv2R+byxtrVWEdMu9Sp
Luicu7cnjt70ThhwROj7mw4K6ct1ved50lrMBzF48uHV3Ma4bZwWrt/DhsQLEIMC
rJf9tryT0qVrXZom6syvtGIDzLxVhHMlZWWCAvH3BzhXViqDvh7xAkEz1D49vFt+
qM8ndY0ws75n4l902MLic/GMcOnQf7jR4m8VaiyJ4EA2KlwfDqwH/CcQXLVWtWUJ
34xTnT1WP6qP6UTuMk+5bKtq/+278MhcMEXMMOojmm0Hz6TflBZ3BGf4pf5nPBFM
WempipFhiFQJ5c2q5oy1DgDcMuBMJ0v1RgR+Dyvwkj3X5i+gwHyayEMNOREW6I45
s6ZCH4xA/7T/PZjOFCIjBTc/L62o8wSgYps+cVKURU5ww065c0K0jS0QdW6phm/o
QuMM076r/mxO5j0hLX61iqfpn2vRdnC0fhLoTYtrOoe5o62mydkZ26kXHOY8Qs7m
6mTLTv1UbDaHpC0SNnMq/F7jMoQnC6GyPB2KCRYl30bWERligvZiZrI/Ee5lD6ti
mD+5gd/u5xHFwgI3C5odNsYb+ilCsMYap1jBhdBXJBxZ77z3zo0CNm+sv28fejF8
7NlAOVP8IkPcaVaRXe+2COMDd6o58J/l35jXJQ2r7EOvoFpZDtO+LYFudfkjYdvV
19/cew5bJQi2DtRPQZaroWpOquhKR5EluUt5nZmWq0AJtzgfhPiEHPLpgvxpEVKj
52HpOmx+0YJl2MVTempbztp3yvieHb1era/Js+RP/P81ArvJmmTQYjjOkyEWO53U
PUniOdOiqAaSR55xWcvWzsQ3dGbMnXfSIgnc6sBM0q/7qBcl1GOiJkafqr+h68wm
wYcr89Hcng08H2/UXU1GJTRE+GX0j/TjASn+J6IIULqfI+b1IocJ54jS3Z3AEVJ4
rREJIuGGzCTRK28peVp/VAnGaM7lsprbgL2jLvJbENih+LafqStypVEUrotFaFH7
4jhLgkZ/1YfHbDzexaV7qo/069ypvoAwjG+w+DKwiAy+4wwQbeRs/r7FMaN7fufk
srSmKk0EevzzokekKWhxjzigtHxUcKiMtXoZlZQr+E2i1vSogbKytQqEcXDMzCHK
XvyFT29+Vc+O1ZJxohFfmfkJU5BifGKXX9z/dqlcdp0VK4DPEZ6kPCWq75ofNace
s/c9BoeBAvyxKpSVfrq7+WLlk0yAYH1mle17cCAN9Nokfc642svueihDO/vYP4M0
CmDNti0w7zyxMC2YUrd0BOrawvWZweGkoL3r5m4SWN1QWZEP2BzasebJNHOdo6+d
+l13MB1rXaifS9vn5EFaMj7MRh4Ja8chL/UJKk4LJfeUlheLqBjt07Cw8Mt1FXsL
lHhNCO6Vyngyp/y8hjXjOecm5Kbl+KzMCIKVkBB5EC9HzEM47CMONBtRjGqJxcJC
IY9wg1K9V++5PZ62cN+NP0tN7G3hpv4hZDLvLZZcB5I4I4pdUUqy/uXTYdXw1+wy
gLL28gPFd6JwrOTY9d6jCobih8PFVaHq6p/Qhzp9zqcBbYJ+oFDbN3xV7h+Kude6
LjZodCWR7ur+bV8y7Sx3BgSrHN53LIJRrBw+lEjyvpemZ+VgCY0jUFws1k69fiel
8fepKEmJArOS2bBfsX6yFH0LT8TFDhq7QI3D2IpX3s1k6jLBm+WRySgViF79uuBV
kbqcrFeTFiN3ual+MjopvaFq1fjfP9miqVa8w9T/nH498WkETp9OjPInHxMl2WeB
yDyw1Nf5cXQQRQJlX8jy753L56gsJElbdCjddYWtiDgC4iYByl2MK55FCNY3Ovbf
9PNgTGljyCuJIBS7jIsx6xbF6E0a3tbPKccFvHDzYGllkzXHbhfnggohx3fukkUi
01vlNNoH6tokU/gbuQBWQRMuukhoDvHicoyqURu5is6886T3gitfiFK1QfgmBtKF
RmDzB6cwrIytWnqOFAdKGdRFzSRjLZDGjKsOOHNbIItabtBAkkuyzewBxXx6WoS8
OWbqqR6WQ7F7CUjC4DDN63u6nEc11HvdgSyldKqrbhPdfTTdIKULFpPTD5R3qyw3
FR7Jc8Z7rU/qaHPa7+4Y5lpbUqCzMlzbhEVxYaO23/XlZLGFgpOXud5B1gSlJubW
fI4jkje4YoHCmVdkGikgymb/jDbz+lrPqmq3fOqY6zsz8OFXxYLlk+9qJObkm5f9
oEi0OOOwRQ9jUuKZlvY/80OFOMi3wSKTmGuhHeGEbpSoA1BSewuDaiTMShiPzXud
3dLFBEqIdsI16AMROaPHG+pA7klq0bXbb0uPug1FUHaWuunqOJ77Gy9Pa0XH8WiE
yjKkz5lIgawSIyBhT0Y3l+29e1e/4NZg8FgfQc+nZilorLDOmO/1SlBY1omMn6lm
P63UphdHselPE37uWwVsw8jszYWAKkEUV9tdsvstgcyeedYZvGOHua/ZQU1BVFmT
6/dgENzzOMHBu/SqpDfQjyxYMeWXpUeM3aoOTHKuWN0XXKTkRXHtNZZwS0o0WPVN
tsu9mSZ7xq9Od9N9efoep5mkGazBX4My0yP46p6wQGURIGiUmhYKNdUKG7EvbW5C
UygSg0PxpJbjS0j8wSKvdWaH5nt/VHQWSTKDY7X0tcAPjAjaGwHsDdaS84QxhAAu
7PJI4hvPpgjMG62CaBnQ2NyH+zw1yaBTMojs+lMwimlCV0odQXZP4jEEcXnSNfUf
WZFvlLO5g2u1qTGarbVPSh9mu+MYJLZDWUeKSwWb9piwFRNXME589+ZXTKa5SI2K
KC3sb1zqGH0PyrF+HuXiwZWUZu0LoIXogrF0xZwahEJNuMbQWVSuqdDKriNkMRII
MZag1mWZU8vZj95gscwypkNqQ0ka9on70erl7W4kkCD3ZEp6LFFnAJ+YhPMeHDRJ
paGz3S/mi76aGnNI9pdIr+1/Cj2y2OJl96SeJhdq2AH82ORqkQyK8VW5YxvB2wLa
KlhC+WKZz7fW1mkdhxBr/Tnb47TDXWoTxAsz1aJ4WESqs096fVlzIvfAjKtiKpZJ
5BeqgAycd7pJ2vcgKoB9yDyFUnsA+Wk967bi4sV8ZRiNg976e7zsFliZn1e39Zb/
Kw9NHATToJFjgKgV0Ht+uQpTXPMAWX8w9kHxSaj5w/6E9kHX+zJG5rx07+Qcyk82
l16pgSrMl0LiApT2526AQLfKNnW7m6dAouHMfi/hOfyddjdXFVWiHk3GY7E2SPWJ
woR/MSss/SUe1E3ElQwU2Kl8LNz6MVRyca9doza4YnCVa8v9M9BEKTvc7tzK1mUn
r5236MwXjJM8MpmD3YRI55FY9R0J5rTLl5A2QwqWJTvUJYHVBfJKFyLRgWA3mh8X
ikXFxcRnU19POzP9go8jZ5Ihn+ChfDqdfiJHyi+wrcf0UjN0yxOWS30P9bNjPwIC
8VfjTqvkkCmC/v1jXkjgJq5osAU/fwS8vy/vcFS26JlW25XA8Y16MLgosrjAkYJ9
eslI1xrX6SuL1J4iDApdWBgcU4tjR2nC4CVNrvYGbo4ARbj7Yl0svl+asvrnWRrs
CXkJIgAHUpyKEHK6wB4qp0hZTpH8PFfx0EofkDzjXjVSEGF9e6FybCioePv2C9PE
2wowOSrdvQhg7chMHBf8JjwlL0T9LrMqCsinhPdI+4yIEVCVC/V4sAXigntnxtys
4XeDvnuNhv80CS7WQTUqLcQ0Lhkug32Bct/McBXUGdSGSD5eURu3b/BuN7+ezT7T
r2s710dZDy/WttnVyagzob96YpQKYCAwQZyF4TCXzZ5lcRr8zPX2YBRMhTOQvPlg
AEXrEnpcWReK2uoTX/XzCn9MIlB7cw0xRv5Bb6UtAiT2eGz9Ex5txDWsoAjSwRAR
sqZlgaxW7CmI50ycdck0Mrm7ZI8ScRkjNR0BUWuJaXo0h2id/+DVHRzpYKZRO5Tp
P0TgHf8Ezw3RzR/4+iepLQXJ2UJlLlwnC2SWB09NlDQXX/zfsqVUbFvm4fNUNexz
WHjv1nUvgkU3VJg930Wf3tQ6PhD2JvCo8PNhbTAtbMwJluG2pAJa06qboQzZz2jy
IeTgaAJ3YlqEEfOA+WiXKEwnsHvLegSlHe32L07fiSsRuXLNP6nfNAGZV11QzEA3
ascFnjihpVyPb5WVXhZ0XRmnp2JZavWtG85gV+F98GhcVMAeEDPzSkths1Agm0D1
BYqFFZYeidTODwsNU07fIahPe42nj7bJH799JXZWbUCIYaLhOkyd4OIv1ziYBnA8
qLWgca9Xo8Zg1+fiFLQdwBpz85HvcG6R6wcWBo6K5H+8sTEDIg/viOKxKeRpBnVt
xrJs4RRt3IAVsm9bQtfzbG4mDVoDLUu4uSIwW3ZCzl58TOoXtx3XjJFz0REJh++k
0UlgvY6cCcGhhVjEK2gSY5hJzZGTp1fToDI/1Io0FkFCgTbbbhXfCFz5Zq+8kgED
mO1gdsHYEAjO2evdX/nT4VU0L6PC6Xj41l7ua7g7pRpXFzQVXco6UJOylDLuvsPO
L4tptj/0LTHL+zIqHHs4313nfBFZZ5OLJM33OwJkeP3RyyDXOhS71S8Qwm2L5lHb
dO0/M8KcKJ400gfGLQCq76S+SMnijsLBfAzV0PtUtiasnBe9/wJWNGIhjnVU6Vlk
VA6lz+ZgvNQOcBbAd9bvGtb4Lufen900tSeNBFtTaJdmoC+lyqn3S3s4XbRB51Fq
FGZ4wvdAV50nJqzuei3FUL9JKTdiDOETPqMCaFnujU+RM83PKgU8WTepyqQ5f098
iRYGQz7zr5xdwtl0npf1g+/+PJG1DDJEkpAd7OS4t6/LagHqXDCsm39Dz/ylfvWz
YaP9t4DPX9yt2sYn6IR1YEn1UxN97ERiu7UGt4A1cYFPtJWOIBN4MVu1Vil0nAmQ
v9njN/Ro+ksdGIk0YMIm+ahp1zQ3aiTWxKG1WWWl9JutIrcdQJuoCP0MV5iNRvch
iFOEqgJz86QdmvvFlnLE/IK41n26OZ8goY6A3YbRIy1nNBB5nvpnafaMW8wa1UcI
ae8JrquYhZYevOtrr8uk+SbG+n1lYfFbuS9XKRn4XH4Tdwsyt39trB5c9XJ6t5PE
jLaQ/aCRrRf/jX38EWebReCwUdyh+dgX2J9+04EZWwiMt8adGNjhsn+UzjGX4Qx0
5tVHCbfCx/ISf+6A4Ty3aXQjTKHuPUOJxogMPBsWNhdsehPQANyTYG7JN+MDxvE0
8duUmyI2aABdUMz4lm4rGZt1cFTmp5t15R7WpaomkGkmI2adYgSlyh8WvjA+GUAo
Nc210E+5sMD6Ul7rnm5kxUbAeOZeB2TGG4gM1rIN0zrjJeBg+/S709x16AfYBHM0
nFMP3NAgoiF2ppjjVTCmqK5fzdUqPvgBxaynnO8HGjSPShjPk3/iYDZtE1HZClAB
IlyrcCH6csF89JYWQ36nmGnxJfryhs9Zv0QqFZVu5SZU6buOUFCenXD+TsapXTlD
XWU6d7G46QMG3XVbUd7igtalSjk7kvmHOcpWmNel/fL6u9eaZsG7jHjuXlGkyHsC
ipLwpyFZ9CQTjmyl4tCUUXbjOxVwvCnxyuY/eApGpeT/LEzRsxL1V4sfyp0VTte5
rlMB0MN5m9RiL1Cwzkpvwab0iP103QQ5Uv0stwBedw1laCG4vAYVBQzq+nl8U4cw
OtPK5JcA8dEIqXqN1aK7EIyxodWgis83qMpEL527NqikTZR4PPPDSo/B/562k6lN
s/tCbUhAT69L4+SfwfDoq61qvx1qg2qek36x+bKBBQvB7A/XN7G8zrGfYVuquJgg
cokv/TG1CcQQvKHIZKXXwtfZIpGy0t0o8MpgOXSRejYy2ua/0ZoVxoSfR+cGE8c5
R7/KbpQ7HucVzZmMIQdZNPn/xn6Z1KaZiXv18kBDmcQovhogtk1122vFBjPfAEZV
4M8oOV91XXKN6HLr03Puy3W6SHJ7kDXI31s6VOd/b8sp+jsTVnHFAf1xfs17yECy
1IGnlibOy1JkjRr2fcfLact2RJh5oefHIhmpwM3ybgEjMCmqcDioXCwXkyu86BQ6
sSmsllIr1xQrtSk4NLpxbv7B+tXrSv+JehMBEVeeWl8+bKAIlQxXGvBzn7Llmht7
C+P/tEFO2CYGU1DNTHW+qnUGgEXGsJiRF1VoxI+I2+A2az6+3EFu0cl5cK4EmMDN
OfitMxMaGVKLs0bF3XSRmW7f1zn1g9jSCT4gx0bgJtUpL6q8WLx66wegSpCkWjGF
WPwb3yqtuRdTpbMT9DnCqE2vydE0lfhqyhAEth+niNbHZyoy6O4pulr7VcSSq/LZ
zXhnB14AVwwhUmDv9OC3M/nHU0l2GSRLuPHlnwZvoPVeI9YE64F7GpF44Y0olqu9
gbObOcs7ATg82L8WMyAOSIm/amLJoAXAbDYIqOsKH1RoApusXi3FabuFfLbJWPXb
jsrsDSKawjh7iK5xR1Mz28Wow39VPyujlDQcdw7hspd/vDlJdhGsKlaqWwz7lC3V
hM5Js9w5dUV5Ai4Hacx0FCP2HEnJ1flVjMtLSdNEiCpX9WHJkrSzmyae9K3D4TFp
ouXD8PWaV3zzW33bhvhkdrSPT4j0TL+J1pb0jMMq9vPn5Kt5Mb4P3gJvSbvmzSHk
3yl4rviJoCf0IMN2PmY8tTTKgkKpN6HY9YziVUeF4d2bgnfiDPLzxl919jDfUThZ
l5+XgtBtMjrQXm6nvk6ovXJuT5Ti5oHoR+BNkWD3yo/FbQ+mE6EtUsMXnH/5l96I
/jCe7wNJWbXs6cUgLhlvFynMjVRD7bkKkjGQ2GHn/GjxySWPNa5zZ/NsTkeFGsSp
9gRZzEq83coieoRaFJ5ePbrRWGFlb7gath7KQ4M74UEYOQ564XJNIOiSHhCbvn5b
kbT6+blboVzXiCo6lQhhiaFuG15CgVq0dRAee9fRBEi5WcP9F9swfmEkqb9jzIcz
KQfifC3I9/2Tln8xtjkbZ+pbwF5dk/yfD5dZa5t0Z561CbzPiaC+K1TLYIVWToM+
ZWUGtH1rwzbekgH16yNh0RisIZ8Z0H5JlMz0hK+7q6hO58ga0DdyP3udquhKrYln
pKzu6Y39dwLawozuO/8ReVyZ4i0qm8b/fJyT/OiPVIoUZ5SbXeKV7rEnzA/QIUOr
cyB6SmalEuLXrPjJPtNGVXjKjx82FbJQPPsTKAZvHQkvE4UeeD0EUgPMIdyShf6t
N6bvNZpygh33dx7zhTp191DCNEEis1bXezwnPY3wqcrQ4wwbsurcTsz6JbRn/ODy
ml1q4UpBuiLmfUAMG/qPkcdZk0e53AkLUL811i3AwzqJWnxLl2EJzpgZio2tQWC6
cUTUd0KvpbaqnO+HNy9mfVahaRe8gOLiIdJqgNdYAGWMQfAGaiyGBLN/nxt4bJak
N25m+2JzuTkPB0PlGfAw4rEa302emDQUZej/5Z1lDam7NTypCjyEhLoZXPom1UsV
yvlUlGapETzYb43ls88GmHYpAfpPocxP0rGwaLYwFF/OPTJNkaJkSDrEcQJa0hYq
DZt3ws9cYWgZlwKLb5u8T2byk2xSutBQap+BIkwipCweqC5SOYr2YnZFUsazRxb9
xd+K8tXKh1ZVhKh3GCmzMsPtN7cPEnkfplqsmWDY2e/ORa1D3XXMa3N7DlzsK95a
MI9Rmq5fILVZH1SDdMv3TnI12UbajZbX7VP+udnXZetpYdCfYxixyMaVp9zRN89d
AxJOTXZP3MmJQYp/DeutHkZf7AyMHbqtOgiABBTH5ID2t6N2ScOnfQiKhgISiHqy
BFM0LTq006HoQ8XxW3h5SEaj0SWb6e0t7eUiyaggicuwTl0xXefGorSsENNV5WuC
xMiR4QUuRYeCcPoQhJ0MmTA3dPdfYEESpwmlipGVncmpvXmMuFGAJJBFpfHwVYse
0C7KUl0OJpdPQQXqvSmVCmsNOz5UI9t+1b8D0TUQpxidG4jDf7DycYnJqigcGxqQ
fY8OHWGsivo1A7guwKYUeVO2qDZI5F0+Fde1h+GrL1wadi40LEqXqKSOZ/VppLRr
8fYVOOl3USvDmSn0yZ6Q9yV4Rs4Y6fg4mDzJJb1e+bSQny/q0HzaKqYNO4l6I04H
HPaA6cPP3bgt6c8KBToa6k+Vw2anzNfvca5YamKBxtlZLvAwXJy2PeZ6t7jNL/kx
eVTNysEF14Ufnx9VRaPJWxjxkSZCpt/ID++ErlTYeWU2i0Egna1E720Vnc3YwaIb
qLtDywEu9xPXaaMezYF9sE4IEy/C0xSAu6A1I0dTHqgFaqu3L71rrCR/zXRZngfD
G0YUyF7qKP5XtN9PxFeDsGdgXdoPN+GixPGN4C/29orgZYVngUII8eY5ltBU9jtx
3xi6fQaCLi0NRHoIoRwubKnPi089LtXFPVye/AM+0BTWVQOAcNFPILzggEmorlQx
UjBabCNWIipYsH3+JxAcUY2JxDSViJgpOhxk+t18diUXcad89S4LKH+EvZWm2lZP
zKYAa2719JJRVd8h7RiBcWmLj7QR58oLguA4Ev5Ih4/kPHoRF3t3UGT7SzTDYGk/
NxyohQschv4uovanQkagSCGASj3joDyHtE3jDn1rxipAJpMxz0iSPEAZHrORl3Tz
AcgNRqow/UwA8wDxr0rKwrTLrdYasafJGxzvrTTrzgHvferw+vkj2DfXuMLLtXbW
c4LwxrVyrEolW7LV3AWmfrXVlhDE/q4GL69/1ld3ffB+CjWyJ8okKbcQXBYo7+XS
V09ODYtSVaGTP8POla43hKFcoRr7cqpP1fnYKitbfKXg80YfjmXIuryztjizX6Zv
5eUGDzwfPM81NSPEOORj2cV/SeOkcE4PZmPGo6U97iCWGhTSWCH1RcjeLSvAhBpa
QA/NzjqMCJt8HbLhl9xkx9oQ2HXvJ2QHLgUnFquJ/OI3s91K39kGiysdWay/oNxR
lSGqXACbbygKd/Dh1OJ54nLjRcKkUZJnEQ00mjba7QOMaBzbFk8QxJIxNIqSFn73
aJDJMyAy6QisNMLiwfEkvX0WgRzYZNfbBNfN7Evm16JlKOGUc9sIXfmRWWapcjk4
oEWo22gAX4JRKlXb/8BI20XmLusdt68ffZj5GNpBZHCxzE/RlTZEd+Q3MZOPM4Yy
TNZDw2X8JznU1LiKAF8N8FOQbc05Pk3H6p2n0O753EeyMIlyIOmuVP5CwEqCIhzZ
nXKrQZoq+Q5jFUIHLs0gASv4KY6le4oY53NisJSddRrt40wEy25xzmZjOoTYf6dU
QBitCWgj+ReDUe8x8S10+jPYgckv6I5ALXExWMZtc0n9fxesvZmb0HAroahfpc1X
FXpQsqppXW0m1ZXpUDQl3H+zKSza8N1r19S+gNOg2M0LjNN86K90trtNu0L4siJp
9j9pYTlf/CebaFOKjDFSCLs9J7R9KUO/4GIVCz8DVK0ZYB120vDwlShlYC+A4n3w
IkrW0mbQRlIfv01G0hfVnITQq9syduNkNhZdycOfbQe9vXJgLCh9XdqzxwYWb+5I
ma7ovFWGLtvary5hXwJlN2bQb9qk+tGXSTivFuFJDcMuDxw5F7hOLUY+qeDaj+mJ
xqnhHYZLIBlc/3oOG6YL5Y4NDTsFgwyBoTjMkKrw9ceyBfFOo05tozF0/yiFV7Wc
Apadm1W7FuLAxGOnt6DO119pI0cjyqIzfImzHiQrlIwiXdC9F6DNJn/fXBEbA4ie
Rarwww9TXxKa/z0mfIe1qpFmVWpdKwUE8gupiuPFL6nk9od6lvuFYeTHw6Zot0w2
Vs8GUidMOySB3yB1wrgEkdFW9rFZ4bQYt+loqXaKLPdZLD8kYyr1/2WMt5iBI9Ta
bwC1ol49vU3LdRLQSDEBy2smzMglJVjaWUJJHExtav4BsDJVqVbESr+TEJm++Dx4
seDpYhzq+JKClotC+evdnYqNVeNx5HIiwuTIQJbudC+Y2L1ThJhcuCKCS6xasHyQ
1U8cSm9zOPYOm+7PQdat3p5oibJO0FCFpPRgRlTsEW+kVBQkMX9HKmofmAWF7kPT
UG5KWNfRGVsznWWsSg3Tm0z1zbCmIQ3ot/zeoeVfXe2pdGHhhcrIaiw1xxtSoJN1
x6TDRmw5ESpPlqXplyLhaTCG69frOinlVjr+RwxTLre6Ld0xCEEgCwADhJw5JRQK
o3ByLLZ06P6oVR93NnQhQ2F7qDG37OeNwAD3myY+ej43fPUnQ1hMa7BCIlWes/ur
7l/izfpnXsP1SaTq6VjWdcNgbf9/xb1szEX+ZZmkVOQwIh4iaAWCIVLRsspaPDkT
DC6YvINqJEiwH/mG6zk4IOcPnefeTHQ/yYRou+5VJXs3LhSdKuhOg3QcanlFKPbQ
tUe6Q3eTYcA+1bmnIakHASnXvNh/bZQbtHj85Y1jLC1Xe5mvv89qU+lhbiSC3ZFL
rRkF/YR/TRczE3KcurYDT6hxOi1CQTfgmBAGKzw/jZNy0LByNrfv5zSsEqkJsNfT
QATifDzjSV0PIbwarpBLEXWN7O9v/M5g54Yl5BPZiCu6txHiFAal8RPm9l8xivXy
lNQYELKC0TnXZz4DFe/y9I0PZ4z4F9Ojy67W5pwvMINnEtQvdRZNxiD8cM7dacsq
0M0DG07HNnIidqKusXvflwVDXCw6sfj+ZXOulooeqcy/lBChHeiV/hElRjSNG5bN
QcmCeegCS7HrpgYGCCF67RJ2G/0gZqXGoNL9nji91dR9LwDSfIjIYgoYzoA8HEoR
INABylX41zNkBn1ApspCEdC+qI8Cs4rPzy9aT+Hyd5XhngtKVQt91zLoPVbXRFDW
6S2eT2ozFV/6ph3X0Edr6VhrEtlbQY/kHxMRT/PUlPw78U6Z7lbRI3NxnQtLIuki
ltuugOZpAv7sJ5XwWeZdrIB/EsKE2GK6zjwFmDHS5tcdxx4oMR5H05qzNKQiRjGN
KOxDKRBBzg+mxxAkiEiN7Y221HHOtC35NS8NKhCyLRfH3qTlF5ay6SmmDsCIc2Ms
BuqiKwcpg0/Qxb8UM9dfFjM7s5BKacK8gV2hWXZgGwTyayJLy/3KUHqOPVRRNZqj
ATCuzaucmy+FrvEpSzFuDHpzB0dmrB7nH81yM1opbM/OxC34zRa02b62uGBUAiuo
Owvjhkq/QhpanhVTjnZI1gBt5FwFEC8RRfUOxxII5AG/mdoZDURA7MZ65W+GTAjw
MpG9kMYkiomrW5xAfpMRBiuFwJVupYYlmiN35cgPJdCU3H54t3+akMMofGwSunue
uAoOOZNQ5Wr9w9yrAnonvvgNT4tHguLTp3EziZ7Na3/9lRnV8KTRVQE/EP6yPbC/
SigBE5/acbvHtZCfHmrX1bOK1vtpyUuBnC0s1HedMn8mEqUGsq+n7J8tZhKsBQJi
kNJzEQB3P/Idbdp2xNglk7CILsHovyEN7bJ4mny/70CCygRykqJAl8xRamjycBIW
KsE0LC71D1CNY0meIASmXit9Qy4g01Mh3WVJXTCxgr478t5T5eqTPrxjeDFNpGLh
3aoQUx02PHCdUFEfBV6FcrI6vZsUm+XS8m8lWBVri1ZzvVEZznF+FdxbU82Vv4lc
/VgI2ynQWWiUXjSm5kFZsLwzbec4UGXZ708RGNoR5c0fpIshiSL4iSb46K/pxiOy
rjPb2AJvz5Ve5eLBxrebzUPMTV9fmPixsDZzabv84z/yuNr281Eq/Nv1LfVMu10k
v3F4SX6xAVB2BNCJVDoteJ/VhqPdM1RvxL1r2NPLrM7vXkvyVGoHL3fgvXbdlseW
MWohnadxbDLIKx7rP71q9V0adOaB8O9eFpP06v8sT3P+um6+8WabZdBkI7fkQPa+
G53yrqM4NPGxGEa8v/DTLoKB3I75MG0Dq/jApm4k9HUrtn4sCDY0nEO/3Kt7Qdhi
ImumjNu3CFIp0Rhk2gjnvsS8rTQJbu5UwFeRKuNMQefweKfKscH1HHXfO+CRFmep
GrtSTAWjZ4zV1P4NC0lh/HNTzVk+GgD+2W3xCHaeDMG0EOcGrlbK7gwjZZtt0dne
PTnkq3LoxmfIMwiNmc9JB0SrUNyDdfOqylquTOO9OxT1s/EM4X98fymo3nXqepDH
9KxyvOEwWxKOrySamjmFZhZlVCCEckfz2ae+WmFXOw3istgw0tVFv6LJLmHxa5u3
QwgXbUaOiJlidkPK1OEoS56ZLUgB+0x9rSPGr7Q441tt4LAdFVJuBUftbXfK0NJP
iNPUU+LECBaNudUcwk7N//bygvfVkplvh2hiJHG+VuUVJvPVMObCF9+PJF9i1k52
YGu4zbk9UMwsn3kK9Q5A16k9hyrYKjlBS5fOkpMZoIupD9E1vnT8t3SaRussDB+0
0CsHB8Cujb7X77tDa1yChkChNLczAPGW6nS22BUG44vfrqFkesrn0AeGUFQotP+I
Yn8CZHNCFvMCNxzM7TwzDS3VydlJP0YE54+EeGS2mJTNQPsQyIDULTeJYcWwuWYX
KxTKfWiDHHKuFZYh7xTl6RLwvi/GDtxueJHpLimZUw+zdAwahvGu2kAN6aVZFxOY
N1eMlfSAyg81ohQc/LYX4YzpT6inB20m2CtLybw/UmdlI5CJXI1GjOUs06vKbZHg
SttNYXrxBISJj/biJJ904FP1mTBRyZc45jST8k5+Va1w+1N7dRG7NhVA1hjGtD1u
K4Ff4Zs4WG8HqHf56ifFUuyoQNW/PxCRXS6TZIgjPYjLiyrY5TEvdYI2CSYCUcxw
8uCi8NLCkdOwrKWnwPjfgy6yoZGvNFGrEghQ1Dh5jGwsD19z5DlkoOyiuvjFwaoO
Dd8VE2gpXOa3QC38p1dvxsuBIh7yRIKXtVtTV7ywjGcLEueDMdoyJtt0maxFhAY3
oi9KxvFqqsdEh6AmJjYHjMdVNBi9wkDUuUgT83DPfevoO8McxzdkZnhRWSPwRly5
cLf8+i8RvrNG1j8/M0et0vHvz5fWQJvyjZPp4DDbtWzwBnnJGy/ibGrTyb1V1TLJ
NqlK/38omRrgq2jyhh9BsyggJv8zyomdMoR3w0tLENiZ28OjDrIkTRMjl9DuqfMK
Pge4FOZwO7Q6eb3kumbgm6mnrCn2ulswFqa8mIEemMr2RqVLQjkNqRbn3TgFCxlJ
lCnMHpdxGZkHWEb+3dSHE9DZqw/21cMYUxCUYe+z7IPdfDRWwvRej4Ab2yubqHkp
j82L1KCAStNdXs87BwsDpddaXsjIP4X1euIqcdH9LGjA5Beu248uz7xFmcNIaOkE
WNGXr0eGeiUTb5SHh6temKcn0Qb6bYI1cVcgTakyhdDSP05MyhJewCsgVW+Hlkrm
kF+48YCrW9uMlouhC99pMUJupSXLuR3ElSpuCUpXvBxqCd0ci46LUygvuB2Ptk7K
lGCzjOAmkMO5rOxIFYbqDLsGwWEpXxWfN2rP8kU8agEEn7MVioKXxxwW6AGdTp50
Cl2zzn1kJpGGuWu6MmV9jrSzTRNfjn2AI+uMQogeCzAiF7T79VCD71wql8iP+XfY
cxX9IzHXf5nVLWM/M2wTgdbNwLoSOPwVgWuQY63HUFyfHH0zOkQvvkU0TSBta2JJ
I0XyWdEcz1GntP4+UZiGLzq++UAGIQ4/M1EM8QrqVFol5eKxXjGhoho8PQ8pxaRt
fayBtT5TFD/fm5nWwnTKHOShoKF0QC3j8Qvpc4dq7UADhVL40GvDTjd2qIsanzIN
NzW14vfF/7W36fcpEN/MCHQhMv2G68bnt0i2YWpJdBLBBmZ05TsAyGChkTrv3KBM
XSAaaQ4O6ROkwM/z2MQCTzt5dPEuSrR2JNAAN6Pgwm4RSNnvXtlQaAL9nrcuB6YO
tQCxinY3qKHUkJG/qr5J+Nwn4Dh1TGTpkeZvV2W+SDwH3qTTbLZaGB+FQNaqGTu7
eBX8tDXcL82C8H9ChkjAjsGkGxUyFnPzSDrca9D+LlrGUksqyjm3eLSFbIygvif8
dCb3PCmswqNNwKRqLRO00CJiSLNC0pElNbplaL2sQt7OjELkGLKlQp7mCZso2qVW
TeFQhXNbwtAb6cTXeaoVQDwrcwX8CKrW+4fDX9s3AQA4Rk/MkXZ62oh9gT7ulOmD
5+Ej3+sMXXCfFeZ0qhsyVWBC8e+4Gl9rDInl2YHO+QOrnayAZV3yPSL6eLfYqcbH
kvvr+7yf2S1/XjKu34SlDMMY+9biO4CGuo26lBfn4P/dvfJ4xj7jxpcghrpBkKW+
+Xpq3MIrKHWIMPTifexKIglEixuoAgEzbM6fmg1xNVZ74PNstUC0IzQ29Ak/+CLT
0qYG/GysD+MImGkPm6qzBi01/jAFENCWvRwdKMQHXqB+Ljuish6l3LHEhrE5TJcj
WCtqfsShnNAp76hn6WzquD2Hw44xk8ym9ddLYBTHtFPjfpx9ADfdOoWxCK7zIFYl
NltW04dJnjsK5aqygRQMNQdmAadp0yZwLLqKTbAgBWgEosQiVlPrejJ37XBWZ/Ym
AEpNs/6EKAwGkVjTPac1W+Ke14ewkyW/oDuVzRC8mYJFDzNSzMyxuufbdTr85QRA
81GLPlI9fp5hp2yOiXfNym0lLik1kYtNbJfXhl1bo3Ah28kpdr3AacuHT5N4Nz4n
+nFXbZX7fIfZmWa6WV3dHsDEV+Ks3qbZImCuFNqaz+BKnxxMonsERKaEQHGKOssV
3TzEw2y4P3rfh7s1ftimetXk0deTUZ12a7ZcvGmwYhau6H1mVRrCRJM6X+bTLQzn
6DJN95MWqFofGfXw5NsiyfunxeHqMoC9tYXOs8tKC5N710gItPgywosQ16nM/fAY
zI456VKIAIogqP0qijQYXxYZQfBah397ln8D4H1W5Ey4/vTmvHi6FVhyEoNed+jJ
rhLhefVIJ7vPKSJRJjs1MQAUZGB0PX97WNS3rUXqJ2vDbbrOqfe8xPcYdvXyyYDP
fIV7TAs+XiVaxScUcR2gRRG9qUe0zEWBoacr+A0eR+Ix7zXpbB58Yfi3mo6/wl5Z
sG3urkTWWeTY35ZaYp8ztD/+Sg+yWNr76Ps7+CHlRp7XPdr0PTEo4Lj34siAYZBO
sT2g/p6uNV3OtLiqce9aEdMToyKobHrW8ZsFCkhKwCsDuYy1KXPkOd3wF3C5EBv2
n1Z0ADb4GdryVLQeB3lP6hyh+SAZ+SqPH7JAj/qkkhHxp4uciZ6lkTzs5xl5hilO
05PltFGOewKf/x1oQCCn0bJs8OKxwilO5IDH7kLfjJFSYY22Ju0aCTdg+U2Pd+kV
/2rH7Il27PAXBT50tihMrWb0IeYP/SPUv26OqCf+E7ZfiHla8B8kY6YeHxxYZzbJ
XtlUrFPwibozusQZEwwjTWvoy15iXEmXkYYAlqvJ35s2c6Er73G6sp6dXVew0ejM
6KRejuTa9HL+uqjxg4lpzM7iP53K+18QZN1R7zJA4Y+CBr7a325qoZ5W5479qYP3
p7v5v5qkpu0066fG2vq6Y+lJL9CZC075g3kncEm+41NfYC6ixLBa2qqoGGN5Z4oj
WmqBoTKclsLjHxHsw67tl+0FdWENL62A1ybAv0kZP2bUSpvlfr7bKjZz1j9Jpw6u
wVY5Qc0kC2wnoXfHnQlMdN0YfN8txcmuEPg1hyjlxGlBy4cD8pPkfSb1fOdx1HoV
EP8qHYbBzdvT4bb2eyHKJcyHxDGON4Pt4B1nByK8DDV+H5+I8assJhhrm0ZNK5af
JP7xF89ZecslQbbOGkr1WguCj+LYcK7XWCLz0bb6b3g318RlbXlV1x0vUy9L51VU
mUY4LJKvBolrgCji6x8JtiTPEg5grbUJCJ3kDSbsqjziZRvlwZxD4UfQcarAb19n
c9lYVC1CKH7OsC+bz8k+lIg1jjSQuQaA3SzoU8VP25VExsLRnGtRRqpubOBDabNH
bv6NaKxIqryBwLVRtSUVsFXVchUlzNlYAIpzS1X2hwNg/f5+ED5V2/mU0zDqZxtl
wPaOwgYJeyujlfGTUyFMHj5e3q6hFxxeTc3IdpPgp7GWBEWZYM5urHX102e+YpPR
SafCyrZaTXu/caO6rilRirQm+nC1Mhj8n4C8rCCDWa8xntxr1iUvmYpKwO5D0R37
aahbinaRKKXgxuRtS9qUt7xMloMuREFWvnBtFLYmaQ1nrckLnVkQv7N8KXmyYk2v
IRfED4THrJx2qVIvims+gDs5wWMlbd/ajhggFXFtMrJjytuEfIhl4xNED76eZRWb
Sy/FpXbjFu4V0Y4meHvCHw+EOMAbwABrugKWEUmvj8raBf2SqPLe3D0Ka1/O+mcM
7Wnu3KiYmIa5peJAD7iMh73rh0F4vulY4NHyiPcATx0ByX5LNs2gcJdiuTBL4xkS
NaiRYn+qMzBp/Mo2xn5Pg1xktrnhYoF7adkw7FResJzGrMG4s6Fn0uSfW36RUquj
v19bXr4+6Ur3i61Ai42OVxBd15eYSPX9YMDodWW+h/dRcRIHbv43aG6TR0U57JJP
8lXhTn/yz0OeaIHjuCS3TZ8CliWYngL//IXrEszwLKpSqePDODa9Xevct+qf9cSU
iNcviF8Wcecc20ySMvdPPHEVxzGS32WbwDGcLg7zgkp/M5ZRxf0Z/MMeseq8AiGn
uxsxUhY7FC/LuVGBhfEoqGeKY6kfqqPzYwPkoo2ceyJabwkPu1uKlwy7+wTR0eI2
hG/+B8q0xPQ5F6mAT41xs9Vb7qzIgLBi/x9T6xgip93/6TZC++n1IKq4rXh5SNGd
y+WT27muHvlS14R5AuavhTf1Kb27zrQjtjsTZwwqCtdCZ6ecMdrkMGW7NdYJx7qS
UGlp17Ef2FSSNoSVKCfrz8Tlsb18epHCJxrPMamXJ3ExzViwj83WsjJmexH/pMHA
3C5p39qGFqFfMZmpC0nZA8Ij9a+UBKgJHuxheO4wHA5UtpcoTucfOPOwKNefklsJ
iBvWvidQelaBfO29qSibDx/dlltZUAuGxgdKdOUdmUJIfCFYfQQvJpve0Y2A01l1
I/oY4B1tsKrkFQgvJmVYY6KXTP0VQAmAY7QYclAQRDQdEWgW8W+U8Y5f2Znx2RTG
8huAKOql4vgxHodsECV2OLMohRay7m7puCb9UH9+jPhOYWf39wDw4aCVNNgcVBR3
dr0gOoT5cSdP/SD1DS2F4emqVlEONDXoBjd4fJZSa1gSByHSRGKOBgfPORMbh0oP
aieaFIy9xfYpwBnpPvlwWAD9jUL9Fv3U9IpFi8NH/3rGguGg/Tg5JQzuXCQZu0LR
GbxfmoxYCjhT7nb2MV3Xo1hcKtXuL0YzDnroR2lxHJU0oTTgfbI5TO7CRnpMaIp4
wX9y5DgaUqabW2v1P7x0MHDLIaDQcG4PkA5ZLIkereXqvR8yIpzpJEOKOm3Fa8CT
8N/yB+/dmCVUnoMNmYot9P3ST+KiFsFuSmk3r/d7iKQ+1zGtgsj1dQOB4sj+dg5i
lzFqJpGecamEQafcxvlDLNffDscy1X+Qo8QYrJv5m2OCiusoYD0cJj2sZlDvzzlH
Cpi/WPY67jrHqQrG38nfig6s5GXpQX+b9wvrxw2p7Kw=
`pragma protect end_protected
