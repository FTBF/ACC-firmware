// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 03:56:41 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
d0EGLrT0kUoaFnTl1M9rRhaxnCDzA6oELE3cpeKiXLdUiMaZKZAxZ3I6pB+3vxrg
Y3WSoAUd7KFM7y+nWrMvgq+ZEZS8QUW8Pj1r2EGvFFaf5Sl5jLSmFk5IvTT+/QoD
W3uOE4H1wKS//lGmCjuss708IVU0KF/LNGXcvLal9NU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11632)
ewV825Qq1xTZ47AFPQZht/Bv8yWJXnhmh0jG4m7AIvZNrzQENhsA1NN+Lre/kog8
IT25iF5Z+Xqg8KzdfhIvEbNazV2M9X+J/+bC19xUrQZYgTAOI5bSIb/uY39tgyi6
cWT4HO6mCyxxOlrudZdOENOfE1SpXxPU4KWguRof7Px+DZNgD36qoybi+BW5NnwR
hvHIAxws6+xmcyzPPsPSJVQFHNiYdPZqQGRl2fuMeak8B8waUWN0w9M5DumwwHVz
gqc7ZYt2TvK/RD2v4cbk9aigFavwlKb2Yd3+xnWgIYINruOu60zAnsDvk352BlUs
NvLmf9p3ZyQtCzICTZQrIMc515sziQeggMrsAi7mDgqfeaz+eSvq6pvFU4m219HO
Uh6/SegxX4jn2W55iePSWRSS1YqIpYMdVCoMiS4iheZKEPOWYpI7aviavjtabruq
sQWBRiKyO65gyEmK6SytoKeT8shm8P9w/R5JLkgJSjjrFMKVYVQaz1pmigGg5+n+
kwyOZE2HhUFAuA0Ofm2WGKZn/zAOYRqjtPa7k5HHkhxhw62wmEdKW8pDr5GdQqku
x7WON6iG7GGNxl9T0iKGdCTnYF6kOrpuCoE9MmK/x6POscnN9wuQ9j/to8aT8ADS
l789wPEurYs9uPpmKfPHHV+lblQbyIC0rluan1Wu2nnIOlJPWQIKQM0sOwBHHC9B
crDxPX6zf0zpuq/vLOPFfgMVS1MoynHl7FZZaR83PNpw5MRxKE4s0IxbN4xdC1/L
g/ynBEe7asZa99UiTvPsvBIp3U+1u/vpAaa6H0KRvzBzQ1rbpm7adC031kE42NrL
I8FvdgZGmDctedGuvHaHnT3+nJ6TRmF6RVxXQp3U2pf/MNUKud4evbF6fv7tyKcF
z6X7ArvQF9Q4saRE1vFhb01aXdGjpIBsaBGTyyFFQQ9rl4qmPoiR0OtKYEsxn1U+
cLN2minqQ3OAAm3coUXj4CvY37R3tqpX907NDYosuoNng9YMJyCWt7d33A9Jh31J
T5pmMZUpsn8OzkaM/wlix/HO10dTuZRT8uUMViYvfBWzsfLWuJRVl08xoSkdhl0P
iCVcqpG3FlaEPfGWJOV5WyNUe6QOZLYGq9SkAqctZzj/yl/ioy+BJiX/QEmZnsda
vi+JV7VU+RYS5i/AsuxPpx9Yb+wZHsJOkyM1xrGDmcgBC09eUAy5UbdEl0dKWf8q
a6suqyXfhxVxQc9SQDjwQa8uJvAHgANE8dHeilenSclB0ZMm1F+uKJBTAVtFmX/T
uiXcU/kNZ7LmyZTWToWrWPMAvA9nwkBz+WsbB4tJV5SRqMY6rWkbPHp3RKJlCpzz
HHUIaVzZZprI3JmI5xhf8zPOAOHI+tD6FDStGeAm+SBbhQEPE0k4gBSDDmbsCQd7
xtfbUchjZMR/ABcsGUeZMlYkSKftBsZouHytx8R0XWg4bpwZPUDTP3ivnLJNN2ph
so3XdHES/JGAy6Vyrey1cmsIyBqLEQQyeGpAbB0hmsq3f3HIKK0hTFkhVLjAG0l8
Vnn9VxsnyGsyssOAcOPN/xQm9CUbq0e4rRBjC3icYJCMIWGjlMZw54RWaWWqmsct
1DJTSffeZDCyLmsi49us7rOdszpiWU1xCRgIYbwxXHs4po4uYprpjh4JHksb/RHL
fiOg9JMSK4Ax57m6jeK01Cq6byGqcT4qeRmRHPuQPAd7V3y+mArm5iZ2A4bcl6pG
WV8rdFEZQn1mgKuflrfXJKyeSQc3XVK8sU/UFySpsfAvQe7gvzxec4mYVfwheMkq
LIhDUrN5Yl//isIBPn6P+DYA81iq6fe5uZ9vwlp8UwYsfRHIU8ANqVuxiMB4KZ45
7EhYGkNxQxqx3ltpIXV/1otFF/TurH9YDSFlyEXoAVOfKT57qQ/4EAbPptHbwZ88
jYDgQB391sFCHngMKYYFFRHxIymv0mc5ICGcv3TRNy6FtcXIl0Z91vStYn+HIRj5
EgayxKIdJNoIvHg8JXQXkTrLM6Q0hSPBwTIw8z9s9YkdD9aTQcynasI1kGx61T+m
lj03LClLtP/HFXubnvGEuXpy6K8OuRy8qhVvgwXT0GQn7rEUf0aV+ML67Osc7eFO
KQDIQIA2m+LvhSHDjhgV7fNxW0k9LPBmnoIk10tSQ2l15oX58AcmZxII1tjgHx19
OIkBSkIOwldlo+hVIcfKRH91LYKsf0jYdK4YCLUUkHXMZLL2nDVcbNWkthOzHEjG
sVMug88j7ria2Qx/BHd7nyaRlH+y+NqmeE/ijFoExYNTyzeTvvBkwOWPZOjJNeZu
OxvEVLVIEGJCE/VacFOsyzPY06FxE69Gg9zA4r0fVmwC64JHthYO4/wIl3DPffge
FEc8OK18hPL0Dun6mQP4r66fXAFLPFtSpGp7e01aTw7k++X39KfY9SMWSKvjN9RF
ZxFhfT6wsqNe7h+PXCyTRWcEs4ec/CP1wWDILTV08DMm8R8dy0aP4xiqBIvH/NmT
21qmYrObQGcxXnT1P9tSbKiYw9g3i1JeaHajeO5Dp6kPxfWYS+e+9+rnBt2CfXe0
CNUXLOXWRGYV78nSEVxDSK8x/cUB9fAKWndIV1wbxyxZeL+CKjKhvLPcEBM3aUw6
ONhWou/b5+7htX01iNKV78ZGk7PFwqfIA6eXLWuop+bddV6/mIkhV0HdUz58km4w
A8Gulorxua50kgaMNCLyCaDn5JWif227l9U1j01p9Jyuoa7apAe+euab8Uv/LJdD
Zyn3E7UC4+/1Rqc9tfgxoLqtYkTOddfGConuvmkG4fE4EOK09S2Dy82ZpbyhgoPS
gOmGUiftWg8COSb+jU74MTfmsq3ajdKTLnKNlCG3Q91w8DRFgqG/06uB6ivMENeD
j7hRiWNvy5/QWcfES7mKMQyLH0JatfY40YabVBAfolYJObAAD6EzEhbLuALJY88m
jHyUKgpBc8Gr/M1sG2aMWLK2muwD2nTSvMFn24/vWTSJ5pMgLZWCObHZm+dg+GUR
EMm+ego52p5RMyxdMztqoEPcuJoLUzXJL9dVIXQGDkFMdQWpWpMPNbOq5pVw+i+A
fTKw30kjFdrffi5e2X6Xc7z406pyW7rLPj+5oOQJauh15vPfjHKEI6R1va8ewFRA
U5b/K36t8zHjnnDb6cF6UiCfzYwZCxMRvlV4i0Zyyv8sWyuWU0LKB/+zKvFkdJAu
r+kI3ugou8MF7YJujA/Edw/Z6KTH3QlmMGqaa5PFkS+iYiD+GnUFzPi/6oFTHrcZ
uNZ99KV68f6vGesPIXsSFyBAs9wb9FQIrI8NJYgX5muJvZ+bhtwoV8ImmykogQ0n
gKldHFCUSfHNJWghj3er30bHuInUOixM7leb8ZV8UCdl7mTySM+orxrvnpx82UWD
3YMxzNEk7ZTfOoRJyfqJDAUcD/E0V0bBAcFjIj7/ejlOHDw2V8jmA4vXJxkkumka
1NPDaDFQ5vigoJ9Y4WIdS8c5Uv021a4Zz2rBETWzpL7IHKPZ57w4nUWz5ehpNtGy
PIZoDA0eMIxuozZrhxzjeMna6yP1GTd64LXoy3r9GF1nEXWBFxCbXglH7GM5vyiz
H74Pr1z68yi3V8OQ7AET982WdNPFbii3h9KRUiOShdHbBSo7GcQ+khrV0ZDBpx2R
EJ/fj8w4W3HsHaags+erHs7fJ/lKDMjhuyE9UFvCBVG62YDoWY0UYq+GFlMfo11q
F5AOvEpr2nlRGf/tvkLZc+DW6jlFqkBAd000RLyo7X2yZQtE0LeV8j3Q5uIz0k+i
aXycgmGWYiKSRUle88fWR72K43LrLEA9KDbj6VbjByz281mw5TfIucYFWrLqzuet
ELicfNXF77I9re4XrQQcDflJtdGEWNTN+ty7KSCMO2+hSrrWwkMzlyNhLjVpolBL
G03hQ6gzbFAU6FWeYaZgrXlNMkaxtGpI6MH9985St4qA1J+HNjpGoaJDHchmbr56
kkF2mfb8tUxcjXh1qa7yEZyYFjAO7zZORkr6UHuxTOM5XTT597B1g+InVDUGYWn5
pDV86NM8DjGN9JLQEX8J9QXtxUYqBW3XqT3QU2ZQouK5stjfribwp7mjCeb86Utn
7r23o8gmuvR/ckVcm5AZc9yWr5vVlBETD7mPQyrhF39vr2YoXc74x90VSYLYuutM
/BV+4unlv2LQhGphXUPQxmgwsvkGtB7xpzjLOsirg5ItzEl2IIYGZtnQpt435A/k
PymLQz4mYHFXvBtbsqSxpcjmFNLvtub2D8T2FfYI14QGT8HoKsrGXKg34eCkVUEz
5jJ7Kx3YdMaS9jJJRYHwDcShxcddPzIdeq13FNEuOHtgfCD8wvnYvQIQIN+xzFKC
Vy7wvAXy7GSEQoGXy6oUFGy06w3t89W3ZaMLoe0hqcl18fTY2BfqaeTkWwa9ZMvp
W58wFIvWo+NKJlV9CTprrJjERjRPBIrlviMZ93t5j7ycx+Jln0m0c4DtD2Fb/jAa
VScnrarx2+/SI9AU2XvZJRFYM9ghVow76pqksRJ5DLckqtObBaH5GMASLVARzup6
Mo7X0y0cK0R7dgBDK0vJ8xdgKClqe8m9gA2NMAnJWijo+LDh1UQA8QHcdI1UIEHx
RpbXJepoG2beVAfrryZLpnPBw+msbpnk5FaqbPUj2J59/9EFfS1aR0j+yOIohaVP
txcQ2vAVcq4xt70xUi6YVZ6WbcDb0WyLJhfIOKxUtXD/+IAyLXLBkXA/VL3V3xyF
jC/ggBmXCqkn868oXAyGLZ9Z2L+I9pyYdzrO0Gs0nHEG9yzpA9zof6e1wFJtjH3s
BK6IQvi0tuPBoYAhlUaq0xjkfAMtIfhOKoz8G3vwOhJmXlZWx2NtlaPuFGPMpKf7
ILifZIIc9eeoZ6pjU+5X/Rwlw2W9tPLubMkEINsEnHRU9mqoOH6lOgKg2uAeo5S/
JKoDTZwMyiOhiBv1YXylPE/6jOXeZ8uXO+jiRVpyTcGGPWCrp7kPoG0plLBx256Y
XeCoo8TWuo0O2RlvVo5mNyyKoO775i15tGL4cWJMToa1nT5/+QEYw9x4uA6cvUFE
qUijmOTXntrQfsJ7wv6ruM0/D4Yvkf00uqOu0Wv4vanK8pGHog/zfjTOhQT06GDL
AmE0JXbFXkdcBpErZ/l8gazv3Ruho3ZH7sEXLZyRtxM4dJJnfz2/p95f+XSsB+s9
6fsPYifniRIn4fUqVWw642bVielL0BRvQgZXzfEqN2iXL6NfFwpeNy+uU1dusXoq
FrbqhrcMAbzCEKBQM2SbS3d78CyO4dAewEaBvnx/CJLIqQ7IcBrsmgBDwHvGhX0m
HIl5rkUt7PuuGgGyW9l4vWrPd2ENfgHgT7MFiB1DM5UmOrpGk4bDd4KplS5nezww
NbKo91+9m+ADp8LG8LEzx+UNCWcwrWjw4PrVDVsgaSaIbGZyGoyJ5IBNeVHEAndk
SlhwToq3MFmfZIFBgMNUBS2jpAXM8RzdhE7PfYXsYlsyplBV0qWjNpmLX+7xsaJ+
dT4qNmHaFDyhwUNdYf3hmALM4axNOZ5Cjcso62Jz5xqNIh2Q5x/DjWApHqfGcVWj
eZVSmaYhhL3jPGpL2xqw8q4ulF57F99YX7Mve3/N37FS9+9gStuWtVjSDZccJmHM
PXizlJZSsIRjqddagf2aCme/lNMoAvd+MULfsTk1HVHm09sVsHZALSVyc87IKf9W
0y1Pw0oPcax/7VIV4NpL+zX8wun3tDghTDAlYrQ1TPJatogurJWUEsWzrpzXgA7G
nYIBWag4QLrPiLzNIxGIJv3xeh0afRyooX1nMNmZ6kp9lNXtK9XLynTByejxPZsg
eeyqsb8eNdjNgjjcDvri+1EYGcTLi/T+1nKWm6FYhFrotn6wlXgFkjnZQk99+IxG
xqpH2TnGRqjY05v4lZ0WUJd9rUOAPGxg75sXolOiUVvyRXvaDhIAFbIP5uU32yYY
FxSxlFo4N7Y8sIwFfAX6vvGHh2FLPq3CSbTGee8s+UIbY6iT7ym1VTfG8hJhFxe/
WsIB86gQZXApN9DGEsEi5t4Wa0DqCtMN6Zi0OsE3buGcUeAbjZFtYPc5uomrbzxx
NgIYanahVV+AgPBbVVwxtDBeRtxkpxGI5pRSOENmUUd23ycTDuxX6xflGXDEW5mw
EK+p2P8HqvhC9fmWL2mTZIhYeaeQuuSxVE/oN9ykkqtYnVFyAQXMoplXbdwxDX/R
eilBFXYvI8bbBzYL6vM+fwDKy5NGJ0jAf7XvSPU5RdoAGcq0QdZc00eb5L5IWqlx
dcQse2xmrs9BXkg9q02XjaLPNE3xMHb49sV5PfQbmv3SGPMcvh88SW+VGiAbkfBk
At0cE0KJnQEilqm5I4XOxohzJMwXUqFJTb+7rz4w8uOMPlI9IDrYGEflFNc9A4iL
jOQeSnbGSLLaiu8SmN76RWCunXYUT1vGxGFl0uCnMiM9HYBrduU9grlwU9BW1E/M
5aItm2Xo4mT7DD1CyLP8nkjd36niw8Efj4xa7NLWgB1/1spCxnyxi2Ne3GDZ7q3S
jhsPaaEjcQAp9ufXP/JEdtSak0sBiqtQul83uC08tkeBJByMESSxbCDCRgDKAN1U
UlFQXh5/kTxEEZSLse28YR9kcABZ/aZsrQYis29YIkPxJSji/ViSyb99kTXZ9M7D
jaekXCeKSGcF6g5mzUepZYagTrsWvjcXZC8gAqvMRZIXeI6NHR6lPVZkqFq9wjHB
XWRs8uI/JWyyAU/BNPa/M9TFCIR80QYlRYWfO+usJh3+IjGyLyks1a01uS9wgzAJ
SFLahmxqSX6MzGUJy8TsNKZeCacEPQ/uHtK/Oo8tX8DuOwhIuCF2JahQwgZOlr/x
vT7vWj4gt3bBUGMvydsj5ZdUfrVgM0ndWwvI/j/hV044OSG7TjciDnrWOp4+b4Xv
Pz5sDX7N5gRqXWz5r6mMmdd63rZ1or3UijrFcKg6O9lrJu9Yp3puo2v18DNkqtLJ
izlvHOqO/JnSfzulOnc+39oB8jK6y+odG1dQptveOpBrEW0SVtDMqVztyldJzTxP
/KemztqgZ+5yV7E1JDqc05nIode+DuNFZmESveKfBSrWRHlHhJFbL5XajLI0BZIG
HQBcK4lH90BovT3xy1N4AfQWVX1s/CTyI1lWeP9nZxSdk52pPkHmfks1LtNEc7zy
v17ye+x7qkS6kWf4cnKOm8UFhrq0Vtt571wvM1vHHztXbYBgXrFcDAHW4vGZdpVj
GKAs7ztRf5vWS4jczRpZbpQpzGga+Y+iraqIcYF5hGEnAeinyZb5ukri/QWrVP9Y
Cx65FDh5Jn9MQyzBk5XZnPGxY2j733I4zlDyzFnmVyP7Xk+FGnfRtOWdzMblk0Gw
4R8FwAmo4AHfNf8OTFdyzFAOgRP6jlizU3WMdOpHf9CQ++/yOWMeHaa2FKA0Nc8B
ZRFWqcG9qt1dZsTIXK3zEwGg++Ax0gL/N6fjZWKcAu5GB2Pej6HUhr/pbaTLmmHK
WAdsu1rxVAL9nFhZCzAl2Ae4ui2x7DLZauHnSCJe1AWXO2JJocbtgLIIDgj6gT0d
uM0gdaEV0BSL6Lme6iFoqwaN++ERpKh+HUP+lYiWtnzDz9Jd9iaqkgdC40Sf7xFC
UYVz7qKdN6Ypqsh2HXlbGQTZF6S4U2j7r8uR5RRi+7v7M/nY7AhiRpZG0Fjkh4sN
MVrBzRrMb8UNMHTtiamFfdnGG0GC3THON24z6fHllHhPRAt4x2gmBq7cqIP7Xy6/
5sX9wD9kbY61jgrsanVQt4TZS7xAJPRiBveMgKgvsO2E2id9QpOCYyz+mYKLF1Z8
+M7/zzqkFQLAilblP2QzwNVar65t85u9WOOsMOHjWYUMTC77h6ciSOt9ggcopCB7
dJj3Oo6z0TnWdQHgndduoYQaxLX6rEX2Ylf4R06W3/QRKMhAzpWeYR9o+oQVchfL
V9fp+YA3ahba5msrU/ViotG4G5amQbHSQfJcE2PChyb0K75eA2yb1FPH+dbx80MX
tR++ncJuOr5TLnUdPqigdBjAjaHPfm3Ii4RaD8fbe8lyMW4+gQDIcRMGtze9kD3R
J1+ylEIAW3NSA0haYAf/7c04alAWQUN8SL51TWMBIO0wWg0vc6l3KKJZIeMLvM5H
2Y03lW3ef//U/1PqxMvG3vDGRkYqySBR1cg1q5uO32EDBkp8UB0KP6/dC9ou1kcc
WZ1KPty5CeGy9rxv/oc3PbWP2ma5QNmQZf7FWzAj8K3QdVsPpHG/5RAtuaJ/BvPN
EOJyczHYR3BiNbxKQ123p4/XuNJccL0iqIG6ekz7/1NbPlR0SfLPjX4MUvrdDBAM
6ZpcwDmE+7DA5XMdOrlzTrZMnogfnObkne4463Cgm9FnFlB7IFXDtUJ6T66lg4dO
P/6T6MkvyZ28KcHhp4ee/ksgZFimJWiV9kMH2QrreqCuyLahohV+tZaSLmJfpPrW
ld+Ui9ADRlgb4EUbc9wgHJrW2ODdMQDMJ7UCrrz5q/HtdGDKxJDeuspEt243WPGX
uqbxhN4OrNzAPjYO/YnAYnUdw5pUqNzIOnZj9XdnKb2rJTiSA7UNCAYYNPIrqa7w
F3QnP/xqPNYTkdW42s49yEabCginoIs1WQL/8Dcg6CKGEyvDaI4/0NmH6f+1fx2e
TCcJKvIqrb+Mkds8T0kgsfmXrLn1SdK8m3QJekpg3Pi+2GqlF7XIFaigL5DdBf9v
48B9M01ySnbLHyAPzaV9BEsuOF05ekremyVHEmDJVwpURg7Sh3vDwyoFqZJNi0Gk
3FPhk1L/ztidPwdxlM2qTNsC+HDEEIqYPLQ4SGwiO83laXJjJx84+fJUEPgR2+ku
NOEb5lSjOzP8Qgex+8i4Ub0pJ/aZtAOWnEViuFwhXhrDiBGxIUslg5g75x0vbT3K
9vA3omS0zrAHtLIl1/414WoBb286n/ZHHJe37tLJ4/6dxuo/eugF3DEtdZ+R7mjh
oFMuP4bqpa9PYMWVQTLaWxZsW5Ws+1Wngd1M+5MiqnBfJIvQC71c9eYfYqjO7T/i
+330zEhmvLDT18hVGH1GYzi5TLQMcPMSLH0ndcyJNptYLY9bO7LMfdxbTCo4Hxkm
7QnCNGmwYj/6aZGACeRFdGhJHhp3rX/0oN9Uhk90n3x8tKht4t6N9AFne+ccnqQS
A+R4oRJqpYvCXkRtSH4uxg8j898Ai87gdx83Nomk5XHO2H2sgHF2QgZPnTJCt+Qf
iNJctXrCKRWu7tWIOkZPFF2QTyG+EBCVLLckIeVJPX5Pn2lfmOvME6dw1l9NbRHH
fhWBCN7ckfYXeTLEOIIIbIxixPoHkx5d5v8wN7ZpU6DylFMpfv14s/5XqeFOZds3
obRrxukz5VFIdok5oTKIhI6kPRZ1FYxEPnA+Z1TZFmxs5tKobUqJ5FhnJRfRfqrB
VEgkCS4PjGkN/3Y6jaVzExKMQW8cDkVmsTNpYOTxSS+VbCFhevMnmY3T4Y8ZlLgW
tT6CRS8/4iiW1r+UcZO1P+Bmo/jc2dQOYOorwcP3/jaWhfYkJABswd4wUty4TvYo
ZPRV0Dju0tU9rlAdoM3y/tOpuanhmzf/m7Dcupd6BZhuRPLgh80k3Y8dlKQsoxun
rY2CRcw/TOY9XmFH7Yscar1Zsr8GGs47wg3cP40vv4Adk5ditlz6XyEXNzz4oPDj
Am5MO1n/fLZodOHmwnSgrNkk8fHzw8Fr/4XcgSmjNX7JigPY5Av9pcnUcZwO6LF4
5gQX5gCD43+oaAW2qM/+JJndVLHkWxApxv9zxma4tIDzKl8+mBERcCq8Cn7VlxT8
P+LMaZKyYJPvpMF3IqUHolkOpiKQErdyJUHUMf3ppzxkpe6vjKRYUrxc/GeXAc+K
JBy4w1wz4EOGIvDAs+Z8akqTMqfuXFIVwQvifJZ7b8Z/58Y07aT7lRqIt+BwFipv
JvFNOw7z2AZBjwWIAi8NFDKB8rHs8To1R1lmUF4QyyWlOItFi6sJVJJOD2Vzr6L2
jYM+xzUyzvk5/OvecW6hVL1s1dp9Odfvsh4e5hcijrQAXPsphz3hHMYjBCXI2mh3
n/IcD5fFCU3zGGx7aqGSq7KCd/FL6gjDgs1scAMqMdaxVR0WWDabvOdZ77WwWMZi
LFg9u12tcuv5yzosfUUj7kKxiJslXYv+DTijS6f7hAbNWwK/LNBbI1Wl40a3iqMw
372/pL3WRtOSZ5mZuP+CLQwxn6+XPDry3lkBx1Sby710z6RGk/4QtJRIItrObwvk
CZa1Jp5tgbHjwBhspObnJREAjAbOKvt3XMpvkwsH0dXLPdxBMC7wLq9wirtMkPP/
VMr6qNWzfTZgrcVSrM+zlRrBLS6UrwSzm6SARmjIugOvLXSnSyFSR8Ai2CDs6O1Q
HcTWF8vP3cVWEIfix6Q6jN/ikGCz5dON9qialjElWZDP6b5qeU14H1n9IRpH1O/Z
oIY97GycT07gjFOKdpLxU2EUhJRWSynbb8AdxkVu/TVjV0qITnyBm4xge0oizERg
kbamTxGhBUpBxGy16P9nCqKmnXGaz0QRtNiAOZr6MLS+Y8qHsJRZQoNy0ATksCM7
1mTwBboe6icO0NThHSsowBTlvPAxiYIMY5ZaxENuCcwxQZGUqiRl21cTu+LFjEMq
AgrBttdc8OqpOfrs/I7ZEc53cqajBcWFlBsd3zZD16pS6ajT2JegVP+cGtt+KoUp
6Y2XCwYoIiBW7QPRIi8jXos8b6d/ZfBFPmkwttmvl4r89kyU8XdmPf0wmZoviTzG
DaffvBVaOGCQwLN3pnyGstZE0zaKi4FSHrlrft08+maSFWHbXPpXTTL4akg9L7k4
em0iaLOqr107Si9HuWFs2no8vEPY8zCRB+EQL6Pq/gyoahcZALMgAUN56TJxRHNB
wH1C0oUdJXPSp/HevploSf3R1htgRxVGD+UheJ+ORiIJM43+kw4kth7fw6l6rJlN
7UYtxGk7eUABxgSaBD8s6XdEF6AtQaYP0t7I3OlFGagiGczLENrLQ0QBt7SpnN0V
LXdhA8RK+AC0g23w+V5oe3vDVkF7fWiWf5TxyDbq6bKbYjlN6YTOjtIEuouMNyP5
ERqk2qayDxSA7Lwu1Wab1bk1qjYf+Erop8MUi9tTmLTk6rmgg0m6Zr1bbYBfIKv+
hnzmEui6Ec8+6a8VGTHwOPIj8DPhCYrjXtL2+1S8V5Boq755el0UGIEsV5uc5xXb
XSfDqYIfXaFd4mKlZaRFlChk0JJMc8FZxcLbbiFW8AD/XUhuPfLaFXpWZ655quFE
9ZiZpQtXP+V1/jr6afFeCqB4FUSECkJU/x+ClcFMtakFyY7WTHX0TwDD3zOygEmF
0wMoyEmW3mE8g9dT2IlhdmwJ9xjlJNtM5RoU1vVpgq2e7M7g/Uh3pl0ek4/y4BqJ
ff3DFO4ZauLEqWEm2NAjVFa8Hc5F4KYE5xXx52+qlM/myVR1kiUuT2WoMbQs6fjZ
iUKh13E9BEmUApZTvomoc9DIdEVP8Piae/MMVF1SwM3uy5B/nAEyjfJnHKLHxhmI
ouWwJR1vBlBPzaRg7fAnu/9b5Qe3KTSoXZZzB+SYxIl4up6FmlMjMpFDQsF5as+Q
7kBa9FiWypAEDaJ7kn9mbTF/IbJU315oGMYaK0MTA9EQ0oXQrnp+wNK0qBChe7o2
+65syKiggmggdrRG+xGf9JMEVm7CwrJ1lEUqcuMSCG4abqPbZgC+7w8cLoJC4A75
KBCRRfJiqLilVgOb1mOI3ukqhB9WLL5WJDjqmsyXkvTss3S2ccxxbn2ljVNDX+Ih
J+Dj69z6PYtIHAh4xSBnGGFKlONkKPhYXlQalJCsec6exYuNn8fZSr3DolXYQE0X
QzHg22eXV3QaViJD/39wpFdKnG7D9Nt/SEFREIaefuq+dYtFmlZKao8e8J46qgFW
VdXsLVFnEamqOm1G6ht6yqv1Uf4oHkcCz1/AhE7Iv+NTfdLFIaNd/mC8OVBkK6Qp
DcEgaqP3Bv7jZRTizLSbZPoNuruQ5pgrLOSX94Vd7bWC+bnk6UD2NVggdchlS0Xo
0j4hixBBGLPwWMuV32vLlNnrX31tR+hLPmt1EN55CTtuFfpmv1nhwJlUfgHhdxl8
AvBlM4DmPwz7Za1o6rSntIJHg/J3QToAYiWuciHEuLfpTzQEA1ZMRXVYpBRpBmgW
Vqdl45YWqsg+rG6298Bm5YXu5fiegS71x+pGwxYQjKqP36m8VyP/e8smBFoiNrC7
CAPM5kSUQTc4hB4DTvIAKfUSWcXQEO3zvfREJ1M7Ax8ecq+g0nzmMvxa6Y+ZYT/q
VMScCsEJupGztS+tyEHFBnUTzarRGuCQO1vT7+ZZBmwljQbUdByzxPcgZtaz52/U
CrYZ2GgZftg7oEf3RMC+Cd8hmIgiBFd8LOVgfBuHoBZIeQwH9FPTYdI+g15kHV8H
25oEkf2w80hqgF98mXK2eNki3NEfbeOgzCDiuUBFMgUYleVhOtdel5Al4Tc9uEu+
ct+Eap8hv23OpDhDRYWJpUOGEXlcGDMFEudNPXmgVORJVT5qM246ANCJ/vgUNPMQ
UTKAAz4Js9t8/m1mie8GMe+zaLDi75EfI1Q+2s1GTQaezn6WdId4NyJmNxPvho7t
0nDGRRHaPEjhn0zGhuo4bilpPtlMj61L8mfFDdUJefxTIFp7DdzF20NobS60UrrS
L16bbdDlm7CV0IyisSMWOpnQSBbwTsxsRnPa41hfUQmZuAs4FTx4GzI/IIOBpPXY
ZN9BRvgsJQ2x5QGJPqOwJk8EIh4rSelhxkcSwTE0RdUfMnOzl9ZNxsesDjG8rPcR
ZYaCGWkCmTorc73lqcW8QAd4tLvuDjyTFkfBpoBrtE7LtHY/V+LwdWdXTTsmSc1k
pUJ5sPn2B9H4RI/bGRveSSYJxMEZg/ULWGK6LHngD22Owp9xNTu0YH2QfzlDR1hF
qFa7zURPARLc7CscX/1A+d6/L3UfEbq2h9iuop4tnZpJV08T7Y1uLyukJt9pRgJ4
9D19HVpLwBYdf1PYOciB+CwG6jru5iNEB9cQBK1nLX0fNRRkphrPqUjDgH+S/ZR8
gdw/rgqyxerZuQSqaQZGT/5cKeoGES7eI5xgQYthELl4ukzaPI4N+HLjYwdu5l5M
fOv73aD/XYUzLiDuTE/2Xw/7GHOxJYI8c+hlUaclEy2lF8UGHhgh+oPP5IIek05+
fN/ciS41yqD8LLiH8BuSdGNDEeJOyb8/56c4quJkGlPqPBEYV9A14/Rdb9oo+VXV
6ABax1zORwL5R1MXpeUZb/8RTFwS/4nysS2SOTpmsn1/gbaINFlkdqZ4iqBZTGbJ
2sKhVkcPkicbFD4GtYqiK+SDCuHTProyws0JT/mS/GMN2MafxhVxljLfNH8vB/9O
z+tSXQMw5R+DkLHKbJVMXViX71hjbdNVXDok28rCP0ilEKD9VJq0MWNV5TXRp38m
HtRHaNfkLwsSFo0jrK6NZqvHnCv+hOb+nnrZn9iBzkM4lnzMKVhanKDGnMaPomyq
VJUmmhECsbZykBYHLxfAdbYSPNEgMHf+Ry/5GOFwwtaIyWYJRC/xe99+6JNQP49w
5Rp9J1Rm9l6k2L+ek2ZYMLbwRaStzX3y8rxcOs62lQJEpziBWcPSkPOtSbr5RFt9
wLQ1SEo607lRcU7xQAsHDziLFQmz27H+myAW0HlXwamVrkiRdKGeJ1MVbVUcpJFy
I0/rwA3Ffev09GwpTQCl7I2HOmoDlEQhR24NXi+BbqobAYa20cae2tfWa7B68Yo7
aOaU2Lxk2D39vKHCJjyelnIECsXonCWEkbf51m1VjnN3yygo5Df3+mrAtwjSVTRJ
OBCqmLaGOW84sZxe5ckP2T6wYUXUgo/ygp9aFVkHSD+D+U26BSGI8J8rPFggBd3Q
Sm5PhFrZBW4ZDSG7ftsyIcptErZU3zeuz6dXV95rTN2xfcHDA5OVoOF7Q0VjVtT2
gY7GFI/kf4DXCxxfR31k5/lO2Kp/ZUN6wDJ1rn4sXWOjGHpMjpqbI5kCRCtsGzNo
lTSDYwu6l21BIdRCkBXOV4/eWsGSZ0CtNEMuFRe2GD1sFFtIkA9DQGrTF7XzpM4G
T3mO9L39u3/07mGkgcGOfoOqlgl3Qnyd8KDKiD4szOrEMZxalPi/Dr7Rt4YcX8Bw
mVKBp00IK9fdsAAyLir7gS6Amanqo+xreJ0rzQXCTQO/cgSBcXz6tozepUQH1CCp
j8JITbXaJq7fuaFZxlxc348/M3WV5TeA7SmfKeHPBXdadRajwhNG9yET75zSV3tc
lAwPrxI+eznySnONPUTst4+TVevBw3U+gTDqPw6aK6BVIw3LepDJxAN7fVk0qjRw
+jHd6sArt1OxR+wM02/uHcV4tqATl8XrBxT9g8sLJ9rojg8MBRR4XvfiCoY0PaU3
Hg95srILYYfY3GQl4CEmndC31fKKrg9kJ5KF4scKv4ka1ag3rAMBfZkKLmKqZyIv
Lc+vyR68HxkhJ2tcMOzR0A3v3eo5zHE10hsQmGFJXSqzfYokY6fgvar00NxRabsJ
3Klzkvw11rfZPmHK7eWbbBoR1trYjdZ+veZWYh9LoBJ/YsYIbpxF5mhzXXl0nfHz
Iofzo9TRF0XCs9j0nviU/d4eIpXesjWeNfrGF/HBd5neUvOnvlxM+2t/Dj1RgQtK
PhKhpP6ftoymdn8Q04rij3VD3yqa/t/LVTzXB17h3TxPy3od+pwF9jkRG2H1xbQf
l+eZqjseu9CBNuN7lGuXgxHfmTtHcao+7xnIk2j4mDuUjJtI128ocl2mvGeQZm82
wQPgM6ATbaGDhwXv5ZMvUhrvdyzMvkZQGklTpqHul74bGoJzQB/PxWexcTABf0OD
E+GIpucUjLiwSjC4CLxDulxdYP8QgMpOrW7HYKH5MNBd1+t701J5xqO9U8Fn5y3Q
lvuS6ApcZ1iR2qQsr6WTMSUSyit1ql/9HCecByf8WqAg5QnWGCTyLAI1X6hosBtC
J2XVVVAqg5mzeM5YywIC43a2ofG1P1BB+0e/gOQb1/63TS2uNqCmxgh5AmVDePAZ
vuQqc7i2HpjFQiKb68TQgBzUTIJGElhveHAhMv8ZLUyC8/dStYImyJu6WGu7q78D
MyLmiwllLSZgJGctXUfmficEtTgofCQAgr/k7lHXYubUuSjWbAx/0XLxRthLGMRK
u566Gml7Zq38VoglrSDSsGbgghpOLQpYMt0l34iG/jfXURikE0ABxGNXmdEOkwpd
aNpktpQCoo/MM142WXyDklYp2JexNrBw7KmIyrHZgfu0aV8blMOO8EHmKpTiYNST
mwkPcuhzcRsvrED0TlEgWrQqRqWW3FMi1mnVaLs9LQNU1JcA52WMPWAwaq9oIC54
uKuxENdFKtdgce9LQG+QPDoUzEzqoBZqPJ1Wnoa5s4CPBxS40oA6+yJ8jIenKSYJ
So+Ok8g37qPSvDWdldbVbjSPAMsR9tqEGK6C2/ml476xZncU5dVpR0daNw15kmib
RuUxdlgzunE/oiY+UW6How==
`pragma protect end_protected
