// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 03:56:37 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tdpQVf+RqNe3PV9nlQe+JCHCoUFIV6dj2zRyoaDbuTUMvxzvxgjBmZIen6hD0Sfh
+hDnTerMnEaKgNjl73Z4RXuMETuxJTt92iZd8owA83wf9YgqU7r5WbuXGbgLg0DU
xL7+uv4AjNofrItZ2RKaeXd0foLnGF9k5AY8Dd2xF/I=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 104688)
8Ojl/C1LDuVvpExpix+y1I2siZbNry8SVKQrehrtrOPHMtOgZXHb9qldJyh+Ndyg
oXPIlGui79NuqBCRB5YfBSNgK5JJhtkwJ91AEsCEVIuRYL/oEgbdcNnbtle1LZgI
HyIuaYCpoI3SVTNKPsYASwQmtZufvocVK4e5EvtXPelZHa/Z674tQmSUuCxnSczG
+I7gIpA3M+PxlrXNUE0mzls1YPf6bWnKX9fq09HDjphU+wFg1qu7nVifEtd2f6SO
SGYA50041rOuWAQNN9HGBYJPawzG1g8/DJg+Vg8INY8wlzXWvKNG6SzOH/1KWuCF
ft1ZFwxLShhT6sHIpAArT1ir6jMGuy6k5GJTOB3KiV7uISFrR06pZnZrnFBUs9Tj
jWrhefwPaCcXJyCbCN/WEnbRb0qV8dvEi+OKZDeDr/GvfuUEP7j0vBmcnONeifJR
R3eVkm4n1XXu8vGyS0qykUMqHxNCO0IhEMNA8BROz9L4CO/WXRA+ARLqZHf3omnA
LiMG7YVQMELtDeg+cZ2+jPdM+lLqwzRKsbOo04obHIip4wuxVVBeeekXR8UEqZuo
O32p4eaBfzH2tIKaD9AgT4g1HQvqDfIEW5qAw6EWuYGheWEuHzSCq9Wto8iIz0np
YeXQPZpLwr0v6PdIkx3BSr+HCgYwpKovsqNXHFSosFFw/+jKWvdgFPHy8+MPL5BD
nkZHunf6AO0RWtn8NjbDyPGyVJiUAbehbNCpZbl9gK7YybXE4X/dPMi9bqzwheVU
uzYdfk9iLeItKegBKLxEmQPgCXDy7Ikutqr9ORiwHQeznT+q6QMFFMYafRaTYJ6q
pcvMCGSwEsGVMn3FRbB8Jdq89TLJlPB0Lfh2H/ebuVKmtMwh6bDSg2hr8tCza7sz
1gREUiLNLfWlH2v4Pn067vvdTtF2K1Q758s+1ElOrteLaNTLxZsP3K+d/AURXF5E
J2fXJdbl+HFeYSYhp+uCkubqayLHgDoV7DhRM3WjUoTr0icMZZrJMv2D9DVnb7Cc
a73GC2h3em3yUyEb3SO7/BIWsMq7wcb5qDJ5ZmTAatJdSDBRdLKUq+wPjG073D7V
iw/DuHiPxxfznRVKD1bdZrtNRrKHAiJnfRpUWG0u1l3rUkwoL3emC9507wjP433M
PyqklApnC9/V8r9WCnM/Y9yv6ONm8hDLLNeQPIq+it4W79ZtsisWOyNXdu4EZU4/
blOWdDEN56+fPFavQs5t1DUKx2Wdwltr9ippMobCdqqBNxiiRpz6vc7jkw440QxZ
SMJqieVzDeubQwuqD7/GcinCkmE9a30xxoEq6bi1OqTKNoJbHymvkW8/FPZVUrcm
SnquJm+x/2BIgJbmgz2VAcNXm2jRmmremR7Wg3M/X+1H50dlpERzyJJLEuLdSsoA
xrwMPBHPw+lXDUJBeEOpvNWQG1Yi1/QZ26Xnt6bbjx7Syfb6l+Ccmp7X4+Sd1mj1
LD26Ps2XeyfH7H1QIXJVuRJa07A7nESlsoKJpaUasyn809M6exuPvplxlroqcjUP
8W4tU13HRcOZNVfGSHQ7weBlB3ykg27U5b4rQPKrRNT+45E8d7l8qBisrMMDr8qd
Sd5qbBJhC68/j7yj6SlJKPTtbF7OMj2CzTmfTEWLZvu4TJ49HvjE4tJUhnZqJ3vc
D7XraYI9EDa/p2zfXJk5CKmU/Yl4HeOOtjK+vhFl29n+5WJdn/8jOOF/AyW6bto1
CPEWubugiA+7F/6VoR0enwdCyGDk1K0UnawTkJqD1Sa00yaKAjJCxsCXzT502XQk
u5LJn/tXr4PkZnchQrNVvGXRdktuKE0Lwa3sOCIYg8cd3fOSCJbnlT5C6Y3g8y3c
WXp8kwzXjsftGkyxOzNCHl4qiES65jKLwWcwtyeEzFK1hele07sXog8/POqRn/WI
CzdQ2OulkFBVpMVOFwBEJjnBWlWcaqP95cBZ0tiuriwLgInZSkqNZjfmWq2JPUQ2
Lu7dbrKREyFCNpAB2c8paoswmegB7mRfNvVQkNNA8soqzHA4gar00wTmLCLmLDNA
wbGKJ5I6weyV4FjvyaTEEmo9+qd99LQr/1k3IsGy9pSsA+lVKUkZBKS3udASGjMZ
/RoFDdK94/o5edqlouLCSeD0tb/12pQj0T0T0uB6cSBxIln53ytWag7oRJcDUMrH
Zt68II1cRlm4fSVRMYjc6syOjcI3fUHS5cJ+zf1JiIvy9RqofKzAP81tbzqAlK85
oW/0cv1ZiYgvx2kt07x3CC8TPMNdi6iz+h4Hcg4qeZCo8cMJKVD9HPU46AI40wb2
S1SG/u6vGC5eja0YgdY6NAKlEQKGBtNPKIKHPORW8XLS7pYAFKQyAFOC6IRWdDEZ
ne5T+TrbDyMO7tMDoJ0RafChkeYkKK8A0C2enPnA03tZ/SSHX08esOVZJaOqVRcf
kRa1LroLAU+lZPxpyKaPboJFXMYS8TRL0EXIbM0UuiXFS9F+VH9iGGxNpwYKKOd6
wZyt4mYn+dZGDrSDcwhIlbGsojJvGayziIw9fsFGeAqswFqUTzSNpPuydPAy2Ayj
Rt9o4EtB7CKDqVE+rMiKHo+waSXOtkkHdKqR3qbMBmH1h547Bg/PnhMgyKB/hffI
XYHgDnnDgZkt7stesZ+ZnCf1ssAGXKor/tRnqXtt6UF2DmZFmYrvlSPwUQyjmQNJ
Vr0A+gthuU8+tms9izQ+82EMOxZquQu4X2nZDbcQahrrzs/bZUMf4Dx9f5IOU7R1
vpRRs3sgg3TZMNgwRMfaUmzDO+itiNeyLe/Ru7rri/6wrFNTptaH416nw9GFS3y6
kA1gwwR3dcySByBlmjOOdqIuXPsuZsupGb6UYxEWr5OfNgApuwfjQ7TvlYRlbs27
YBpcY+7KNsk/mlk2aE3O2zROz6ZZ/Qrvm/82asH8q7TCKq92OeJB1osN6fDJOR0z
+ixIc4Hnl3jE6z7eAX6H4nniZksK564fAh66Z4Js+Bu0XVn3pbiCKaedXhrnWWpn
6zOxsQp2bv7svEBXRS14RFaQzN9KxsuJoqsVD43HtoijNdo7IK1dkTFNWIGCXL11
uoN0R9eUdW42zgtuK81rni8mF6XEbjfRTIp/D04izfbcpgcf61ZACfWs0zA3uPz4
Bd08ND83ktM+eJwP3nSIt5IjOv/PKD1I1rlN7sGCCdOwrumfkwy5pr7d84EldoZr
BEQd6i5+ONW+ax2JjXyIOvTM4YLFtuViL2vueTeDwC/UjLv/7k0OHqVwhUISY9DA
ALYDflppEM285/eRFhiFChUx6BaS/p5VGeMxVjqSsNzseoUD3nOuGG2o+BDev9Ch
emBCPX0U/UQRrLCBbBIeZL41bW5chwrk7IsWx2SvY6LG8kB43qqvYFm7RlDjdj0s
vA468gHmnJO7XLcDzdTkFyGY6k2mflN4Ztv3XK5VawfF2bskcKgNRkkNGfq1ZLKz
nTSRKFftDSH9nXImlfHUcdTDkwKa70IumJmWdUeRX1H/2LMcT916oEWq6C3BfFND
2tya6cu3rJF5L5ISTYfDPqhij2uEvZrSIh//qrNljHaanXlKzgMFLMJ/Y8htHDgr
gGq/gkerACsNlrSa0mINMorHCcGGAYWaQ/HLqNGVq+AedKaqaKhbB7kp9hf4/Ylu
gbMeUOPs75vqxBZlgi4mtzNEanfWE2urCA/xhH5z+P92XSyKX8MIutZlIEzugAc+
XcxG7drVYkFTpIFGzGJlm0FJxhbAR918mw1tS3LKItHrioR3HKdhoCIRtpMzR5v5
3k3DLiwMRvqe2IkA1kH0IXNabMtfk4wADPd9eQAThuTfJO9I4/+hpiELBHq+Zslh
UKX6YqzA6XiaPiwosYx2HUHz9qrs3IC/OIl7EjWT3b+WXH0PW0CnAVwxyFNlIT09
7cO/ZKDKA5/bQGsWG9ZKvmrzNrrRH91vTY/dVy2R32A+0XLcvkyxCigeonl+Zrrc
UwjuD4ve2tIqCmK5/XcfWTw8ImGrOWbKuRI9M6hIG9jKk4/ugvHWmjnZEvfPY0rn
EHZDtzMd6uXM9rv24XB0rfC1Kv73HKg56EPwoEiEf/BflQ8pMeMCQ9e0BOnY/uzS
NH5cLk9fCkGXD1TlhmuDINoCgrfUxyTL8FrAjXE2QKyyq9FFEtMG+yxqSkFOCDPj
MzBura63+Z1QM+ptLgOZeuc2yuRFJS+V0t9Hzz4HfrEQ1pepRcs1XmWGMI4KPk/A
e3bkWrF2crWqB6SaZGQZ2zXeBDnLJCrDzvzN/K5k4Pl9DgcZqgP53xSdXqGgAzhW
s7018vqkNJIAe1KSEWh6FVoEKgacV/DUTBnNVWYoJf/lSEL3MadwJvaTUZLSgCVE
sxSCIpVIQV5WFAqJ+c1zsC1hhsBM0LWJrrMYg3hJUgm6vFvPFYf3luVjwDer1ZFh
Pd5XKYF01uZ/RhIamhzMsR0FGKGOysErrz8xFjx7CgOAPYYDKapv2lAGWSa1C33V
PU9rFcrF5poLzrTAfwTB9zI5CafNxSwbw98O0H3CN9Odv0OGvuJKSTV7Nvq1OBon
aRRAxv6u+0UBq2VovmaiG6FeofPIbDROB3g5ynXFvPmLTSPuJ/yyaV9iNBIdxUxO
3OPeBJEE727E/xWvRIsFEgeU2px3P/Wc0piI3H9Llj6KvIiEnGz/ZTi6ltagggO4
wqQhi0aG1MZajBVAAu0lak6bdzu1bzo5bjeCUc7Lac1LFfHYKIirJsM4GbBkVHfb
2y5gAMOspxbEnAunTwQgM+T54PnXT136JdDW0RIZT2tcPv+0X6XtojuEdsBjV+eF
eiJu/owMQHGPvx2p1KhWVJwmHdvnLS0VlAszWYprjQ5eZp6ZN83HWEWDie1MDutM
zT5O7mnSyguL3NFgIgijH6he/W74MfnXZNGI1fS0POQ6cf8ZDeFPb7tI0Gt2GOkY
rdwXIKKK9w2USi1Yt07SF6ATJwH8qMHFZGseHHIBAh5BiIKjeiWqofQ8xAjGoeWd
OyW8rxW2vhZBtKVAty1GSM9pAmMhi4thuh8rf4oh0QCAMOgN/aVE+uKl/8Z/pZyg
MuJ5b9PcFyaOy7AM9JoaRmFWY8HWCpWor5uWror/0+FzaLXPZOYqRNQhuJhThEZw
oWYULhuFPGruEG4TH49zLGQ1ps2PESVfq1CkrVVfcyg3fDhV55cO9VIbNqCu6c5x
1bA+wft+pYPyXjaoU2jdinzqxJN36R3Tu2+iETWDYRmGJ7hVJAqTd7rOG9gVI6jj
r7YA6YXE69SANih++AEAGsKCfFD+2kA5B4SHCdo/WIGBKR2ObYQuotueXjImF7Ge
lj1UXpI2CbJNRXw28mSwgmG0D8ewBBBu8z3dEJpuVE1RVna1oTdHrrQIH4cvbBU0
Qrfj5pYL/gLFLqDZpF5QisyVM6bE3nISJ/Zf+ZDDxR6QBImJzREwZ8X7icjI2p0+
zlTxB+YXKhnOlzk4woL2h3r4NB0oDzH6/V/uoo1KkciLmcGls0yYIFJXV8l8rlmS
Cobn/BH8+6Ie4PIa0EUaBRpNrJ1Ld8rVvEWLirSK7I/glV0Q9DHOE/SJejRDTnKC
g6kkfqRNSXP2wFGXDQCiJiBobxqdHW412+rX7H+YOI0ovzHk6p9dJGsuDlkRm6Yq
Aj5Y6jxJHwsFeyhqoVq/oAMpAunYJTRxc5wEcqQnZ+awkGiIp5NgQsK02swcCEYk
qHDF01K+sxzg7V49bxdBFXm8FM04p1i16mjDVJeyrtTy4NFgF/RP4XxZxe+XbEyN
xYifYExODfOBPF3krXUFkg+wzAA2orHv5G6AlzlEUoSJAuUnX94XyjTkA6mVnNz/
hXlPC++K6JB52YewGITiF6hx3k33GU547bDLwz+6IMPYzaZr6HE9GR0ACwzPFxSG
kyxjCpDiwOVbStIZPP9e0aKdjb4LeI89opsDdCuloUo20qS7/XcDcSQ/4w8I07N5
JHGqguh62VwloA96tms3ou9TjZ5VukOuPqWkm5R6AHKt1FlF2qKBrrFVdsEtZryN
xkEINPB9Zr9JQfvSTZvOi7xpxELghp8N6RutfEKGTuhidGiAorBPa9TfM+B55S5Q
yqS2ktF6MH56PlIx8NwRDr5DXnuMCQWdLEVVWedf6rt83BjxxwH5l96JaFtRfoes
ThtHDbVxW1ZXET/D7Uxx/xieACHOt+6BscC3M7SwkyK4MtVoExNvn3gwfnnyD7M5
bxKGsABkff2fGWMgFjJ7eZxssjkdIEM7GfDhWqA5KL/sscYbmiktiW9oOo5Nn7aD
6XpypzJJcb6awI9VId81eDSYtC9d1QTDTjA6fOTpZ7YeqS376YIUo3OB34H/+5rz
3i/iz8Uq8IH6TEFm4k+ScFzFedgam5FSLCgBa48R/eV3L3HOaciubVJ50gT/Ymqu
hnHNuvT29U7FZ+TaItFI9w7ACarT8UvaSlGIbcWSS5pp7UiH/F6oBzirGu5UpOLc
fVVpVS5MwShZHG/4oKRkca1YGiTn/WaMYM8M8cWyZcK8hoCnlvZEsqOPkK5aR/S2
7W2IOrqPEMa7LOZGJDhnGa0+jhh30NcxNH94LFW7q0r2vdUTupMe0iTnF/blolMd
/5mduOTKfUfhmF/+u6K8kvxy3oGEmm/eu7y19nJWWeRlvPJ39iZCuehC+NlR0gMR
AwGicAIyDTimDhQAicItdN5XrLVjVctw7GTo26xo2DJBqk7/iJGBBdsbPyp8QhDz
JsiTNJkLzTdgwReqhcI6hUh4sOCN9c6Q8bzzw29t4iPADnoHlnK6dyolaELEAwpl
x109fku98N13KkXXYxSx9jesj6S+RiH9+6ObAm/eZVWsKVaEB8MeWeGROSzXipJC
tW5FRPNnV+T32GsXgFbKVNo9udALbO/QI30S5Cd9IaYiu98xB8swEONs3pFzdYWq
xWujYTYV/BpRumnYwvhnLWbgrKdK3Q0oUyObkU6sBqN3W5/6p41zLFcWDXCrhFj/
cUjLUrCYZeBUwVRnOd4ShSZsOb4eOQ2vDoHnQ2fv0RkIgky9Sd2Klmlyn+8MRTzY
TOxBn6Cbu2tF+JGkobXZjLKEikPTY3K+RlVW6ZF2DeXRLMG+epBeUy18m4ZnD5Ek
LJsoaCr+ImN+dNzvFIkg5gbO+NOWrSzFmPpTLNQkDAVz8atnxeFfkqPih5Ld8qhL
6FWxvYFNY8WnCPHNreqOB3cmBjuqsFGA2FB2WZMYHBIP6u/UJBUnMhABGEeTzB8y
OqbKcmIda8Vo8qOB1RpGgZfRTReUvEqgxgzToUDhjkygNWojZv087put3+UeYQY4
DlkvxW4mvEzFt00PF/ZsVfMRWR0E7Y9XmjiXGK57lzlu/6gY+vJA8lMbB/r4NVP7
z+ceUmNp1bzOA4MbWu2oTBu6SkMGf/h5/qj+eu/vmQwhf+FW8+Tj7lfZPHmyi8jK
IMCmk9voVRxekVRzbMxN5k9m2e6/QsTdzBNnExPOAnwLzhKgoYoA26PYfLQtYYDx
yVmy9M7Ou2j+/EyXuZqgLH26I1bAUydT4vrFW9Ief2N+a1IQIu7sMuh759VEZnTg
Lg2JpOR/Zv0oulT8qlGpCKVT5W4NzcIbOcsAruNFlt7LVUFa+B0DVKH6qCDwlK1t
BkURtS1goIdJK5eR+mb++Y+XjWSZnKkAwo2H81PYL/RL8sq51No9JhY55jG+NHsW
uUaBpCjTmYYGBTWK1JePY7utMIaYG/3IR4OkxbaOPP1237IQXuqWgHUW2JrNTpic
iZe8F08csOCRNPNFwVR/DYk1aDGlBkZSMMGftYyAaOfDi4e5DCCiEUmFMtCJkzXF
Rp5Pp2Mis3+hmHcZxEy8sDK+Ov0FuUPccYDLm/s4Mo3RLTKZzKthBuU6/zG0RooE
LKDkJq1Fd7cSlWTYGUTa1/+CfadkyQwWeev5CBiWD1XLaMwjfA3blLBFwDPdhYbL
df18UH3WMSFeJnUkjnbTTvSThxPW52DfjOMKDjUAvitA4fvVJNr1KGOoQEOj54qj
C7nn5jjodGLm7sGSkt5f2lAJ8r6WI5dVlEeK8Ri6I1rJbJnQ3YDaLZWNfZxwR0uA
Y0RhVGFLTmUhtg/e2h9YZwdkogZZHknucHQ5ZNEhyqYsjB/jWZhefX5sU8f19y9/
4go0g8c0CqZ+oZyjIswtkTGJvg8MnbDiE4ak/77ZBgJ4LPb7N/5aAm3VlwAL9hhk
2hu/qwSzjUA28sCqH1if0xm3lgOIJnd0k4ixzUzlhmgFQZAoXJxHHkQDTd0AXNP0
6H3TX5I8JUVsMAre00CFjboQHF/6x9hqy/DTWgdJngGe6QUELr8xJBoqJvSFTf3K
s50OLB3hv4CLwtqxkCTrWOBabzSl2Ho/ojD9BlNe2BjHlhFFp26QyB6wEU9582nu
WWRazCgw7j9YcW8pE3mUyBwTtedeJF15trEku1yhtDqMkGIJeig4IN8Qz3cIafiH
J10mPFeUTXb5k7Z3jomtOAyC1V1LobRyTYqbHbjm3vBzg7uYPTudkh/ScmTajvbi
pZKhGhKqXBCehVOP69jyhVJNeK5isJs62qR2/tsstkUbvPzkC3BtoKXdqhulYzZm
pDNayuA9u8fid0GkOFzkTzlvtKFtXeLKOobuxwHSqtyYqqLtp1QU6+/iEGo4Z3ro
0T7aoN+XCUmT/dvyRHQ/GZx4Nyga7UwLu/5u32cxQ8XSweOQow3U7TFbvQAPatvm
knehl6yfud10VhPUtjjWBufR9Pcs7DugCrDdEFsqpH47n4UeIYjr7WEWdItu6KOg
oPl0dDqcqA4V8CkavBbpGMjfqBdQyFCPe2LUQ5OK8btzRIWwJbab88Gm2+SYnKl7
e/Ej5AlPli0lmbxkfFb7DC4Uqq+TtSFrnv8h2hRVO84ke+V4YwEVk9IoRsxbEx8n
rqmnVhFwzPiCELBl3DYOgoPNaa0yZeFYJoFWS79cgBDTP/wddXNt6QKXIBlB2BHR
FiEqepTx/EDJUBlZ2CuWNWqbI5bFyz1LAV6feizEJAQPobQh2x19fDPDy88po7q3
BufWp6CWOIxUolSX8hCIiIoo+GBAzgw2t4eVknncxAoAU/IATw0EIpA0RVqYJycA
7n+uhT6yyOxQHg95T7hg3MyEEo885jMUSCuXyh3pB5guAKkbAdKdcJKQU1r9QVnR
bGcMzWfw5/F5A7AyfPwj0Fwrp2tWwv8nOdUQN/Wkz9Hg98xWs30UpMAP/mnxcqmY
kng2VxDK88GDlcDgpOo45md5vNWdeOHCsrmFvsCYaakxZV7qy360Y/FVp43keZUj
a+Hxtkje9CYv3hK/39THHTMuHh7QEKXd7n5EfVumvx4onjRWurM/8fFsl/SsQFKI
L9qoZG5lMqUJW6lRPMkUo/uwxQ5njXYWEs4vhyyV8mCsigIlI1w0Bjt8QDFqki9N
uinxLyjZdRgy6mAi7XsJNgNCTUSCDWytuLiWbp7IT4wemmB9eoUYMYJmSqFSPDSk
VRDCBa783wWQdTRP84+vMutzZzI+1052s2xYxfP4mYncGfOABjSh2Nn0dYy6Ui0A
6ypgYCIloqgkwen/JhmImYigUhJYNkAg5wdQs9V5aLEKt6ITJ3TBmN4KOhoqcihe
VB8+ln1tzhx/nuS37vCrWnSnhe7nevxzkUiZEZ4UBvETFRNMqRLBdoCItQmYI73L
A7LoA68SmitNCIdBhlu5xvt3o2mifB4BzV+4g6NDLEqPWo56zu89xnqBypyamOaz
3TdhimnGgD28C6/Mr8YZE23w+GO8SqI+oQvHvTzC6GjnxFmm4fDWf5ui4pSgiN7M
lmPIQm+c1ZmzGvJo3M/exXhUkncWY4M5fiyw0kU2s6zNOVpaLZ+dSPyZHfqUrIgP
71CEOKvAOoYvWd7M6QMHZ+Zh8Qynafcgn3N8mcK2UD3UYgjRPhhQD/VJL8NtKMMS
TVVsIC4oK8+6kGpwL0s6A4MzSCLEtH9o7Rod8rYbQL0Phag9RaVs7eHzC8eVRT/g
5SFGvGyXa0I1vzRQ3L5X/VssRUaBqay3Tvs/8nn4VPjIpLcB7UNcPfCX9AJuMTX/
O2r1xHa5QuPmyaqqC7d6JPgoHjuS1FNsA7/2bTez6ZQyXdwAmQM96ZFMn53jqHVM
+N/AtR7XBCr+rYKmm7I4VPIqC9my69QKv4UmGTMq9mSLJCRbd/Zz61ITtLh2TAQY
d55c5Kix7bdg9C1Y+9lZ0irVdWotasmhDLnUHk7dP/u2PlE2hj9SEF9Erpf0QkPP
0+kfzcLZjJnS1qT6jK5wM6uBE60keyX47GZGFmTGD0/JmIFNYMcZQ+hrUC0A/RXP
+D9CQD1nQdEtu8epa/nDlQzj+UKusALKq/Oq1o0zXbBlqUmdM//uccU0yXgfNH+e
5bIHPYeMBf3VX4CJG0YBbWMXv8IKoCcC32IcIAcMl68CYZkl8weJCP3BX8upovb5
f79aeZupDWDAuXxkzNpieBDRZ6hhlQH1qMR0EqhDWJLuLlOwXESXTLmNEj508exy
0Sw3FyJhNhlHmwsD8l0fY7X/J1xZkHNRFbE3QWeIIJyKDXPz9IQfb8DtcOaiWRxE
UbnnoQYGgYBLWD/H6tRkGB6HW8olWfXvnpN6jYFShKdjJVoMmiP0U05fUO9yaImC
Y49NvORdvsifMvT2bEkqaiAMIm9GRFXNi4LLAfX9H8J36qzn8zlAMJ1x28G9id/E
kQCcl1XI2BukWtT912o7me39L3BzKeuv4naYbdKw6fg4GGmrfmvXi9KNxffLGQ58
JdREsdJ+3KZgVVEasgjwMynjpmftzNbHrLa8rt6NE4DdTSz1IuAUeqFLSabsXBC1
Np7lpof+O9lkhwpXLqZThjnpMnuAlA0OZFl5cLF8nGBDHf4Wv4dCHB1goQqY7f41
jtMwA7zMXWUddrlk8qGPGL7ztv/cm3WYrOBKh4YzYFC9CgAfe3iPENlvl0kU6wcf
OY47F8egJimwOV+oXyGuFJ9uPE3Nhscut8Xa1S5ShPosi0Vt96OsJxHQF52FFEhx
97BbYKaQr+J6BFy00RjqvRYJSRLRO0ajo1VT64BNZ4T5sL65Q4aA0RCGTjq+3/k0
XlVZCzHgY7H8D2A2fseMKflodmUxgOXoYdPpQ++h/0QnCs5JxAi4VUomBcWswoSj
kQjLU3DFq898njsnveo2Wep+kATTl4UEq7dOzxEAfa5frjURqKNwiHUfvEgbN+r/
J7D48Taq8kkIxHZ1SwuTYwhG8zrwooN38/UNzBGTyjKEI2A0dZe2xZUVNDgUjP6s
RSaZqDcep95jcc1bRGrnCZY4xcRjqjeGKkLDQ02F1XN0EhLLVwjtNIW/C7KQek5u
yZp9yUo5A6s/nYnt5T1IqxobupAOgVz3AVzEjdqPLtEG4YDXm2gWAEDo5PtZCC/z
pKemLEsSaE1eTerQnuEcaonaIOciBMLg9jk0HeK7y9ngsiq5sjlJo0OqrPUtm9a/
l65ZO+udN+CRUfTIXveWca4pVVSEkfzYbr6D8xa2VtQEV2JDjDxv3H5M/hDWg6wA
v4/+S81UaRe3bS7/kDnwYbtFJ52b0BzGLDu+YnrBHxC54Cqd4b7Qr+8LMs+G9+co
aIfe0kXfet20PX0ZQpzU6VzNphC14M5HpgEZO4Zk7xT+GGoCtx8nx853pOYlYD+/
P+o3D7QdLOHR5bLInUEgXimnjaDOSmyEXuTJ0qaVZhxrZklrZ9l7+0p37l8cf3py
JFIGG2M2vJsmsxtvpbs4njVQur2HxivuHTylGpLvcRoxMwut3XcavDka1wTHYzyv
OEs0qn8S56KiJx79NB2ErLqyJ2TaperR/yAQ4ZX73axC2P4GuaVBthVg5Ugbc/Pa
1/YwEb5IpeYkNyVuJ8t3plF5vKvwj0JdEVtbeOIju2ienEgoCuL++ah7c/dDx2/1
vRBKNDW16ESc9Z48vahG6/w4M4yeRI0bdB3ZFXZlGEV/Xc6qw4Km9pWooK5bDIWI
Foo3Fjqzcac3m3ePN+hv7DefwJXFwm2i1MhWYS1O0TSmSVU3mFEowYq4gZFahUxM
njLVMOpuz/+CBoGxCENLoTJBfNT6zt8TqAWgob5FKsTiNazkrDh1mHtbkOdEAqB2
Y6+zvZxFSY1Rpk93svElwgeokjLtgUCaNQOr025Vv9HbOKPPQgIe6SFVUfpcB9Y6
0xSaYBZDgG4Xvlc3Vpk1oI23fo+F/ZAJ8EXTneEQLZto4oitNbhgunCINAp79Cdn
HHkCEewEMqa5ULzDtt243tnyPVZmWtVExzqTkGnCOokpONPoRffjkTOAbzUwDLig
pkMNKkDz+NjeOR/BefKlScVp/3hX8qoZ3vEkDAIOIjNfo/JCYxn7SuDsZqgvW6UD
k7opfWUHmynssDZw74Bzs4XBPzOekoNZ4pMYTr0pTTxCF3fg/ye98/2HF7xpIayC
jEyMz7+4gpofKU6tQP/3zoYWxJD7XGXABmfoaeT2LtsQKLO5awWki/rUzqYIsNfG
L4/S/qUUjhwTQA35+ekOWg0KnQesBL/sQwirhxW0OY8WrBYogDjDnIUWm1Q2LAoe
bzPZm1gZycNQgSyGp5qiBJzHivXMTXROxzOqM+/ky2iA8bxjrrmZwuOI6RpCP9GT
EkIdb4vglZutxzXP7IwowMoZfZzJ2M6PEfZZOrVtLuBl0oIs5Og6WDZoGT2ZQ2+/
nutLvnXywyomXNnyNpTdcJV3/VXDqhpJcpI+BxbRANULMmB2f83qxxAkxEXu+8hK
HeWr4G+guqzeDIwenZXc4BAGmNMFx10aZbXFAVSD0Erq/UrRfupgcfoNJy2N+KB+
LG4+rQUVHWtNKARlm+H0aUha+45+QX54MmMxcsy7P4G5P8E4O5XuSR8ii+buYfC1
kvuJoiTYriPZi4jRLX+iVBIOgTfJDtIgY+SGUAHyWUZZ2iy1LQ+YTvCQTUC3y+qv
mF/QzAF3rwXOv6OzVBi5gBjUa4YhU2JDF9gNrTyVEs/Nuo1JYHx7F1UdAHld/5Bx
j4jf+MLp2q32itUxwqvD9YcOcSN2AwPuqE5kmINyj9DMnHGklA3Z3j76213Iu5Vk
UFMwFp1uQxd3K8hTqTpnMEAaNLPxeccg0EOIqPX5UeTiNnuHosBepDEYxj+jKr9F
+++rqql1h1TOaM3EZ5IHu1OOndLlmTb3HRIIMoZd+OWTWdIqY4xqHrdsfz/a5kH6
S2r3r0g48LxPg37i41bFAcU3EO8O2F2hcCNgUahsesmb+UO4yD+GpnE+DHXk4z3/
xVUzmOGd+3Uly4gApcZ3oSDfqPXaeidYhhvbWqgqCH7cOpLmClevt03RfKMJq8U6
+sHzu/GbQIr53c0S005UCtht0GwqM8eDSKhJWtSDGjGSEyceOFYxKK4g6FN2rrKN
ol67Kl81lXv6/pTrZ0tTxQwDIEFEa5/jEuV+Hos2BYA0dgbyuB+rS5PLszmcXp/f
3DpqFOWUFJsA+0Jb66EsYA47Ds6By59ItitCHCofykgFc+jbt88lWdzFSKk1cUWe
FdMvoaDHUEeE7wXkEEV6ku9pbM/3DAZrFO5Z5tghn5gN1E9M5Bk2LchtlFzBAt41
ISD9SHPPpSXhcx/9Y0ThttNtegQMbTKozYdrkPfHDOADV1pkDesbONplCM/ivKdn
oLOn6EDYDxEicpalCSvpGiqvmFnzIPAlvHmyUlqk2zO0FY70DuXW3uwKAczPvluC
1KHRXk83XRipJfUxulO52Aj3WsF62G3T1YC4dcO5cViipMKErvp17Znd1zmUi+rc
AgFKe+kZZRCZkqXQIKiCzywh3fPicnRszY1E08X1bwQfoArOi/LncjtpwMpa/ci7
Uw5zPoOdBUYhGLcRSX5rrbpLP6kjq5aftxnvNEI2vg590buietIZ4ngV/P/eps37
/e0rCeAsifA9Hnd+ClptQXedurvwybRfRYtizRCdYsRM+RPhIayMoH17Zkh8LdMl
xO75WHIjAyzVEMBzbrvwAVJIBuehEvTBbaThUm43OiQJs45tyiHNtCPPnyNtB4ga
2t1NC6gxsDTi9arzX7R5fIk0KaIZRewjSZ55W4kZtgEAB0orwVS4LptKuR5ydN9v
+FX/zwlG0UfhhVcPmZyr0U7+7gcnbxb6flD0gMSPjJL7dT3c5lSYU+KzFWFJCzdG
n7f0PGfN90eWDRUVpc4hRt2NRrkOUBrdNwCNDepnYEHQZ/QwPue8CSaCSsbmYlyJ
0Cq6Hh1gWey4HVSYkhcuIhZwD5MzqbNtm9EfTQwRtdBlhFYFy+GvdX+ZryT5uRYG
jM11H/1/HBa+DL+FE/3FSZ1IUFvJGBEmf1jUpAcobHSOmQD/YVk7sHlOlgQ/opy7
JCAyNpuvt3NnKZbvvsFYLJ5j/4w0PXVRIbjr7rOhrQBk6ABU/wKYres4QdraPIN2
OeGfedI8Z8DfEpoRO+j0thA/24+9gTDlXCalPJtr3o1nqSLYpBqUz+t1GQEuRY6X
eIJtRiPwc323br1e1CpkBo2SEaNDGIy1HwBtSBHTit1i0RgnWniLdCVfRwOm1bff
aHE1ITow/VyOHhqr76u06tzvCFECqN6E/xvdThimkIN7g9cBWdiQlJlLUQBWlBk4
6w9z04tNnYbSvupGC5jwp8mseyKgClWbFntcCNddEyGhh09V6RE+ffhfap1Xq8+w
WuZPHhy6zTfAg/jjhBBf7rNxZuGX17WHqNkhZRzGkyp/0Ge4g9aBqeMpw4TmC05U
nuslbx/9ctL09POAzbJFXUmJDnif15E3H8rooZLIwf/6vKPgPH3pQjFmh2zBG1IF
TZKvtVnZauDEh9JcuWdnYvlFwPtWMgnO/ZgqCv9m4FSkR8Ry/TpcWwkZ6YRReO+N
FnB5pwo780Svml+mmJHRiDwQAVIsHBfcE2H9/pF/+LkQoKdvgjdPtiNZi0t/K6dp
t5G09rkERt489a2RDOh3qk6DUUKYaDqKs/J1L/tW4/Agv93F9Wk4YwJPRlsx3imv
F9mX7MPla1/SPQqOTZAI2nbSuZ5chwC+rwZEcXwDMKmtZfUuJkjuCvAUtykwvPXR
iSZ8n6ZszlcNPYDQRp87QIz6sK2SFJYPvvofFK1H3gkW0exDT02uqnOamwcr452W
gwX59Dmk1fVUbyNYMA69sr37PG6NrJXUSCNPtetLUFEWT8CqQSAxbm6+7IjTcEKJ
IBgG292WubIKoC3SCIWStltMr+5hNpeLa5IBLxcFwzDp7875ACDklMJWDrUh4fof
HHM2fwIiKtI/SOte1KnT2ta3VT13b7aNO25HFPvjdvxlgj1ch8++VSSimKIKfLfD
bwSfDseAchyBe7yz54i83QxG+YCH6ymKVAWiCrnGMTfkflDqc8vagT0Vye0p9/cf
c73CvweszMbpfoD7rhnF1j41wmNAHzUvJgSYJm7OuFYoIc81HsYpFVMhpw2LKdne
2WkbKsqlOpUb8jTrDYM3tjOjHasxrunb7rcSqLC0ll85PISUOH/H7cXCRI0js5ij
SJEWVUban/Z0WMCvMIPBYU8AQ73zkrkRXJ2P//T3wq8Cy+BM5Mi8rHgOKAnJza8C
vu2/i4B6S+a6Mvf3a/Q+Tr2zBh4pZW2Z3HeCiRuw3Ge9z0cSYhuFQkppkHto+lZ2
Tz93l93oWiNGE6bMmvpEkeD+f4jiCX+VCx8CAQ1nwoQSpxSQB/V0Rb//svUovcaC
tDL04n/1Ev/2f139098YUgBf5kkllAWHAD+GTZARO+8RzroUD2svrIVhkNus7hXa
VLwXcpRq6J2cZgwFr9u7Diz3UwV3FA1fPNVW0oQpH9mpoYMpya8g+O5LuWDzCa7f
bKHIYJObLzRvGxxk558QlW1WJnp37yalo6Q+uGp+LnYvewXT03jyAkyucPgxwJlv
/ZMtrbzByst7ESn3NqxJMknLmQIKkn1hM+iI+oeh9E1Rlb2TT46t6BLpOh9Ovkii
kVVdU0YIy+E8u2FskBM8eBUZx8HlaAkbIFV4O7vvx6SyFMABGOsrxNi4zUjThStg
FnoPNGxOX+Y++B4EPp2ZeZYZsaQKf/+1A9GJTIiZN5sjdR724lJRJ3fwwvGIoK0g
VM3eD2/GVAVXS+AaoPvaArWjKeidcy11Alj5xsW6ykDYIyTrnJnr5sV1MvowK+I2
Kuz6IzR9bi7xx6CJKFpIPuL9piZBt8CuIYsTpJpiCd9ZeZYexizBRzs9sb5ZRELY
M1hN/fr1Q5tSkqgzOQkv1+TUdwU3E4KYGkdRi0E1MGF453gbv5R1hDD0vJcZUNFp
e4kP5LZILjkjf5PLCURFzB8CuFu+oBtfItDAgNw/4og03mA/jAXD13bY3lAAuc8o
T1bDRt5dSsXppdwMVTo1X7zVw4pD2moYy8X0bQj2UJfc73worjGvWGFcv1e/YZOP
T8Fj4NWgHXfBWM5bTCz3QAO2xRPigu1+Z984KLgTbWWsiGiX9KEk9KX/uOozozyq
ow5eBXWQnLmbzlMwyo1dEPSNg1ulyzKQ09WjN4W47NtIBqFuxMk91J+PRH8juDi8
IuFC9BsqbYx5BvepSahDVr5BExKefbbjYqM91XPT1mk/Hn4nExFK0Im0UYBr3uLU
gXg2EmQVGnO+fP7cBgrJnSgMZU4fYMCewoZMIauZ1Tdm2+1tg9FBctIifkf+Vaip
lSRMWgX/ef2drb7eIqwG0b+qHiyFjgF2AkxG9uCi6go7dQ3nHZDYL9BREF/3XHTf
Zv15oM1//EWREBMq18A7h4/0GxWDy6iUH1LAcXA9FqtcFGFcVKPfZGIozrJntcwH
4gGMFJZU1/96XPlqyxfwlyp8L5cOO9yqnXZWL3p9zwpY8br0gyl7dtWoVGKQfkLi
gxYBmM7m1ewWtL/n1b+WPjhCuTJxtXWj+Cq0DnKsETxpFACErbvAvWl6DEMw8S6f
OmHF1k0DQm9gs3VCRq3N+amRmbluijpgYueV7JAyHU3S5vP3mqSNSkDXAqrpsHAf
OMLpRIZI+AzAwoj0tG3Nn15hZX1xL7CWhX1mcR10HJDGwewyhdsiHNuWz7hrZ1rv
qUMsjVKvrdsIFjYdbKtJwLqGbz8agq79BD5E2me5SMgVar3Kh+vqsoxs8YLEBBxP
LcdhfKkoRRsDfe3cEfyEqJb6aq4eU7yxlQuG2lBVhvVwEDNaVYog0hygy2v5s+rK
lWGLvk8bejJRgm1LK2dZWxCy+JLEFAGtLm2xmRU5B06XRyff0pQ28ivqDKA5r2wa
Y5IVjWCiV+Rc7JHSqyumCV0iagMvQ7q2iR/ZSiBwx7FffUc9vM/A4fTmHtOfvaB+
FkJUwLUJppDeiLUCKYA/UwzrP0GXEomnzSEqWG1hQfsx/haUA9vdX7QxZKd4fGOV
jOQzpjwqCVlNt+JIb364FaXjHn/C8fI51VzjuUbgIH04BVNMpeWCLEnfes2ok49z
FEd6TC/p4528WSq6Y7HyZ5BjKMHJkD7Etx7T3jrVQBnetOj+yiXoVgT5GVviguj5
7GY5sTRgWYshrWqbQ97O6VqKt7uv86zfTmeHUmpHlwA+ZIMY1n8OQZe1FdJuodLT
fZ/E1eHC4TkhagsYG0xfmbJXZ7totL2mnLxKE9VRjTZVJJw1hGnnaGL1/3AHQm5t
ZaI3XxgZ2YJdk5H2fAObl4Ge/A5RVOOTq1HlqLC+Do6MKKlM80na1HbnNT/GUY6r
meS2wnFOZ3ckT+zsE/6qaDXdq6V4fHXWGUfkKSqOFb7yLlvhC5TiD6hYJF8jK3eg
gSanLMmxKi2dyNKeWDKB7tfZ4bXf57xlAuyzs/x77g8J5eyRp5ftvmN5DGpZnlzs
8iYVgk+wdKQy+V3aLq2Ms76QP9aKexfUXNEQbJFNBu41jdOnW7PU0P7ZyvRIN/wz
xV+lz6DftvLGyaoO5sw0troTedYmH35Bx5BNZJ0WSaydLiIdf/4WRHnjGcnYwJY+
z8h2vdL8W8vGxJkgmaszv2xss7gA+/OJ/OmslJ7h6gs/0e7r3l97xeWmErJTNe7U
sRZJ6R7IIWOEPh/KdHIM4X2KsLI7lSg5v7Ud1yH3sVr8zgDMZW2I3oIrw6XUD7Z9
ouyry8jwJWfxI4NUfXzvCQNSo5KLVIry67qObs8pU2rH4gxxrRpe6mTl7ZnZy9L3
qKuovx4ZvnConK2HHhMaiG1siI83qox9zT7UWRiJ5yvDV645663p30kL6AKi3B3p
jp6DjqGUUXkOFVjrhEDepGKlHDj1ar5qK2jY30yCkMw4KBJjS8PUKQTXpRYHalJj
UhURf6ZXApXTFapcI5M8SSBEvWO/eZMOOdffzqH67HI7kCRo2yF4R4r+51E9h8zu
JMhvOSbRKQ6kxoJFSSKCAEOotwse3WrJw1R4/a5Jxu3LlIHuCCsIQAMuvchRzT9K
3mhqhotCkg6L6CXwocvJ+sCicvPPLsebEliYUDhca22O2OZz5GR1Nppzbm/WVqbB
D+Se9OnKjS68wXv/RG4aDZqR13xwh7Tffgz8KzqVy1s0x3kkU5E7iI3fn8CcMK5K
MNqUu0YTKP5GacQdzRNKv1HsanpOe9BVY1Yyx+suv/J8bKc3AnxaFSNXAhYUp7Pg
oJ5R5tp/4Yr8Qlj4TETWHYO0xU/tY9CPMl4EHB0sJVNMDaHOhhurXxltbLxmEN66
STOIEfQe6bgOv34qcNf/frt14uznoqwf1GTaWI3qid3I374MUeH3M3BcRAIIkJr3
r70LR+0AEK0lD+sbp70eOmSYo1ohr2cuZ3wK1QewHQQF9LmkSVG4+V3/mO6JrDSe
GduK6yWfzZ30NP/2hM5tqvSdm5EJC2VGEQta2Y6nu3GDe1qSeTU1ABxrDr+YmPWL
Xiqa29RJ/9OlMKTjKQnVuXWPRLYAQqdiGx2X4bdBSkJrGilguSHm3Sr9bSkmYDzB
vQfnvvG/GTHZcbjH/IWcU4W0UaWdOCrzP2QOzEXRD+cit7L/QTCyrMTZoVM2luug
qkyvZ8K0mgx7rWBfVhkbM3DmytDJd7PaJpfbkNcrMAXLyAqubAZkXvMBN5qAm8do
whc2a0J/V/Ck0WK5n53iYgGCahI60icMA8KbTaXMcxQDle5a3pCHhWOrS28oxbg7
KRiFIvM/t8F8huBFjcEvPfGacriGCwmsYwmD8/2MFudxPDR0MQ1ISw4uZnH5smFU
DMCAOtksIG34HIKjPbmhG5jtME6IzcgwZGaB73AqyjCUbn3L6DWfcqhoV0HYH0Qo
JU1Znw+i3p1P4Pi6Iz+2JK1DEKHHJ6C2JpRN84PCRg500xEa3kvFrtRhnKdkc5FB
lQ7MjqeEXKBp6sBZYy2F+kucbV4XKpvlEp6r9UAjeuSWbPGiK9ufzumxsdDZ7dXJ
YFBzv/fRaFACp8BZyxeATjVExW5NABF5MzHgmdNokRonCcv5An8LUUze+gZaSiHm
OqkolMwYXZLap2WHxIXBJJetsOqcaBASTIFVPJqgUosW8No4zwLkyYvpF571y2WQ
KFojYwjknh/ddEJpAycMDr5gcRv+iJGmQ42nm8giyXeWmNQSCCg0frCsnMZw1juQ
J2Nt2zwVoFIjPQDGTNy4N0z4dNFMeO2tnSte9fEGOVTvoOUgBFciNF8Z4tCfEAxv
Wi75IY6jz5+PCXIAr8vng6AJAFYe2ZlH80qxVTRNzb96lM9n6LJxhKthOtBaFcoU
W6i2pTuiqFICIg41Xzjshyv80ZeTjF06lSa3eL3Uzt0j2VH0pAue5XWK5e6iIwS2
dLKzTF/ZxISD2p+Hcky6slRciOaf3N4+t2CdXTy0tQ9By8TW6W0gTdOicTJyTkv4
+0tm9koNypHypRlIdXGnrj5WngdhUINWB23Fk5lnH08V6uwonxo4PGk/EggZGhAg
BJevmbtnl77m5uNHl3Tl2410EkWtoQAq9mLV0Z6+THejTzTnM5HiLNwChjN6eUNP
1uBWKiTQxi6FIRkAoI/eB5e4uWVyfKvWZrofP4KN2NjyG84UqrASNvVPbDAi9/8T
YA1Sx+efspoO9pPIPoQAyVAkgRW1R7YoxIHwx3aaHKMw/fnq/1K73z3S8eYJpADZ
zpx2fPfIUTM3Xt9Su1By/malwqFvWYjYqera5PtNqYNlElsclVC5V+anMM5qIqA/
9SsGzecJWasinKZicc9sgsSe6ac2uoVYjJcjIMX6JyTgJQ6Z/JauBzhNsBQ0KJ/u
RtMX6yQosNKky5X/zG3CeSkvSlGy9eSiH85sD57bFMH7tMm0x2P5K8ctQmXaQmKi
HtPMxfqWG67XQVoB8VL+QBjhQMZLCAeJW+0+gU9S91Ddfw+zv1acbJ60FiWfARmv
Flkwfny1t2zq66et1uU5aZ49oWtfbyfakGaZMdXvcAkfgIEBzxUBB66aKaiHj52I
1MGoUlSyAm5mCY2pfEUR/S4kL/ZYXtXlgD/s8QGvOhnSjwYN6xJm0BCU/yogdqf8
ZHfeaFYWrGU14Y2HvxGTO/XmJ1QzHd5CDEMpMhyoVjHgEqY16qDsdFfVYLrh/Aay
TAv9Q+ARnepfRoBsK8ymlijuVh1en7b21VpVPvhy4ecjfO0sQJfEYwDzgYQoZyma
mzOWbdX2/C3suzO/m+RRWm4Q+kcbInOhx6cdHV32GIlXZs6M/0OLciOsnwe7SANm
+FPZbt+5FoSiVH1wx9snaikWVjwpCMerJMdAUwjHA6Q6kWNiW/akZTEQxPoaRlrZ
kE9bFUuSDMR6TuLlupc3dU7MSFOmSHqzOQuvq6/RLCE18UVMj63veOVTsEeEAQJS
B96rFZmttS6Mu4TQm2fyLXVP0PuCaZFYv9jBh3tIB84gelo/BuFFBiyQKpMFYFYd
LYm/+osPPAkDdltvcOIocZPBJlAwEzmBJTN0SkMcbCPGUioeW4S5T4nYDaT21I4B
kh/hilxDOUFASqt0J0TOst8fs+ea04Cp1VwZisXrsT1brLaNTEWdchphPrXGxuFC
D2eUJ+55/npCo8RhQGDahYkmGWm6T01uFf4WYk+Z5EEuTdJd48hbYk0dF6Yu1Lp1
hGjojpOfKMR1TbE5xjyZ/ILIH+OKaJWVbiis81Q5t6p1cmgg2blIvvwo4x2pn5Og
1yUjZtUWS7+ycONZlLT2rpb0KrMsA4i6dwGXreM2X5rjLlTNS7xbeiLeeRO5zXYu
e664WDvoTK5bBnu6+kvWO+aGCIS0O+t+SBrnPwmwNHsWZZWA1BzEHV86gnH98Sv7
+sx2nYtFCQhejGSLJjE3FH4MpPG/v2mAZbD+szFuTDJ6DeR5SEo6pvg/1/I5FYKH
4VnGWsGsRc+dmpmRE1zAEvWuGNQWV0jWKDTmbSgykDiM1J78a0BsS/sZaFy8gT1s
qy2AasToVwsuVaDaxA2e5kqG2Ye4lseUF83LhgkKogF+NMREhq94ampN5qWxa8cq
URMOyEdSAs40szJ4FDHJBF5PyAuslTPnf3YG09aYLFdHxCVyk6vXguP1m6OsN6hG
Wu0JozSDg6onKCQOijy7xuw0yxqBDL01nNqMBpm1CRV1eDtghG4hEh8DDH3SVOD6
Hc2bHf0mylw/KpmOVPM/4vU0d45yvAzeQSu2CNF/QHJ9Wua5wtUYC5XiLeUnJ8Ar
p/vwKnJN0uf0t2IXdmDZQL5nWetFhQuuzFeKoB1gxOfDLYbkpSOPzMpsxKDIw+U1
tqsCZI2+kP5bKpccn+GS95PnqinuwX0I2Zyj0SW2KvV4CF3460Zy8WsOADiyn7Yz
8eyyg3BCn9FnTl39xUg1+T9US/Cqb5NZHmMDjQMHMtPlbLlsdW4Bjtinc6i1SOE0
MHlupJ/mv957pLNMp5Q+UXdkxIoy5+qRRmsbXR75dUDsmiZBEn9h72dq/7x1O54B
/p81vM+QSQIJOdHOVPVlwYURCsyIEsccfrypZFPx5NzfrIgrJE1c0whAa541jdLH
Ht8lVHbApA/dQCqkp8M8Al2RiZZ+2+o/CkZVPNcdZOIEaj68n6eVuma3b01S/cNV
DasgBxiGf8wcLudpormNQjQAf7b3atkBL88BsrPFV22uKzQSKZoxIYoVA9aQK9//
eLNWd2DYf6HEWkOKRhgEv5HSomh7TZOS+k4ECv/+rNsi6jW9xi0WdujzCsN8ifLb
BlyIE2UdCprwRDFNbuUWr/88wHsFH90YSTMScbzv68JE/2llpCPi9MGOHagWhjAx
B01Fp0zq671suwx1I+vkr6OGyg/5CFd6AgMWMSpjwpkEENMJ2eaYStWzZKBvEBVA
RvBKv8t2zu+OQ2u2A4JM893EQFCkBlJQwWCNzug1rVvxctbOh4+2CyMCRrJ4a2BI
eNTTEulZoxuy7TosuoQh5y3f4IxlGc3xRKLz0dR6I/kq0H++l+x8sb/aAl03rjrj
szlehRRFq/3BtMz4VPtb7aC6JZebY9z2NxvNkei70Ca0K/SBZnnSMrrI1rJ1wklr
WN9zi9uy4QmakyVUbAzIJ9etH1y/kQ3jzPy3RpUZpXHtEneYVqoKCnCP/gDNStij
Wi3mOYSPg+Nj6TsQp3ajI0HVLwxN2WFky1zSTqpDt88p5CK9FNpM5VtKjhA7kndF
ZadzIea3ix/ywBFk+mRHtCgVNhJz4YYHwFzHXB416cwH+FUc5VANuN/HFqw1woAJ
xkLhsnVmJpmfOXTbOL5kkXP0iAw0H6f2TLXAlf8tVXsMkF6iW1p002aFHyQ6oePO
xIhQFSLJC0gOLz1fYN46aKAcDpreMKTYr7C62v+fnVd/JG/YsfTBBA4EdSFsD1cK
/4y0omxxRJxQG6xCoPmhNNdTZeAZvk6a4Pn6VpiU5waFfFtAsua5EdV+1uOH9vlZ
jqr78ZWFYG9P7iECUGrNmFno5C8qkaNNZSCJw6PDm+Ck/944LqUfhsmp0zYHg/1I
yV4BIwFG3fnvnWAaS4s7TEgdQAHdBsNbzvZbtxDV30tkyEkUZNCjdU0b8VqAdaIZ
ef/l6pIof3qpfCr4UL1BnYzsNlHYYXKlh21EgzqUBtemDeWk2CtqCPT5oHh/iNzf
9lpV42vkln145uLGVOsWSUwSRewb7NnEcGzAClGybBaihPdTlsOLxjfGR/bJ2poT
1rkwZ54oEgSLWwh8m03BK3uFtuW3CutTq6ABdxDsqY9T8GHoYHEjOxaKT07iaenp
/JNAKLdDYTN52ISpSXvgWxY5fPXO9Ch656VU7OWp1xbXgigia1KQ2XNzbYcbDElp
WCV8J4mfflJuRlkf6Kh5GvHvv1nVBDoqHaYTzfTQaYmVyb/WfC9hgb0RtmJUmUmH
S7euzRmCcJ2yGenbPW5tQpcP5zuba6/Bo7D2Ek8KBzk9M3nJhirQ2sgSDGMybtWS
lP7nkb2arhAhFReMlpctHP/GyHRB0qZ1VxNqgXEa6VdujqnxfHzgJ2+9TG3bIUps
U+wWTyRniLf0Hd/ntnDap6394jSsQ03rySKN/QJfTcPywqDtONAJqiiDArUkYM+X
BOtaO3ys/mIcdK835v2a11cPpGug7jreX94T0i+YCr/RFa7U/Kq+xkpl7oX4MCln
JZ8hBeP4QmcIuM6Zssh4jY9jp2q/DXLBCxzGwEyqOTccB3WE0HoBjnC0TjTgfI/m
OamlaQSHjDmVK2cdtL5gJigBIhVK+GciunAZOaSdb9gxh/vysDf9I+AUsIe0mRna
pf6NZUaOYMpRexAIaAPHjr94mas83K+6TN4ZYeTX6kyDb18nzDd14jcIQF2Q1CGE
4eFYhbTgyKisOdOb4lrnYx2xH+oBo5ZBHcla/R9/uoIkdZXrH5VLEcfs1Q5pVqMl
fCsqx/31CwycHGOYsOSqQOnzW4Tx66MO+5tj3bsVxVhA4Mq311cyOSCb8JcPsPPG
VPDGppSK8Tp91HSW7o6ww3ySa3BnXyWy9YOLGcvsc0uSBnuieI/tYXbB4lK15XhT
zayqDf3v9rdq98kq9/1iUAcOpKxAT/zaP0385yKHY9eJQXCh+mP6Bk3F1pATH841
YzNKkC9OvYi6LvtuhVFOpvHyr0cD7o44M8HXdvF1zxHNM/mraufhh+QWdwygYHSH
5dDdPnB6FVc/fWUTg0O0usIEa5Da9bMVr4NT3ISO0+0QsQ6WhmnoSAVLIploBIlf
Mr7H3LsIw0TI860SU6nsWuawTDQw9N4i41ACbUMpqtSzRmZgLDCB31PtHricu/2b
b5d9NkPorM75hwqFBT5RuHyeONEI5zNwgz/7d22/Emzwg+ccOxhGsnXQW5tA6z6z
Y/P2XPw2fQFh11SQx6jt7ss3w1IbKABfNLnUV/3oy+JjHzvikVwNuTgmr96c17sL
xTPHSzz3lB0KeyfN2KFXURSyysoq8iEk0D33c5AFcpkT2zAyfCvtpqFyr8ek+ons
KvCuvBNT+MqotL4Mv3uLnpfFGu9sh/lVUvMubR8tV/d89RhypCkcbjPRKOjPa0bV
1BX0jo0JiO5/vDpcTUXuLUGqbH3ujlx2P9/pYN757gVZuXIR2HI+v1clG3rNM2Bf
pxDjKBAaT5g9EseeDAKQ3y1vdgneQl0HcNY+T+oqG+DdwjBQO0OxFepcxArMjUT+
GggQW5amiBYMNfTLegWweKazjRk0U6F2ogSbbn6TV2E1IVMxgOE9IZteuZMuQHUh
SYhWr5iq1QU37o13erhcnS/hi1iVkIgQgufhTkQrXARk2W05fF6WTeHKCfFhpNa5
YofzQt9RAHyyUY7p3Vtj1MeTwoAj882UJZW0MMMymIymTBpl0AsXKNnq5h3JqgVJ
qR+Hncq3l+hhRXVZHPdso9WPBTOLNIqdODBXbPqVUQB6jZpKkeUCUCoVMk/gV4Hc
u9f+pVIJgJn9NYmuNCvUyW0b+qEfMeBIluWx2UdW6vTvAgiU+hrXFiBlBf5MaVcU
GvyK0JQaP3qeGmLE7PYY9F1dzqcZvRXgxgwnpjQDdYTRO4DYAP6/xGAXnPutHP8P
l4EYovs0dhbO7msFSuKzYkLjRllQnNU7lHW2MS7nlyYzE1/G8KrOfZYYz8x1x7iQ
prD09Mr2lVF5amnjDceXzSWnNqNi5icYB+9On7nPLLraIopuQF0o2y0Z28IdHfGl
CQLjKG2j1/rl2ZZ+ujLSqs/cmPvOuE0AIp83p54VXPhlOYL1YUO9aUkMjOy+VwFW
NpcMylrm07CJAiXXl1gCNO0faxcjCeaFFZBPeqREvgnyHLUSc9kKX8aHSTwguCME
MB14BGiCrdH2+S9SdOXaV07VTmqN6FbR/u6S66ukTdEtLPqaIWxxtCP2JagWb8L5
5+JtH+CWijSOohYnwDVXduMTpsJycIRKFKjwONKK/W312cV5GYJQpbZdriBTsN3Z
f5jBksaLK8DBt2pTMeoOYsMV8o5d2sGa+WnGNPm7DzugYj0A5150meI78LBciRSM
6SxjgBaldSfhK0ulsEkbl3J6fQMevcNKGs/K6JSZf5/8Mzt19pKgwkGP6p9t+cQ4
eiqzapLui2MHxVIFT14Ljotuan6EotL/QehLS+hoj6lcHu60eW6qdjZx4rfDAyvd
DyVIpp+4xllkxIw3WMRh73allt5zOFbDwjwHI9fd8AsvIpvCsuuF+6gW687xHHAC
uuyO6grGklQpChqurXOO/8nWWfHtqvlWoJXXuIdXyM1L0Myddjxjl8BOtEF2FWeA
H74eM/PIFXcuLjN5rJJ4IZiKJXdfLf32pSwBBBwe/A1q8kPvVa77csbHz6PDayUf
2MhKFncZJ9JhmpbNp0TGyW4xRC074SZ+hWSrbHYHaJvl3m8ODhN2ZgPBVF/kQTVm
emDa+Q66lAeZOsdHDVyH7aZ2ToiiBHRxn4ElQze5JvbybNfkZVblH7wCXiJFjrDI
Glue8xSHqe/+mQzkWS9tORNA/PW3zt0mvR0qClnT7LJTdkyekcWb64LfV8yIQ/A2
JxfNBpIlaUKViIaEm1UDlrI8gT/pdIsSbGzm99soyndQaHJI/YJC37OpH7zCpOGf
v92DIEcp491n1njR10UyWuWAZHNobDtbegRk/x9d70cS9RRj340YNk0quiUtnKF5
K0eAIWT6dL5XZslHvR+1zofaNjJMq5XuDvSRcB+svkYLaUdOtuHnGu+Gh6lntmg4
aO3H7wnFXEMvQYMVdFR1N9Pio/ame/ZT/UF/kmswm8/lbjfv2irOyiUznNBDrGZa
YOQLX2m/ELkEAdYE+Mvur2xl73765FgtW5vavOXPVH6xH2XHQr3/hNE2bLISIO22
9Zo14akElRS2oQryLsYmN4JlezsFfYuvmlypUVQNT53iwmjGtZFUxE+iAKkUNfod
7jb/gBlBElumHlgvblfozUaRhsEl0JmE3aFRZ/sjXA7O5otpDGSQ/gt2xJ9/usS3
kWnDuHeoUi2oodRbJnGxL2ZYWHoqgJMV2XzuLYOwJeAo7WWB6hRy/d4IIetnn13z
XM+20g7TOdGRpTTLm1vHJTYd525HAVms4m+8uCI+Y3xqj/ii8kB+JreiCRzf0yfZ
LR2PFylDT/YfORXarJTaR5oXWNFDfXfYhFiwRgh2XDUilMKOFsuUauJkRnLZ5zy9
2OPjX+4cyvyztuivZbWtHqVqEmWUnc4UIVJ4NFF6ayNrgwwRXbNnZE8E6fHIvy4E
bUdukwih9tYmhpVrGh5FBleIvX2fFI3eWhXwtsKLMimVwgdIXZJ7jJa73fptuUiO
R5czcPGMKNHKPe+bDhEwNNMoL3r76cHMofx2E1z9fzXXhw8Cm+c1p5FhbeFKEl/x
6Th+u0Kgo3XcLKpqhRnhP6Pfx9r5CuBh5VCA2LadzVqjTUWgQPpic0KmFvfGS98C
JDWSXVNAY+AIbW2161HaEMrNn//i3RReWq484ki/REF4DbnP2uW/56WEjuGoZugd
+S3qdxi2ir/iQiq/aRle7wXxg4VQZeP+erieB8+HesmAzwFjeyEj3jns7eNueHxN
1o/8zmgGvWQFxPLj7haExRqtFmKtFU5EVpTQUnxZmMbdPOXNZqAbdsUHLf0Rv9bu
krShGemNqSejwHp9p97QdCd/pmqqQFHWhoYo8s87rXo2TqsycTVJVH6BVcgevidX
Dd9GRBjUuluiYxgRFFgC4WiOKRVPYSf+7FI7klsf/2rsmnRd1QbJHoqAjO9wNcXz
tj8XVkkkXRkyou9W4ei68AVVe1LLPnIhpbSQJF4j6pkq7QnqNARLlaRTOLSi/w/J
7yxWW8+K9e0QMBd//jEBmt4YrTZBDabz0A/2uRYc9Bm/36Y1wRwtk8KldmZPIY4K
JgW6zmKnKzN7plRk4IRazH5q0Cx3wl5Mvb64Jwp9g4qs1NwybNsLc6Ts5ghYBgbc
jtNjAfjOWc3Ngr3b0WV+Q50nX5dniOKBfxSgyE17hketzwQOkhaHxqiApy2m6RBm
aeMPUvo4D1d0CkpRHedddJFoJilW5M0i3aC3+tIKQLKuwkucWFycJWAI+PaZa9K1
Z69JJspMyQpt9qxEmntLRYmfTysIiPI4QUJCxG/glVWEVkcu7fIdVXPzPVjJyDOS
NiS9myFIzNAxlsUb8H9D/GTK3cRGYs9DmFm0uh6bAxpk++CkhjvvTOSC7oN5SwBA
VnFd5YzubA+YiL2Vi2F5GWA2oh5blarWBoV15Yj/ZqtRL9zNQIe/bYzNBQQxrGF2
4lgxwm8/62XIg7A9C7C7ffHJwtVGDefGOli3qRrfpD4aUZKrXjXlCDTZZzHJkfzs
jy3qdOwqIvN25olLFzPmKioYay/L+Tihp798D05A27YmutdhFn/W51XZjY/XsK6F
V1Je8HCevHdwvluweTzka3kFbgqEZTZYvSjTgB3fipsdBCrm55nPaDN4nwxPx1tK
427xhrYgFd4No1mGjrO6BJzoRcHXS73OR7NiAVzxZoxQAN9Gl+Vpe2yaTk8Sle6A
WGathKTUrcBlP4hhlLU/eirhxcJ6NLsBmOHrfCNqGxNRVE/K+y8MBuyYatRpqVI1
+1W6D9H1HgEG5VIjXqUx6MxKEpGFHEH10HKd3BAVIt8fF1UBU8rXqSbcg6TwEga7
um05h9EwlKta3fT4JtV1mYhAsvUn2GIaOYObeiHsHrOqdYNh2LhHlo4CxlAUehXL
r6IJLq/CIZxv/7dsKk06f1SzT6R2Ca6b0jOvgjvAodDjse16f5KbF4J75Z9MXaEu
oaALlN3imoue6+Vg86phciqUOui3krO8I+PxeOjVTEBn//t5PubI2RJXUJPkZJV6
W6vxaxnDx1aSQqq+PkjX9LCAXoFlm1Q13W0vT5242I+r6FOzKLSMkciemQyKteqG
5+fHjvEjTSLL4+CRJgj98HpZW8Wq2Alq7l76xoOQ+IpVLXWAVkwwFE72OSqas8Y7
fIi00fP0fp+nAIy7/OYrPIYsvXOX1/XPdPLOeF41j1kzzTwwyHF+5rwCet3Udh7D
PJCXc6QMPYY1wUR/jXMoB7yFNOqWK3qI7+Qk2n/ZyB6mimMwpLH+XE1YrsQCIn8T
5vdLo54iwQIrKMHv/LhnD8xRMOUo771Uk4tLbS+6gnYpFqKv9bHd5SfmIQa8uDOr
ELnSIRLpo/sqFWvzJ3B508MN05XdNSRUzNeSto8IUUwTzmejSPfq7AVZ1gtAFann
h5mRIWnOnpMGEMk1SFELb/MLJDZuKP6+dFnETNU0nCKhosCbRVnNekcTgxXOAb5D
HAosmNnqA44K/K4fBJWwC6/XfUYMgktxFAT2phUig80zUA2LHzTcGbbNzrdiIUf/
E1uztElqtM2r6mc3IVXbezMV1MOPko8agOuK6pFayPXwxOPX0jixcaPjhsfEvM3m
4RQijrk+uYc1ssHT0P9KrjhipCQ09qktg1knTdjiEBArrIjhsc2qXgzEpObT01Q8
ZsU1PX2HA98NylO6/po7VjUkandYhAzftido9jfaTedFYDZ0iYi58KX5yBBu+8bs
6XDn6eCAcQW40U5JOiyT9ecXz7TOhPNhz6lL8MlgYWEiLtxyy+xEoIHBrE/u5waM
8wgk8ykmppFi3LI+LjsY91VWEFhsFTchQ4RaaSMqxam5hvca7pYomO4JwD3DGo6E
C6GDYwegM8YOq6U73qjvxmUpVWPzByFoJ7JfVcVJC9JBOR+/fAal9DaRP+0HAt81
yNH4Q/dGiencbhow5Oy/QSYeFYr3FJUx3l/PYCCU4fmtVfIZCGoJ4eTDC6IOiNq3
ERxFET+C+OXM9QIasGlcAmZkap2VfGY1sloWA8QdrMu0uNzGpb2/cIM6BNLFMmoo
L74oQN6BhP8AT8OPGPIfj4M6vUa6COhcKOi0luiKpX/XJBvcLzT4W3LwP+ZTwEuP
fNh3KV5fOBoimhlYsreYt/z6fEkZE7knknCK49AVJxRHqzBa9EUK7Kg46yO9Oe/k
ed+5btD2emVk329oWkEeT/2l4FMiAnWI7lBxX7ui2UtsmTmzDZm/lJ2dSgd8sKkb
4ujijhZ6L998++5mtNUsaT43/0kv+6GSz8QKRvAC8yEitgm4SkCaAVybuubDcOa6
cBV5Cg6lpjv7LDJMfg11gKHJsxAMSZb5ada6TcLiLskF5JUmB7V1z7wXglZKMY/k
7C8fT4yqdWPSGC/33InxffZSJ1ify0jkgsq/V2M0e6edoId9T3Q7xemMdTbiMeaA
X4Cr+Nia4YWJU7VqNmAK/FL9ekBeCDgtVpDKA3W+Q4qLEt74oNe2kcHSggUwFfQ9
6mPbT7vINtdS12v6GxhtmjN4ddDadR95wimIfHZoz8fjnRj8eBAEajk//+gWuP7R
tBDOjS+Fit+im/VWYGXls/0S0U09LsgdnuumR5HXO3vZ1U8QSHDHgAOvUJ5TXHis
w+yrOhKK4ZPPRXe5lfnIFhhlJQnUBF6ZFqGsKCEmT0rAFgS3JWK3yv8VN4qscBHm
9JAKIenP6msdUukNJZJKcq20wxeREHZahKaDeDBiLwC878gG9UWINfsOSkIJhRIs
3vtrU9fw9pCBEKrKEkyxBIAKXEw9U7NkIvW9Hjj18U61cBEsX0vv14qBOQ1+nMIp
R5b552Dj0stbkyXpVKy4mcxHZdpijXUv5HVFpv3QRRCbNY6VgAswQEqrQhXpNyu1
Tb5oSJWExYAu6HeymWOeRW+ZVcv2pOoatNVdWTy8QbvXf6wtSI05usgYmGfzrdVm
Mrj+kP1WlnmxQYz+AnMuMGEbR+pFnOuUrXI18+DW9tWjgggpvsgkJOQZeetaI8lU
esVqyqcvQ91uvkO0y8yw2+AKt/DN+FsGPIzsDoqM9BRarS57VYHkr3lk3LD2mpf/
QkW40+WzNZyFgcd7+NiC0hJ3oYQxNYoJS7OF/eX7oLtk2W5YdiLzXkunzU9Zkxxy
PBdWm5tWoNePYOTt+MebMI3NOpsn+CYL73HyZl5KSjVJRq677EFYd+Lsdo7aqKHl
Py5LkvgWx5/5fOHVD3i8eZM2mihnjbS8uJe7Y02bgcOPqABeliYWdpAsTF8B+4Zx
va+ZSn/5z9hsIsugl4LBTu3HxysVudeG7j2wn79V3wMW45fYoFcxD+QgdFYaV/Rb
WVsJMWqUN3ZZtYlwc4zg0BbW3PE6RC+TQ020Kx9gUNXX+q6yc1eYw9B8OkettMUM
moIkRFf6gugTViQNrFQkcL3IJXFdxK8ApQdMylm+sFHTu3CAOgRky2nrvhB9bszH
VERnXdg8hMRgxwN9HZvc3Kj8JrLxa0Cc4nkxfzdJtXrCDKC+nWkAGlVB+NmxZ/7N
sd5eOu53tSda0b1ctO8Oa7JcQxkJ11cXdl+ToVehwXl8gtBVdK2eE54VTIN/fIfj
apJbKyBydyHrGOyrDAikx2IPGH0TRPV5OqhZuO/M5YSkmCoYPNeqbS7bu75WIlHF
2y+w2fH75YBC90IIMLqAzvTbaT7eXHD9bUZBy/hXLCDVbDTR3ZI2UGSOVkRta+re
EHj0mFnzYAyiEzv7vhPri5bYO9JAc/ohC303USr3ppDY/7vbkJhuAwuoQn7lCGOm
PQbbnZfUkBThqv5S/wz1nS/igMMnZCTa322BSQLiCOPEe2d1HNLy+wttkIJQt8vQ
9LwuH1VyAp+g+Y7MBODu5elLXoQinDcL1IbWRVgKvjKdEryZcO0z8MWO5pYu+lIZ
OqIHNkyxftOIs084/zOtsgFkrCa73KvNiSgTitaG2p4XcM5K8KI/bfwX72JgN0IP
8NA84chgQ+V2VQQjpEzvVTNnDSRCsfkA/KCZhB23mMrGKzMlupfLln3IBEtbvSno
Ab7YdXvl3PyKPyIxdmgwoc86KOIMId2BlLh6ob5DHGGexFyyutt65q39eOqpkOYJ
MBobAAVkzVAmZvHvY9awM/BAKx0sOjM4/2PoAHtqek+0fqV0vHUubqjE7Q5i2aQg
MFkMO6OeUfGhanXVY0s0yduTTifvIUV9AS4l84B+B/cD8ECLHhtTOUwswDs+nzg5
fUKRKfDEEjiml8VFfSeJpuLTQk+BZx2MeCNH0rdexkyrvZeSjxIQYxtecM/aOXwI
B0tRJlwJbf0MBhOL0njK1gKgDcCBdmfAYkihBNT8qDxpdvqikIw2vQ2EELbW+NIa
4df2CUW2qJhnmqZ/1MQ9JmF45uIEuZouzzHH9A5C5JqJco5L4/GXUr5w0nF1pC5w
Lu0rQxlrsd1QJjFhj9w3HUhQAxDsMkMbuymqy0TQqQH45fjQi3p0JUUTEIkBpjI8
gjxd5cfcIaZ9kVFjzF+jpEdwwJ9Qm6NLQIGZke2wdeMclqsGsM8qNJG/AS1G4Mc6
w6OPp8IVh/d6Ne4vXrM2wj5J6J/6svkvKAndBsWKuP3pvZfGxL3U+4UurfSHy3Ho
lTbBEWrm6TdxTUulOBbe5X34sIIofTY1NuPReDdY+GHJBxnr/SA3Gp6UZuXrzH5M
L+vM0aqzkM4ZkthMdrWkG2fzC1SxRv8dgpOsT6S3QhuU3Wv45O1+GHHU1gs9sSRz
88ibm3bkhkXtPgHsXTbigSZzEr6v7AOzyH8d3RTJ7Yf+dNDmpNFT6It/6cfFeMYe
DtnO18CyhCv2zLVDbhAOz+45t3War+hLVimSyjnXEd0AGfcXTR4OErCSq5pMfXct
D5Dm62PCurhRC+McKarRq3ek2x3Xfevw5qNKX48HPne0d0CNsaEaV9SovKfdyhqd
sFEuAwic996v9SpRRyUgeE6t+utLdh+hBUQtc6KVVAEqzqyhdoscHQ3kPKUFgp6/
FIDogiygYMokh9/qEvIr1fIfYi7+Dk0b/bJYVgLhv+QGgMz5at468LfKjdnpfpmD
HEj2+q1k4RVs0XgbLfCPM7lEqteNJrKh33OZ1XMUm5yY9EFOlN7e6GSJY+TXBwgs
ieZWH768qWrkqrwB5fUdLnqwcVBSiPi5Fbt7iX2D3PxonKdrqxn+rstYy32NG7dP
ZXky8TenH9Xodw/yG2F5IlkGAOXP9SqwXGBGEkGvIlMf+cKX9e25AwTSD4/Ujwmb
uaTW5P5YOAo4nBfgt1v3Po7WGzqTwaEOt6gE9GjQAWgR86SSEfbI4NNNAoRsrSOz
S1WOh9Z+s2x+oJBsA4pFjaju4AwJq/aiKZ+JbOqXrSbLRzUdP7g2GJW+8RhMF6V9
8f5RzkR7p5pW9fCqRfy/prBcc7ZpgjgYpAPBAbJqGw8ZKPbSYjfIfX9yuH7GfIil
DTdCpSV0eOPttslJzOPSDL6zbn1h0w7Ystc1XdjHKxHtWF6cPjVutk4CaI+MJSvb
yS2tEC+yclZ0nhqdFQOJ0zogFX/HNu7PVmwhEnBV5zxL/TqeSvMi0Q6j+VtffpoP
NqE1IZQ4nJFdoM1RKId51gnDjGlpFWUK2H3DRkbp6uTJwYxq6jqezUfIhbxHIlJ9
p/37JyqAh+wg2A0ofhY4ujOZ31xXnX7Ix6uh/oo+a7gXo0zaRGMl91EL10ar60Ny
eN/0vOcSStg1eMz+wq+ZSYA51LUOAk8RZXMWiT0CDdphhYcxIZ1sWu0pot948VsR
P5wc4ZGM0zRS7u5f8w188f1gQUJNUzErpN93qLsOWS1+kl0ELw+AVA4DU9jlj6U7
PeU8LgyHsFZ3/Mm2ihjwqgDYAmG9aUsL0Sjs6ZTTxyWLzDnx+tANBZZDyKg9W86o
mvObpQ4rEyCZmNRXUBff08rYRsXElxQzjTxK79RQbWIUDTJdAeax9J+5xth/EtFQ
ycIeTp5nDy099nnQp9qP4c79N7VtpiBuU1+y/+dWuM2Ee6YRBZ5Z+aBdCt2u4fz9
+jrbVJu3brsga54SDE/tmwcF6hILAG13/miLOXYPERjFaB/xoe5qFk6l5gm3Y/v/
R0YY3fCwf0KUUYYLJjWU3+QfZFxN3FbNqbIEjLnLeNIiqsWDKT1ZuX0Iixm1K33v
wsRGkTNZUgGnTl+HSYFfuEVfklcFGKfmVUqqPumz+Pcd2N56kbKT838bcV27+dxO
cKhsxkRhLVvvCpwp9P7XBskHsTWjiEUWzAhxEEeNC4hYHeT6/D2S6KzTSOiy+2xp
wSIFnyR4v8sl/5067uetOkrEfYGghJsfsGMiIJq0AawsaSp10T26Z2KB9lzZxM+u
kt+wyd5OX7pQxBzfQvtCLCW9aMM2qLVvmEaQJSqrxEKLsSi5zEh+i7l+waFXmi7J
JZMkw6pK+yrA1P29BEfUV3Ej2vtREjXFApv9Vmotfo3eei1PjnmTFLCu9ZyD0pQp
zhEga2jLj0OysJWf7Bywn9crfOu/KYX3M3XVmzyZ1xUaMj7VqLpnWv3BYQlGHiD9
r+s/eQB6WsKp8kGEOFbeXl5jB1Ijor2T0E1Mc4v86RNvgO6muLdqabDKsKJW/6zQ
OnHNvD5mCS+EQWFV1BWEtAuCGHFQUnpeP8TZb/5tkeR1Dut66SclSc43v7l/V9jm
pSZ4G6tjEurKVLC5wHXqkzSwxToaWr+kaNIxGPg/WF5emM7MheNMc2BUKrH8wdcI
sMEWHeTAsgrjjI4U27BjD6I6yt6TIwuNXkvP4SZ3g/0Ob5Ua3gmCVb6OBRL2LT68
x3TRa4+QXJKri6pNyzfM0m2KtVqoh/uGd6ygm4ffexVqA0QjD+fhmjUTmLfRa4Tz
2/fGOvzwBC3CHDcUkMGkWRxEvuhxJ0eHJZ+4sZUAU/teEFXlFm4rizopjxeoWmQI
ZIyJxBG1dGFS0qqgCfezoGJrHM/9NZU3guAlLsBuuMMXQFe3jhx3vDOOWtI2Wt19
8rW5zVRvGdxdJ/+OLz31zSpSSv4AUbTMA/tvkSHwgkPk03FH5OSbB8B76a3Yr+mV
i0mAFtAE+nU1Jc9HWzxjzHXNNg5AkTaYP4rL69zcUmkdPwSbvifJeo17ULKeVcIS
HTI0U1qsFntX/imCqs08mqV5KE/LEmQNlwAq67HzkmhPFLIMYk23g0gKQDxlri74
gFimQSQTskiEG+ExL6kRKHQE1FXHn5Y7V6gtEkukFLrAw2rKAwL6S3HC64J4dkXS
yYVPpNAsfQDXYB7r7XExX0lo5/A0sHYbOyXXw+jdjLdJn+2Xe1qHGkqF4XBGC64V
g6nZldu8ZBLSUqdoeVAt6DvDpgKnHUYPRzyLfl+/xcav1q/LuXg3J698jKtW+XD+
VMuck553E1LTwfZZmrTAZ08G1QYSm5CMzkSC7Da4L9iDlDfOZNiafKRLCVaaRBAw
xBCc/AnsEnEVPl4/FHd5gy/+ppkamqXw2FowK9Ju078Ow4H4Knmste3ly70swdT7
/OSBd3eX/JXatnnwzGk1sRVDClKH5pItLp/BoEReUoT/QZaxYo9ecSVXtXrLZIFz
+tqvLtXBTpnWMykc9t3f7UPmx6q7W0iOmuoYVPQ2uOUBMLnMp8K5Pe9cgdGizslE
bUDQ1+GQGGEwyvel8KlRWiU0QhHtPrEqSlUucefL/00R0wqSUZbmVVBxSiGFi7h6
/rq6zscPjfS79vM/SCNYMjmevnVa6yVzLfBQ2LsuPZGxyL6HtXxt/IjVG8aYGqp2
QtGeaMintqgkMdenlAqps50W/MImh0Nvdl2qksHFQh0UaMbCAAqFWheRxG+sXwwc
1ZH4IbVn6lP6VZ7u14iVtNlXplI8YnyItbFBIXVKUGGxMGBUp07RFRWYH4NA2Jx4
/c4U09GkItY1peH7Mn55vNqwK1cXMP94/WSIgXhfVQ8zhgxc+n+PAd9b8tOx31MK
BRtkXFsqGB1Un8a3k8sappLpBKYwxfrJu4dsFFQ42yUDbKtxBIiDUl2j12hPhybn
rLsp4ScPBtiGGmzMJaQjKoJ2dHkifIKd+zAqfjAesqyVQysUvkiCIwi+/Ze7sLVX
hHuVjdS8aD5pZgEQ6zudOrI6Nit8hUmbW6P2HTk2lSkmiGH6Ife4pMfiDfbx5wsG
5DkLDHVRBBQsJAzpn+JWPm3q4cTXebMAh5gwOK0P5qgRnB3dmvR+pWbcnW8EKg9+
0ZwQmpQLy9gyDjfttSokRy+xMC1qQrdMxaCoDm+LNCIw1la/G3HyGLRSyjbaJrMf
7F2nHil5o5ziUkwazMRoC5rzLPIjq8EGxuBruHqRhdPyrPppTPCWBuFpbiGEcoXu
5K3u3J2U3WkJeV+G9y03ji8VLetOCu6poG9rlYWBCZkrXieAyBiaVx6zoqDbjgb3
a5IDB/hVAYlOaq2jogN2QKfOBkxIDTIwXlN7ss8H6YPE/DQWl6p8geNFGtnHSBTV
ZXB/mEY1SuZjtnuI1ELVY6e/bsJvAx9CUYPDy+jQKVegBQJuae+vB+hanI0nykhT
xJXbejUzONhmhDTejQcsSlcHQqJ1iKxM26oPzUzdsPE93ggaGvSLQM/OgItcaek6
Dw/7Oz/pLv7bwESo31ZPr8qW5YTiqMaq9ncD6WsQfOVSsLWSUUi0T2RnGew+ShWL
z78hqqs91RFhREjK7cEAO50bEG7tdeNNe7mBlcxW6RSZBJI9yO7ZcsR0usU3ixWh
ws5/Yv7Lr/yV4AWZKOyLqCe8jK9dvV/XEQ2YOhKLZDmUQ2iPLIn0pkJ221WIMsy1
jXuCYsBDAuEtYN5V5AXgFl/jioNJOD+f/Fsrp/z1qP70pbJ6/Qub46/Y5PSgkssE
LZholNpIVdXP1T0fg7+D3NhzssPZJiiJGZlTd7JVLDWiCUk3Do2+LtmD/HEfBSqb
Rb/Ty9pMgDUeRZZC8PY/PPVOYCvqfJYCOQU+/i6GFc/bBNbAF3uZbxI4ChLnBQOy
lZmhv4Vs5uVvpk7kb+eIpRCIP2iVDdr3jPTX5AipSy0bz1mn1Sekl7SdfzsknR+Y
5SN3paCRrUQlwl9R2CTPUdNL1qa111Mq84tk/Aqh5xPGnFXnVnEjn8KxTHQEas3v
P3g5XLK06YQdOFJWMCVX3hvfi3K4Q8L3kUzDtgMeQou495MxI/Tu3I94yg2Kce1P
z0jtRQz5IX1/pX4olTzpC21IIB9WJBdlOP/vy3MTzzdXSKYgfL5/XIFJBjTeAf7S
qS3zlc43IMkVWzbQ8XED2RR9RJlxMR6dulvJaUeDRuTUSgPulVd0CgKWZ5TwE+Xa
lplGDoAlyb8VVMz69/xyzIqpKkebnbVtqox2m4TPezVUknXcsWUFp/BbLLl+6J/e
47GX3eWcHJPBmxxBHiyOU90NFw4FE0R7KzC12c5DL59tyKDyYdh8cujfUCZZesuS
nrSWxCDvuOWcz/KvbRZAeAGDUqMi3p5c8CT1L4C+lfaFsLtyZHf0wOzndoP4Z6Ht
Ld34BK7lZyFk2m00XeWKX3fjJKYGVY0mIwyqmBEDQr1tjVjNETAwIICNUKh6Vs8p
TJGS2x3VPcF/tpa9y1iLfs34+7qO/PiftUSZc+wONeMyv6ajWOI+Z+5LekwVEJNa
kk96L67hlbUyERX5UpQRbpblgFkpdAFnEzf6O7Kg9a/LQn5GRgahMiS9d5DovW6E
l3aNOGmO92yKcgP/+BtE633jiqWrkv1mX7Lc07DRrqL0nRi3x5M7XCysEzy1HwcS
GV4O064L4XU6htSs/rNZKSoYCBjuQuN/Yg6q5kSpPoRdreotlycGShgiHlRO6f/5
duyLsBH0xvfKgQNukgd5R0hDiSSwOPWDezTFG5Opi7NW20JaG1iVDmdWOgO1sB9u
JY59ah2+PrfjUypQlvXgJwhX12UhAnXluGW8BokXHtV1+anRzI7Mys7Ncotxw0Ev
m9BBgf54HCQDzEKKGRUVEyXrBbOGNmVM9EXJFXz/scvvB8vJglVnbZGeBL8tsGvA
M/3Q1L3LPAskxEzZGzrlMx0z31SKFpf2tSgwlBw492ceMxf/qQaUTMznl0YeAT31
6CeIKq8PJotp/DsOX6Zc8P/Wp960DMQjjnnj+3deS7Ia3ihl+VC+3Rsbs259sTGn
Q4Wr4Oc/J5FrbcQzTKiIbaAoCMp9DGwdXiWHdq0MJxkmZiJVmgNOJi0kVN9NRWJH
9XZocYI1rNJyzwbUKjQP8zgGEyR+WYrud2KxSVgpk6zEVZIpFocsH9yYki3Mkclk
jREU/lFluqujgWIA3F4Fa5Z6O96pT8ZWNKvP+BN2ih+f/oPo6bl8Stewjjtr/Xe2
GG3a7cur48N9qhoiw+ebwB4r0bJKbFSL+Roa1et49R+Boh+tNcr6A6wuI/nUSKH1
LzRPZl8zH6M3Nht8wiYsHJmHIb7JE/ToOdEEv7ov7eglQBbdQN7cya1ilUSAT7Rt
898qnXuO4CJjNC6y5I+t5LNERrXtrPONFHzpQBEi/7Lj2Le86NVxpNLzr5E7b8b3
ccitXFvyAeLqDtow0fQ/Z4kWWaTAsFIzJI+Veym3fkTy27+OB+T2KMNaVWRNLxHw
DbJsqmM2ybw9u+0QrK3qJX7Ivw6AchPPFhKp3YC1QrnnMk66CgKzUYkXCJPe8Tnt
iNSyRBUfOnysAylz+93zRZDwxniQ/cx0d7ejhX+vF21z7LzX31DMZKeOdVs3aU5T
ET2X0nzA3SiX3CA2b6tfJRLskF8u1A5EQ77eloV/qOXfK6qKel7JZkUgMhiNjCVz
Bv/euaPDojA8cz8BSLusCbrmIoFf14Maq3Oo6142/o2iAXIqVPrX2F995uOyW3uL
EmEBwTe9RDWs2HgzOYIepQMUIZq8jenbvtB8ecjOd10GgSjlqeZXtOPifFBwpASr
xImxR+Tc3tjr3ZdSla+4Cz89OQJYo33M9wwBg3aHvLpKXxHhuJs7sIQC8iFxG14c
eWZaKo9kohya2uFaK9qXBqxaA5uxtnq3tfoe3RkyWu2SLX+IR748joMpF8S49mW2
0hmyQTG3FQMwurumY3qkdCiWS1HpH3dISgCrl1yRtidzx5YHHPmhcUFFc00nzZpF
y8jrkqgZuV9O52kfHV6mUqbdRW5VuAsCtTE/ipojZ1CPTlYwTbiimB9ccEW+R/UV
B5j4ZDgtLRyraF398ONehQFjjqH/DQhRKl1JhaeB7CbeXjix3gDfDHlnc/GwPIkG
FRPMgkb/8TSJEPMUzgX77FZxnEcM2QmRQC6hhLCVAzj+q4/HhVDAjF1eIPbN9h8z
4EyiHfh+oVFlhuwXLy/TitnGMpfnqcCK1FQvehOOZbJ2f/pJVacICXq2GidNwuBi
Ep/drwMaGF4h0BzKZf4TJGDKyV2V1nqAOj98nxG2tMhU1Or7hnAC7qVuRIzP/7oU
YrONYPtlDHs2EN6coP3wPHqz2RskF0xdYXLP4CMHZNimAumRgzoU7R0Od+qqntKQ
mHAmj6miNHLNp25h4i/0URDdTZ5raG567oS3W9J2hrK/9fkQijpi7Pl93IkTaWSS
WdUP7MLSCCwYv8fGxoiKCe78OsI4HRc/2RPUAxMDFFCEhfRi1oowYWuAmCw94cuf
X/pgVXpiLpjZ8cYTeM2AEWO/uWK78aLVZ6KY1fKgfjnDMC4tror7PBPe4LtZdI7v
5F3FTBR7K4foSoH59mMe/sP00j3qLmvkbgaT/24Z/ihTmpE+e7KcarM0AX6L83BZ
DFR0CsF8/MHEQXv1D5QEf95TzNdleeFCsuG49wj5ckaQ/o6QB8tOcEZ633C6YPK2
Z79oS6yUCLk+MMxUcXWY2OF35HeYhChTY0bz9VrjxutQGPcERRZwlStzA8sVbd3n
y8UfeIQsjWz46UzadNmQKJcf+5rgu2D2cNVe12j9+awhYLhOivtztVvaN4l8hX5A
ii3dn3V/6K97k8ojaWbgnQQtoy2Xvd3bN7dM3cHyMemj+1zaUrG7x/S+QaTNcLIs
n73fuyEGAqQfTmbM0zzdt5Cj50spPcvGJNMvVGYQAQYp1gBYuFZ/lxTdg6TdfXw6
6EC9ungiAxVfOjVcBU7FQ//m3B5hmtq3ZU90VNi/Cbha79xGlgztYZDEvEdUh7Ma
0NNgwG37hH3nTrgvJ5uBvTasx1SueHi3dUktXRB8koU7f3u7p7KqDPgU+o1BT2Sf
K+6CJMJ8cDQjZF5NrV7jDqY/iC1cun3NHk1iYLkuCdijiVzl+LFQcb6yTNCv37Eb
W5rjSrz4wDYlutyTzh2iYcw8WbqM2lf1VX1mWfOyfgDZXNG9JciscCzVJZQ+3r+T
Q/buBVaZi2ZLkSagbYmPBtSyGZRNuUghXtD/kq9zFy/BVv156rI1wv8eeJp+e/QK
rT3ptS11X+Ojw6tIIu/KxZm83fY5aO2VaYOsKKcQYLPap9jWXS2cWdYHwXBqdNEj
6T4Z6XZpTPbJOsIYRtI+AHD0dz3S6Z8SZZ14GC+BQTyn0MU/cZGqxnkqD15G3wYJ
lFSs2f2UK0SINzvsxHNRSSL9KgnwNW0xMzK2ymrQu6Q1Hv2GQ4XpILsYvXPlRCmC
DeHYM9VLXr4OC2jlvmUfOc9q9yR7XmsBycnX/OPotqyMWlixmkxKzVsd3a/cU/Hi
s5WebcmzRBRnr1yGMMQUnl8VUO5iRxicbUCMfumB+C2yyjbCFjJaohjw2pAIKnqD
WE7YV6+OOZ/dh/gzfNsrBFkBgBqWg3yx2riN46no+M42mzxsEgEffLYGYFDXDrUh
ZFr3yS8wwI3M0fv0nyggWvTNjRKEKNoBU+SvfvAt57W+lCRsF1NsEuYbe/32Ay+n
f+IMPoCq8fUG5bYW5k62bOm2wQMtmDGPha8OEbkNTPArDzzVn/N2yEE/d7pepNy0
oKSsgu14+8auhNc65Q1Dxaqfxj9QfAsFXntZ6OBUHzH9oSucM3WWViMLZCuZYyKd
3qMcTqqRxvHb/zQaKaBYsl0Af75nDTlDaZPSCZcgiNllsWonfv83QZfS4/hVNfFu
6Kzm5QGMpWmSILGy+MOlYSwCniM2amgLPYJ44GTgieedNrz/LrOKn4ucH2IbUfMs
M8As2DhSbpZ3qMU9ruTJIuI3oOfGcaPTKpdcjk8ErRrTeWBdBPfk3W3Qykmng48o
qOL3GMRw0jKiabNSGIoDTsDAy6sDY9H4fv8pGwH7GaFUFS6TdvSgyT9E9Yh5bk3p
iyGfyQgdWV+5bR2A4YW8qMQS4EjUWiYXMi13LhjQUuBqUsHycBH0sY5h31sIEa35
CacJwmWvgpHx5xeVUpFxK10+/fowFkMovN3AA7iltSyS68fLEy9ubc73pj6Sc0Hb
vzozCwalXm3CypvJ/xkg1mgg3IR+WXm0YNOl6WxlrWkfUZsU9FttfqLZkV0Ox7SX
HmZvcVmG98TEviCgtaGU5CZbl3FrQgHHS1RGN5zq9T+RjD+TsGwBtxs5NvbXp6uX
tCuOCVfbYImgeU66WRq47F2+7VO9WDC8VBORnACDCsaaIrR6+cvnIR6+5VTm4EST
ZRJiXuWW5GXXpqL2l7eb6DNIXgq/x0sIseZWctGptIvJDlC4WM5gmH/vCoJDWIN9
WB1R8Z2PrNLQglPbZRtVXsiImIAAqG9HFCakBmRRO3m3YMHEX45uBl17K82PnVZZ
WCfklhjIEu22i9s9smUnF263Iaj61lqakZAkAPzWQTpWq5/B0bKCf/Y0lQf9HD2x
ewT6mbgPnjdGjXEKZUyfd2C4vq6ZTuOa1SGyWiRR5UU22CQ22kZhvP/vzoBKhFMQ
0Etinxw4HMpIjIGlfew86wDWIBw8NSvp8Oz4qnAo2sYE1w4gTY5/g+6Mm+SfWtso
jaGEJBPaX44JZT/cDscaTw1MSjBX7t+mDTl6ipgBYsGCEp4z+C9SKPfuOvVgFcoc
/mtu7TmuA3WtG9IZagVyiILDxqKUrX7FVNH1WUlaCBi5N14Htc1HtjskdLeLs+YZ
g2XksaIhR904hEJsenvVt1e3OknClRBUr2jP/JmF+jZDpcmPs6ktOySBWVCVVFmM
w6Bc4Odih0+rEyU1i1gb8Q+Ul5LVjOamThBJDYvA/OAht1dNph4ybog9rGFECA+J
Tp988bdxnnzb53D65cenFvNIbQWZ8H29jRhireQcx/B2STddkqLKAmE+tQaPe+da
5m3gD3sMbtJPJbSbRmfdvZWgFrEbAlMwDO26skMlveDJ+cMw4kGIWFwc9CzdJXDB
jnIB1u5sj1ju7oAvcaOpxdNXszkFsctYmB0acsv3xFTf0MbHBI9SCo+ABmQK6YfN
5sqAEuec1TxssMsHb3leNT1Vr4Abs34GL4NyKggCmMCUy0RKCI2pr+uITy61xQmr
4/zD3TtM713cZNR9L0aBHMNi46cUSZ0YKkSlooizKV44p5kxOJAKbZz0tne/TCOq
sqyATLeDLyXnvQJazn5GsakPIkxf8FCkRxg/f3jk2dXb8zSinhV7aYTz1uIH6epq
fvEQ7axZC/ALy4zK+30jiaHD+0qxq90iYqha2DKs7inwtPrP8mXsVn8wlj26Warr
hMEB7RfsEtIadqEx1fvxfMatHj6MZL2Olfe1D8uvn64Yt4oa6vQh5j1IfPNgxPiy
CG5xBNfAxW/S6xYK1M5dWQKrxoVicR+1eN+7JSEnrzEYz8FRv8euRU0BMxi5C86V
thR+CXqp8Kq7N7Qxf8iArh2lGJ2p59p35la1yI5kwXdtpGxujQPMLqFGu+HsmG0/
+32gkQvDfli4UqaDmMajMs1JAksmEEg5MZ3Fhr7KOz6KFSj88ZxKonJdIBDUR0D7
lTPpYfYUGRktq4ZBQnCDwtV/ww9gs5EvhEUgFarvv+gjOS9NFPfwAPU8tl0c+x+w
UzGvDvdVoDjbaKLlADCBGDhzwRi6SO8hMY1CHFQzrpB4tdcwVDOoU3HRE097n3Ji
MtiCL38yWnhtD9qBpNP1KPJZGLw/4bVDhgI6JWFRtTR00fs1TlMFGIYopvvGzQ0s
b5cfogbSJSrD7AnYmXl7gJr+061SUIm6MzuTDk3p2t9tdedmNGXQ90xVvGYFgsAW
E1IgDEevOCZnOLPrtD8ltzrlSuirX28N8iKof2dnuQVO9LXfJLM+Q/swGhMujQKA
qtpl9ZeHq67z7UX6PCDkESN5xrKMQJgCrLmDxLNwGnaHSNDja8uhwF07ysm7nnB2
14OHdJ9vs4DSd3UNYfmI/MH9361Qk3zofhkKhsQSMgNUGKa7YeY61eguh6DtPsiK
Sbu3x+NTJa2uPqGH9jmFPTt1yVdl5mGysx+4f3hOtOTGoF2oGh0Mkes0w1R/SLO+
IiR15dMx3zaihwIBRbp5T3CXlxdSzMtHg7Offf19Bq6j9+NB6+J0fDeUDWzdjJ5q
fknGFdc42hlHwkAvgw2zwSu/UNym4fCXNNIhKDr6n65e+GHMMHjn1jDSyNmGnBL4
5FkXWFG7d6EQ6WQ2IEJe65nS4ALC19Rbp4khRsymfgqgcSch+bJ60yoiEuzstn6O
6L85psqlilClM0mYbLwcKXkQKv1NoM7WlziNrMzlWjcZmMeKMPQAtPGn9k8q7yfF
AHQ2HgwYiwO2WZ0fLx0DHNotG//E8AlP+kBh99N0zEZYLFyxEoJpHdiLkEtIyp1n
UAprQTwypZSry3OmcYNz4mMNATIDsNtmHw2Pq3d8xxjMdxm3eV4BQpt4lM+0VIcN
OKk4DsmSdLNSJua2gJbad2lGkjo3Ny3WfSp90IZmn4dw1aVa2fJaPZBK1BOwlhFr
Wy0v7n77YdMUjumL9JrawQTFGFmLKMpTQAzvoZ2AK+JxYXsyTN82F7Pr6UWWIgea
QJ/gYEScCSCf1vdtNoAdGr0M2RV0dvIML/sKSdT7vCUhnAymnWd8p0oNIo14i3gv
PvhMms7wIRZmv3Yw40RtfueQjZ+6EYTqWfwY180iEGyO6Q77F40lMSKBfqZyFvRr
CAND4ywuPdJ2zUSIizD4dGKLx7RPwy5PsA+iRhD2nqn6jRtKuyTo49J4ajY0UbK3
2sH6L0AAeaqn+WSpt7M96dcUBuP9i2+R4dM7smvxpCAU+nL8Zovh8dTmGJAzcxxg
JnBXWcppqYgk+wB9lRUOQqy0q/CQJdQZI5+Ple8SEM02bIOL28MjRYnKG29M0ZA7
KoblVNWeaD8m+rWgyzCK0+IPP7I3l/X+F1Y9r/3fzuxBoXtdxlNlLT5dg6aISlbg
sYuwalHqYaB0wIk3f4RPmLAA4BlRH9p7omDQGgVEQslAkVXGibMhf1XKMKR/0glI
LTxYDU1d03U14guQluwtS+b1vBm8lNG8oeI1VaD/VOw7kWdOQOf1e1fz3yJ2mv25
tJxtF0AHoKCNYFhDFHKf1fHLudhIJQTf5pSAT4q8mFaTtogWhU5UgKuOLt148qQy
5Ns9kwgXHnWoqzn3ku1oadthKMoPbukRS2PRfIlUe1gqRPfvhyUtt/FnP7gu0O/1
ypI5QRE5f/eKG7YJdzRKd6/WDSGbQoXEybZOslGjfamWIXnM4DUa90IntUSFeSJI
El4lPLuHC35ScpR448DrhYT+/NgBJfKi39NPCrn+zAUov1PQbJwvB6N+02pie87d
3WmTLsYGAZtnkfzQZPCq+j5+AJK4IO1UjoISqhzo+DHOvJUhmrsaQrIb6OpcBOCh
5nwcPLtmT5T0RtbrDi4fPqVAa8UZnElQlgoo41GYsbeHRFD19zQZlWskAbKrqvP0
mQeEHFjvH9nDC30wkoE0hF4HZCE2FsG/kXfuAkQ6qspERZXiAInh6OWnEP/Hx+vL
O/npw0fRMZfvZsoBF5HDIuR58XRnLaY7jV1WedZNf+NAqMF7u6hTPj8tf9yvpli0
0s/kcm2pWdyD/Pv40MLfPUZa+zEY+C/mzf+55wZEhuxmlB++TokLZfbRjusvrqhc
bz3gLPgnReUF3qdZCxBXNFnPVpvxWbTgsyPXL2w0Q8W1vSQBdxlIA36qICouzw5K
YwB0TLGSSONxHRuOcsrRwdx1alVhiQ0DWdeUH7fDQzUciyzcBg3J3//iySXfeIqx
uqpmJb/0smoFAoR+VT5lHTSrRRryCSwwgx+fu/1dIrktkKc64eC5uRAGMUiLAqRz
Sk8kNrFDypRlUIy47sQoNYrz4WRFWgaRYlS5VWyH6VD8ifkYuX07WD74bkFd0Nk+
q0943+zvskFyaRZq5DBnf585AHbK9KiKn0rdVG0G35FbFZm2ofGoQehgRcJS4eZv
87JfGSJztlrvzfapTChCunUaZUON5wk/nToXF+zIgJoJpLVngfm8bz/HSM1eMyFy
ARp2lEguTIcEt5Ty4f6+AWnqT53pZxJGs7NBWDZ8P5pvbm5pS0Ikpkqt/r8/31Vz
UaOyztSuUxgFIe1UWDOZZ8sZXtQ8DGj7U0wceU+34SerWKQTHwewOGPdrnBs6Aji
vuUIgXzlK5OmU4COTWsKTL+MNiwR+RTzrs22VEsFSw5Sfl618oJ5XT2ImHev78bQ
H2u/3wkzIq0/0kxKPr334P65Ho9QvTLP7/D1F3igrFrU0l4BvrRP9FSstj2bR12E
rL0uh4s98Jgj3syMuLpqJWEpuuzJ9zMssFNQMemDL75x3ecBKgtQr3i4neXLswP8
M67aut1ISPM7Dd5LNes7XJasNSFdCX0kqbuJ583JYmmHrzp+03NI1CjQovCufvJx
9wrzUGtTW/bVxxghuLz30yJe49t94NtEBmSZ/5wb9WxVWvUEqS3j4wANEHCLBXL+
rbIdQUlhfK8G3YHoVNcEcS17I3eLtZ9x5gRHVGM1lXKOxjFxQoziQ5nDBdpqXfZJ
MeaBTgr1HCGp2BwVC7x1vgnBEWGP/nbuq1J11BiGCap1dOAqI3tuX8ZV++Tn+TGn
6ERDDpKighJjhblABeYK8A2lHj4JgUhr2GtpQxhVDmLfdWE7shq2nTLqPXcCUDxh
LqdDwwxwQ4aMcZMngyfLZFzAUsz0a+7NRCCmWJKYgfaFDJwaBa7K1dQEWFaiIYBH
3+rFKsNcxo3hLdh7PmdWtAYWGRpvMcvr8OplJXV89k1Ti+oN3m0ZWPlR6fMkqj10
o1YfX55pQzmvSgVhI7bFrk8wO89CxKWb6TXcGgpUH2kMXX6OgUOp0eDwQ9c4RJtW
0q3HS/DyEbSYPGbZTp8Z+C/mq0fPUUw+geW2EcTbDFsWCY6GKyXr9r2/4jc5orMs
PNPiZQTrR4fSwWNFgUagpKI44g1G+UYcOgSj1syzgzUXEPogneaqJfID09R7x+b/
WEPWteNOq1hN85x7A63CQUxSjxZ43Onpwr2xBD2zLGADK0mz1qwhwZXYszAM6FxP
g16EN8hLKB8oJT7Fbt6vWLWpUBnXLKyyB5ibwlRX0GS7goIObYu5KxZ0rp21SYei
X3cLctirNN0iJuaaSwPglx+E5C6yqWDM6qufoJketYx25LQYegy1sjfSsPkuSguJ
llxEHb4XzKi0hDgIDDIUWQKQaaGpOGBYhZi5RY5YwiCGJDx4GSnHDDbVnDKrt3lZ
/HLtAX05NGCIg3QYUeGrXVbGhQAzyIPBcEzePtSYat7mnddGei/a4pVT1WP7BAaQ
n6mFaURZgjCyzed7r9koPvQL4ORooJYTKcQqrVyhzjHJlt3UL9ikIjK09t7s/WLJ
lOmwSqzZ705Tn1chdHa1oOIhc07NlgcT+aRJ65/PKC5HtlflbNQSm6g9wc2V10XQ
8N0mhi5JYQURx1D+ED8MPyn7bIRpdNSsGGPpft+XwyUzPrZ0d00c6+MjxhvuQiVv
4CfOeBjWTFofzFI1IKANS8LDZlrlkpHT9gqenJXOd70dWAvHb8D7yIuGCNZNVJmc
S0IHBqJdxVgnmpEIqt7wg6mRKh3/4oRUmfJWGD08p/6z99YPFi95428XNdbtUqSr
5MEioAttbvu4Btoo/07Ug5YwjHFFLiRzxO26e77rxta4izkj0sQgAxO7Zh26m/4L
3+IUtuGLuhGJipiA8UP3Poa+Lp6RsehwM34Mo1RPaL/2+qjTQjdIlIQm6aUfZZqP
iWEztONzadF1bZFIUssrv9efA2Dzn9Pd14tqETLFTra6II/hOHrQPT1KZb8sDpxh
ouCPv6iAO7njKenHf/Du18pEIf8uA0A7GuiYeKQFIjpTawCQyjsV9H9DTYZskoK2
wocmSdNkzzMm2n32fqzayhOuROzgpTWe94F+Rk6GIQyxjFbuOyy8y8MiO0ECfHvb
IUVlwKKfv6VgypfrUg2G8IzZ0AcTP5oWUh9S85PCqJ4VBnqbuDoxIpVnKrzsyb/f
aSp2xogwoYF29I72DEKq8WdPqXHnZwvOaoNz3W69m/viySsVE8RP7fU5JA4VVeu2
CZY+uiw6yWVLg0+xAQ5yzuro69IzYuo60nbCsbObrszbWG/Lw5Ay83EC9Q1C/e4P
3cLrDS2NWEsygK9J0Lg7M2R7GAYynMgomAFB0d5lPD6/EyUgP+kSDLOokz7+A771
1my3+WOOlcTCLJ4+rvTFqJ456NxCuW8/l0okRhahWND+gCY9kRMygL82ctrdDt/Q
CTR8keTn0wrMGZhMxVzNfAnW3yS++jdWtcqP1ZVU9DsUYFySakvxb9qXhVmUljv+
wF4bzzktiW9EwtqzEfyPweB47mN121Zb+KeLcX4c02bvrQK7BBt3qoNszao66zw3
ylf87lE7zR6uMTd1xVBFlXmMz+zyPO3nhUJZM9Nf+Kse585ReMuJocV36v+6fOHR
0NTxqPOuBEaPxBBwB3mwqIYC/kAan6tb0DYyKoYYmLE9gJMUYD+fcWp/9UVy2qah
br8btxxPD3xNiYcqFeIeOM5r3+80/3vGkUHX1kTbitlaPxPJqgHlsk2/DhVxBbbB
aD75JUqa4eLNhnHVOgndazJdrfJF0yhrE7v2hFRByNlMz75zONCenL9cN3r5KEFc
JO3pbo35t1+vLJmE4VF4GWVt4RCG6f0OJp1FyiSn3SWSlIGnxZIT2ALez6CuFb2X
b7YpLMuIF/IJ8Saqwide57CKGBD2DaNyuGkXSlkjHHpU04xm3pQtcN32ejmmV9nm
ytNw6DNWDZtqrEjLI1GGFe08S1gAvRpyICUbHSpBUcu2TOuD9bgt9mBS4v8mno8t
lCd2RNXYrI6PBEsAAcGyGnegHCggT/Ku+MZiboDhzH60NL9d+OY3ORTUoCBtEFPB
7YZ1ARrJDdDYvo/zuTf44AmHDQhYPPClABwe8hgqf8+Um7p1LI560JIZirv1bIHo
w349qwco1HTmRwe/wnSqjXO8ZLwzapwpUQDyXNYSRY/8Cy7rdkvM8QrW3Dby5lzk
OMzmgywe5hEb20/mmOreIKidwJs+pYR3jN6ZoIRlnsLn6flK0HbY1wbk0xXlGgQH
2zoWuWYsiihQm/AQ51sccLIRBwZ2aDxi2AZNu15gYoBrrFP4voOKMFsiG9caqU3y
Zt5oU2zWTuVu7PK2KDftqwQmQz3F+hFhn4MylnlcKizara/pOORUwGCl6rBen+4r
Cat7kt94BYj+DrlPBAcgv0b2p91JoB7g3FeA5RA05NQNS9hd7T58BFQSTHWKLGFw
0sZcYLCgWUxNgMsLMwqXfs1PvppKVUfuHXKdLgjYcdK/EUGfIFcOSa0nPzNjrLLQ
6Ma/uhbLZvjWbxQeyolY1InhzkdyE52jwUgHs1hM7ym4H6goFHOJmkUYMyz4v9qB
DkYLSvUkvpnFUzhYv4wfoWy6ZhGyNqcSXsiI8QwxQE252DJDKAGQG9i0M07kmQVC
VnJwi/mz82jJ58Fmj64hAOZqZotIAnh1+3BBbqrTOwcPOdGic4WBS5khZxXNkWDr
p5SMtp7igqbbKQ9XXs0LjE3HPzIefwEr2tlRo57noUck9ySK1Z49+OaqaoxUXB2C
IoN06wTmepnhvSlLn/1AxiqiDcyZY538yS2hcyNP2L0fGtYmZI2qoBMyoMkSXrkr
Wp+I7xSXzaqUcpJpugdtc9GWDNHUj/oqEcUt4kg2AyzlKpDF7eNmUtsRT631BA11
q13oVpMbJhjALWiixsz0jo2aSddSCkSDXoFcGcP1E99zf8kb/1SaHq5mziBJfRLU
Enh2z3dirqBC3bVtZnsLkahw+Pk3uCZk3ucjhLNF9uYoei5h8qwqfeZ6tFKYja7x
LSzeZEK0/HGVO92Z6/x7P44XGHWQqHqYits1eV6uRd1psM+yYtpjzLVznImTL85z
7Lmm7b+muu4o3HcCvrev+veYZRcHEnRrSarGmFwkNH31IFTka40wqCJmSIh1NAXN
72VBZVPuwqWwMCkynxuLaINX1VHb8t35GKnK0rRoJSDpWlNKRWiTAmeLe235EA8y
esLhCcRjlgbfwf2z1JEXxs7Obw8anxO83iBHfnJDpwHgwZhQ6jy5nUVxYuwOltlz
ifyaZ7TS36zzOKfv5NZIKl2gBHUKut0YitbGVSB6JB/Zr5czKBqZ55TwAXRpDcZj
gnv/ewA3v6bIahAclp4EzJm0R6XMttMSJ53W19HL5EYllxTg/hwkGbka7MMK3w2M
XUcIBAdl4v/ytgBi7hlEWVj3Lbolc52ErEbwg3Ze3pp3/EsTVnj9cr+pb5NLL41e
jgPgXxNz1vhaHvobg+WT8D3eOM6NMUdnjNFT8+7vJse+UTAO+upvSn+zi/Pwlrei
GoEJ/y9JFsNOgry3tpOwnGu8xq9+m7EppqcTKKVhdOh2FENKqDxp4N1gBw1Dei9R
3aR36GLKjt5a37NkoN2+OOgewUP7RSdSrenbXBFmhMaUZIGSiJh0W+P83ovh5qEs
dA3NjlyLCCIUPSAvPj0Si04rO+NtXLkObmcHOMWBFDyc+q+Hn/O9G31BaUtSY6YW
0U6yfKNTQtyzgZ4zyiPFfcUCAq3/PQz3EP1XvjFXDp0086l3gaNhZV3P7oWtDaCR
1ySINFAThGo5vExCgIsT3KWc3T2XV5PuT9eqW9g1tKFnmU9Dzf6UYWdy4OuC23sj
GL47fZU1ipjzNarkeBpFJG/KrK7tfKFfnxJkPKcaWjrElD3v9ckpfpcU/aSWxLTY
0SE1XmNizoo1tojIe5G/oROJlxRPLHoLnKlBGtLrOp/Q1eRl7C1fKpzJEtJjUs+a
aGFSqdDHYjnwWrSgaGyDSUtt7aCqcHv7cMfm+oF4/Wer72Khvrl+l0AyOoKBlGsz
sGEzpXYpaPLqP0BG1BiN1CVlKQWJdfuXsBrkGNwJMPobvy+MU3B+2kf+8PFWc8qC
v/Eg4Pl7eDQslRUJGLFSY2gnZVgb+f149/v1zqTCCscHzRsU3kTEYhAgDemGyLZg
26ln8rtckdds2Wrgw4et+RKMXhUgJ3nXcSyghch4O68VdIZW6LI5yuSAz02R9Rpr
tWEN/VH5Vj/m+Gnw8Ua92zyUC1C6iCHnv3LTgyYzwUJbReZgF5Zz4e3b0c1F6xeY
AfCEgJs8SYDRoSJNResp4NYxRM1QAW7evY14smx0lSYNeRGCPDtB5ualZXj0CNCe
t4op6rfAMu4J05sRK8qkmbft4/Go+rAC5i8MroVVfqtcYs7QaU7TGCAZV8hmHCV2
a4sCdMwybFrBlThyEIcc3zG5cICRhDhsdKEPmeWNZu31CBXBUPujb0A8jPBD6X3A
TYDspcQLeYU5nXqRQEnbpiNN8XFVPZhXCtCyguCan4X3gkYslAfPkALSTu6V5ura
TfIryyLn4S6NKJtwC1Y0ucRz88QWPpGEAWcr+SiCUfs/MhYLaiULgtYyaEbyfVd3
aZLMkmCdq+aoY/NAnJNPOsD+NQhcBufw1CQLI+IdYYxUE66XoRqVJUwiTLY3alfa
Mq+g0ooASMfZm/T+SLF7velnKMwRWxfMcoKFJW74SHM2QnknAElpKs94yNQe+T94
KQe/dCzmZxXicyLZg/Sx8XHonVuyxAvXuwgLK1s02z6VQZ6iQKXwnKw5PpsRxcS2
L9HLw1zUUuycKJ3U7EzjBU+PWYpUckfNnZEZ5Uija3X5JhcZXXsunS5RHQua4PGl
X40M8gjQp74Ykt5c/st+oBStFS7leFZYEfXYdsNBMo/AIwusXz6MIxxGpS8NYhlF
LgbZENh78qFKMZEcP6MnSbfcUEtyiVcQu/smrRkMXAjQBLCkEIJD1PaH1VJpXnD3
CVcNbBo6uqtayvjjHPYkWOkU4FEp7eq05a5P45yxf3+ePvdYbnM5JzQCni9ljiof
JHuXAKsTCon50WQI/VxxvhX1TEkeNNsTX7NDJb3rO2BZ4lATBw9noJlhzwZOkX4b
1+FpxHQQ284zINhhrLrJdPoIg2Rs2Ld9LEdJUqlmptN0jAaNuPCnwhEUBsOXkToZ
tip+7bqn+a8MG13qr8ti3+iMIIA49M3ME3WVCvRX6WoAHW4GOUd3Cl6AGpqu6Sa0
RK4MP0ryf3ajhOTvNz79m9R0qKvCVgjGevbOVmGPIcA6UV4JSCSVTd+Rncn/7XTI
8HsNS1Tg1fn0oAlIItFYLenpqYbrbU3IGNm8Gm0mF8WEb7q/NJMDcVAbHknfBWSz
gtdoEHADj2Hbeec7pDLOAYXru5MWBa4c4RcfJ3K0eoaiSXfUIBc4kUdA3Zk6KEnC
EUIxnv59ltozmj8555IT2WAzOJCSAQBYjRIeWn/jqeJdtXJJV5lPW9uPpbtklCGe
oHVyO/9sTPaOxWjMvmdkI8qS3VOQhEaD9j0n8iYOkO7BDVwb0JkmZUNA/x0Dfaez
NfUUaLzeUvetABVDoj++Opm7dZYznTbv7wP5bjfgTXy6pJaN2JZMFNnXtFJ6Bl9Q
hUw2/W+2UvfGjzbXIf2M4WR/jx7Fm19PuZMLJvqBAZqlepPojrC+KxVo5FCrAYxD
vUtncG23XnBYZyDTRjfGmZBrOYO/fPZSpZlVp4tQhVuxpkUNC7JctmkhxaolmArL
dEIMOYZwwcwE/r3NxnffcSENyjy8jTIiwaSRCJ8wfM10gjPgi+zKSRlwyRLkTtrj
AFhPMVlrHsdMpivFrpS82VVDlfrvj8giPrHhljDl4JtY6YCIeWelyrqEkxgYxxsQ
+hmejTRZqOZqp/Wk5Pvyr/S3FGSrb7baGSvQG37hldnUgt8zVtJTEa0gwnWqf7x2
WyhXVyrpY3uMUo2Xsnm8iHZu7RCnbl+tloyt6IubekJMK0W51I3/8LFBaYof7eLJ
IarTMn+cgWI4O/ghgVzmIu9xVEKx/lneAtBfs7vwfYktrRs/C2HI0REdorST3qXD
e0rDrCJLs2Zv4bKHLmX9u85n8jsouIXBLUofJRNIknJwuHdxiMffURe5YqIiUu1U
E5COknahpD7jIW/D7WU4PKS07cR+IbrmF/Jer/4TYSYYIzQQFclDWAk1UNCen3xA
Ngv2PGVaEhFjBk91ZHkKNzudGP1tePy0x/mTuqYo8wjAu8ZE2KMgAcLr3t+uv99h
8qzwaSrxMFZQ9bK4REd618htCOZXakuyahnvSFe9qruC4NJ8Vxh2W19mKZhrHHoe
xufdrjgVHdzdVgh97Af2vBpsmvylbN6pGYOENvScqyVqKyKzFuF4NETHopPSWFkS
WyNl+WtMkJlPl4bWE4jUl8zIlPkWm9DXmx9Zo88GYBz6VVSj+8I3lMZEWTxfrExS
iIVKeuFfS/tjtcuhjeltEdRxfLFojh8/etdyqP23AwQbc8OmrnsumhaKNr3A1MGy
UQkCNDP3t/xPJ5giRyTO1zox8bUPSV+mfIjj5NlXJMmC62Nq6sBB3BVapmjoEdo7
mpbr4u6IP8+ujQNMKoFkhsBcHZz2nWRDHwRMupRPQLSSHcNyHZftAl9NWoNvkrcj
X6ILZTvwziOO3K770vu1lreuxrML/eO7yBGBnE5VPnqY169Mt/l+gK4OsmWrlqTG
JmARh4I0LjYPXQpgGQJS4ru6k5uIeQ/jy4m4fJXrMK9o7OMrbPhr+vWjMYnKaJtO
EB5rdzuINykPXC8oA1g80lZa7ewbA8WsBsEWNsaU4e0uu4r0FwECXIyWlMT2WaAg
SkkaVIGpbJNbN4W8a7kaR6Ef5NXFPsHO2PyItxUOWXzZ6y4N/EHCnrYU0k8ndnHv
5PHp2ka52S+kSfm2ifHCXO8rgKijev+6LYLxybEE4LHh8ALCSdi+i4C+96EigIBu
dlE+MJL7e1PkCYrCox0cBEdSM2vDhoRoXHasqLBtIQ22J6MAzr75cpt2NiGrUzJO
ZYHo0CloF0tGxG1A/IS2rYPh3QoC13M17Au30+mV3CXuqrL40ywS3v9g+ZRPvUcB
YUsJ/OBAAgX09ciTKQOkcUKMpLSeX/5cFGHaOcp7Nmgo1+W+hA1jxJ7VO9Qf+Xzf
FSXGPW9AKWd/h0KYg/CU348RyLRhn2RJN98mBEbQybqir8ieSe0WUF0UG28RZnPq
yutlEEkCQXNRqkWvRxVg322RGG63qZ3QR0QLolWIsNhlqkrIKW4ETt300rnUgvTy
MEdwiJ/fMv73Vat9835hjZNDxSEhBARMafemUBTS/5NTKNvNYd2/aKfLZUbX1rm5
4lGeJKJyDXzRPaOTDp9TaQddhmHYTlngPxeBu5PG+yCGLx9Q+1g7gA4PoB/J3Udp
eztooC7YjVlUxhRbUNEcvApanxY28lHMurcz8Tt6OXxP5GVzC2KEPRoxwtfdjMRE
PcawYlpGljEjbjBCLWnPt0t2yj/eENP5rRN6U1pPJlAkkTYfa6HPAyigEmNBdbGA
fJLDXVhDzwpd4TK0Z+tMjoRU/RRS3nhZa9wAB+fZbi3/76O2OvHNM1v3F8HdV3qY
jPuHznxwKuLrg1zixDgmElVYaPr7VMxRvdEvuFx8Rlk9avhE/AkGhKrC7JKCNYRm
2dauglOfygoTqSr0yRuqigkvf3uKhlpmz79ZmzukB1yiYf9GJSQz78Q+kkB+ZL9+
IIMq2jLrOFWsbCMWaT+DhIUyjqQP6JIFrICwPqJPRT22urohZy+bvNycs1oAcc9L
eti2xLWNdK8wuOriwYLobTJFGaoTnp5nIU21RqavVRK43l3PnVOJtJZaRSUwfZ5w
Vt8k+GxC3Zw6SIfp6f6dGI3PXiXZXDC6MVAHO/cpw3Bbjw1BjKK4m3uOUyFTlOS0
HsaqKca6YmJJyls/xNmZmn6cIYxflEyh4sOAYyPNHuLtYNo85rZ3DxdV9NlBDVD2
y0lM5sBhZtHhq5aK6/UJpvVVGPSVXGaFvopiCAUMj4GazcMHJocNgb5CvowUzLYx
j63jZUyNSHQwkzcHifHCksafKw8ZVHkXSnt+eV3ckbVCLNLVntaXGtaIYbInL5JK
lqi7Vslz7U1eDNqmO7sat7M8S3xFfEAtr6Rl/fYYcvWVc9hlLwxCUxHCZ5GLfEJa
os3l6Fu2c5b9GIKLcJO+fyGhCfTY26PYxM2WVvth/5TLVSXwkHfhXKfVkxwkUISF
4GTdr2mEunUgZPPc2fSjVhPgj3AieGYjGFGSns2RpUGEN9oJ94XSECSPE6LPPAwD
pBzyTW0YGydOBFEjC0toq9S47bIMQnVCE6hwpeHKoLlgdaOCQlUQ9g7b6nvbcGNY
kuECzzGRdVttTi6iOoVFofpQUI/hwwrECeEho5XZgAmcloKRZoBT+bu1FSs453ck
OGam/0PIMZ/KzejrotW1GJ3IAUbMhB4hMB9hU6CDjfv4MEck2cCHhHQcDjYfl4tl
dmGaC0zY6TJ7i0joyCJ2w8wM3nRg3dI9PsoH8tGP0fWsgLjadxhKneJIJgssLjg1
eFaFhZBtwPSe6D6NtS0SYEmHM3+Gm5ABRd1huDEudZUCuhziw+98L5Obs1b9uW8W
My1Au1t/Tn7e7QW70G8jOxRke1UvhaPMMWv5tFXywiOGBPewSn1XuxIJjrAbXB99
RdxbiQR9//wNtxosC8MvPRdv8FNnre31h29td9tKNNfA2TfOg9ctyDZNmWvUejDi
4AG8ZNCX4PEIgMFNexNhgHaaW6eHl3F5mmlHOiTNez1rkwEQ0VKJZxZzlNe5zvEb
wHSGag3bQkbzmBMeovmuxD6FqmIgk3cyU89dAacUYJ3mtpjmVrmmZPYiO8b0938q
Yet2XWabT4EbLgR1u7G/z1Lw1NC2zNJwwBnmKTR4hKBuxbHnchbM9SuHFjWOAoEi
ihvjeMRlelVAtkSvctg7wC6THXtRDe/FteWDTRXiI5XgxFexZk5w/zpVFqS50vWr
3gUYjV4C+5mhtUHMtB1ctmn/e6b087/dQSoCK8MzZihGEDgd70nKa4DbXqGY4FUO
LASDDEbIPXtO8C+48Yi6EyKNc1y1mB+lgnWOZDbxdU/b7uJRMWYxBAmAToRZAYlB
DUtEfPg19fnKaNoRn/bG+LeaXNvcgAmVhloY5SYruHpU3GKaNGiN4UX35p5mTSpS
mN22C0IZuJahy0RgIVJZajllZX0f1kW1DRtlFWbF4d2HIlNqe71x5OnYgADDDFYL
M0Xlxlt5xY1L6IGhNrnACUxnxSrQfsjeCmR/bQokpv6aQwaB8xEllGD1bJvgd8ao
uOk4rtrAsbnlpKiYOuRpJhsWULP7ZkkPy6Y6hD7LSpZCzphInUDHFombzHLSWcTD
YwHJeEeABK8mgSLqEY6L8zi3xbeGil7HU3yve4tGrFIskX4hZ7NwFqrVAduoApDE
mJRIVabTrQ3JM9G1bN5NGkNXqIBK7yrH5XGiCw2Ne1nxyCHslVlI1De5ZXTfp4CA
dbIsS9LEfwv/YAP7ugeWWfNN9v3YwideuJWmXGBo0hTSVlBUWIc5mkKZY4wzUclL
7jMWmU/sIim8KDfqEWxhQ0XTrBu8JfArm7x9DGJBnP7vedPcEvfnGRgtlAoFcbHc
c60jxUYuaAv82RguIf3U4Zt7r3lvV2s1d1uBzrJxpszE/AqpqIDkEE+3o7dWPtPF
rCra3qd0sCwS3kqtcvX4HrS8As/73jc57XcaMU/VkCe9/mupMLBm/SRpD+XE7OIW
a9VD7HkaoBKyH6FuCQjQemhPY+jSwZ3GJNM0A8huMXdm8odxJS6JUyqIAWTOwj+P
iS+YvNeRF3VaI9dhALKMEJ2QyD1l7Xxb9LB86LDRegS35KKqx2I/blGauqCqC6Es
/8KsRQib06cADl3Mdb7h2pxGwvFB4M5A5wH2NXhn2pTUZHtNt9yXJ8jQ3lgY83nk
6lalm9CjzVyLhj11eVglJfzzwt3DtUB16Y4ADeoS4CaKK36mS04sFj3BeJMCwdJ4
zSsMr+6eDjDmQAPcYkPdfE0EllezTxebcm9chcQyIHrxUGO1bRF0r2bNJHlGYSZl
JXohJ+eaaIAz6OMRwhMzmW6y9UssXvIwUDqTwa+c3hc8b4DG7z+gLF+4YlUGZzKM
/lzVX/I8FPB+KM4aG4H5hvtoq6FsUbraA0C8AxQbZmCxj52vBtQif9RbWm0H14D0
cowVID8YhnRXZBwB3CMbn2FYrJZoDK/rHaFfG6CevxTrOsZZQ0tJV2E79qeMiErl
S2i5LkODuaMCH1fnoEAoJZr4+aSgg90NmA4/ozCVBiwICItF5baSt7VzOQ/vIitq
snFTaymAPvz5VGc/ZucbwwdjsXwval74Hqr0MpFG5iwgvxPD2Ittl2KKCl0W9em5
Q7owsc9CPeAHj4BQMWB75y8Iwb4hyNutaAgdUM2RJR7JD+rVQUcTNkxeptCm4YTa
fiVwhjf7GQSl7QekMvEwq/xunjhnvOi+wwI1iGmb0jiMf/rHxOT8H8tC5gq2+Nls
kPLu+5q01D5/nf8on4Zkcu6jXN7cAFNyU2w8/AmIVQh1is5QT9nJbbA/lkIVpnMA
HRUgFdBgZkDb/5km7YbEwZVHNqY8raPowRBYTsq2terlRc9rsUedw3zPJ9ewtm8V
X/N2Mael5pUN/qg/gjjpJ/twvOaGRKBm2rLw9vsFzbZMK2cqaFfvzdEt8Cg5smBE
eZZeUCedQrGoPuTdl5WQ4xMmZlksoHiJjcSrlcwLaucig/eVoaNrqB0bg3hKFvp4
BMmlvHIyDLKijv16RCgUP4fo+WKWDRTMMbhuWCydxf+tPOfCLmsZTEOyPjCyuPf8
NhI1FH6TqZhkJpR8ZOlpAGM2RWhTgrUWadN7OYAzv3n5pfhXzzYLH93S5nXEPoNC
7szJo8e5vnnWaMObT8+eaweF5Eltv9y2GzYguRhhqLdt+UaeXzbNNiYDv6CD3sT8
4d6PM7nNpWPB4tXPV7evhyV6bZbIPlXLN5yCuwMbSwcwV5KaNFnm/fXSDpTcxxXN
ik/TnIRlZPC+Q7eGTQeyGuW6n+LdeSR7c+67ZZArwlBk3WI4vgF6c0Fl9MbcoUJM
Nw2iGgO8sCzIErhaD4JkRsy1txZKPqnR4lEteutOpI9Eygo2iBwGgME8oK8e3DKq
uAjEE+ru7/E+AO1wmiDnA8KnIfI17kbdCq+pBBZGF4MoS6nlREenCLW0AkbHCNoJ
VLWCGnXP5qSM7LQDY9WIvaLKosEXe3zDYTHRvjM9sFPFo7FkvLykmvrerqLe3xHN
z6iYbpVzmR5mTymhyjSFN6INLjBzNQxSNwRBFHYZINzahPenP9TdShk2WMAhWytT
8yw7qe61usRksrJgGFQ8BeXQ0EuKA0tpGocHmTbz0sttudJyjNtuUwGXICz3blQG
LldnXzgzLAWMHgwJxI688zqcE1RV5+r0deQy0OPF2lCOiMGfPoMJdB/MX5T/ec3c
tZvkeultAYuneVQRdoRAXLIx7UJJgvdHdqMBjD5p+lLJ0OBqcviR5w7U6ExPVDZj
Cqt5kB6GmtVTelAleoSodQb3HKSSqDhrmqzzzHbkO9T4oVODdIOenEMvIDuzk7ad
sJniODoEvZauVKbvSVna8RnT+koV1ZXcJ0oa1OHQz+bSZsyJ+cMxasOqVSpIRxFr
1FuL/BHUqkEFIwI+MObu6oAgY7PTdAaNCtvXqkuvCplIwZ1AO1iQ17ov+47WrWHm
fknBW57jB8JF6KMrQ1Hwf7D6x8jjVoHvRSr2PWTe6TC3nG6PEZHWnRXQSD0zpUr6
xYFUj6jROJdAV17spigVD3M7Ns8WpskVzlLXsqmawWC9P9psnxz1Pa3f2p00Fpqi
ARu0q0mDqMlU80zDHFR2YuS/L0kjK5B5U1gatMgccTDKjE6qrQ5HMjjzAiE1kPre
lehCfA02I6wTD0yRyaDzlccW/s3lRCgrFmELI+w9A/eVc0H+HDQsWXe6E8Vg9gDX
okv4TB0BQOHDKA0H/MwD4yNqSzIDZxapYljkdusbopH1fRn5SFzV1ZDujbQrH20f
RrC5ryFjFxvfhAjL/29N9FP9fVOXAmdd2UkYnydy8wIlEvNNsSKmLGgJJNusdBeM
3VRIvaN7k5maTwA8H8wJBI0h+OZg644wZLrtOHAao+wvbrWdI1vt+Y18aw5aLuZS
v1PH64PcBIIoPM9EG8jb/Xzh/v+DgbQVuJ8U6AFaGUG/Rd6ZZ1a/HOn1+myZaeOS
WN0O8tQgM2pCQCQY77GooSyWN406EEGytFJpJeWoiCaR2nUhWhCWq8qL9+Q1FPXH
4CeGBvQLU5TnQLhHUtsAmC9/uE2jULSxiz9YDrKD1Yk0B/dYyNrYv5tulC7Tzpk1
K+wOatS2wPlV1TmKbCOqnOrTm+Q/lxBwGsc0uhoHzT4o3cpRirk86M9ADKp5x0hq
v2Kdf37orJClQpCcpkXJpDqNqFXPMQIFN9ub8fTZ76tAlbvcr76PW2bbfWSbKvHH
0vg8RH8jLxChU35dp5sI+WmlzlDUlmlEElyNSuvUxliHwvlnVcvXpf0KZbpTJaT9
h4FbEsP1wzuAYTWRDhT3o1oKWgjYRL57Ol+gix6Myul8BgraaAdSEJsMbTH0AlVB
jSrFU20LmMP4Zlgaer68CCj9YJGS6A8EXb2F3EZBtHSnURtNjebkuVAzTYhqY+AP
Qac7iWX7NSI/vrQbb9ceuHLIfuhVdLJUqisU1L5EDrPwq4ebmIblPTUISVZwo7Px
Td415WXpv5y2UsNckMq3ZYgz8wikUY96A0v1sCFU0JUzMqak9FaARysN/2YmTBES
l61lSdLk/Bw3DR9hhv3VVUSGZRBZPM5uUCdj0VPGB9EY/m6/U8cZzOP/rmdnYube
/v55q41qMWfMJgJ4hVZ+FOr84ylLZ5EH1ke0fRIqquHhPiq2XRmPwJcQiMeHBQWP
p6SYy6WHRSPzbNELnrNvSQU0qg4nvwdroXkfEnMJT3u3ruQo4w5E+7OtlAcNu4iI
OXgmtoGFMj/4v9pGDovDZmvn89IKlbIExFdd+HdnaMtLrboflPUFwE8/G8BnOg8+
v08KmYxzf7N9RY64GW809jBLJNzjnK12k6+BcnxQnMlPmgWsvQMCy3YDImiQ54GT
69k4Phm0cswDHf1SPSFD+B/gCU06y6ywSR5UbtGDPT8n16PZtWrh2rCs65At2i5O
y7k12l/WeBRavAVcrtVHyVvRdyxIoRkpb/U1bdMN+MzSVlvV2zzrmqwgX8MHKV8P
bTuBevRUQY17P+1i7asyilkWOtkDnfQ4N8z0Wj/wOLWUXDEoiIDE+VwaAQOL7nTB
CiRuZMqVwH6xsCmwvpgGjAlV7DWhmAG2REqk4NkTeg7TDJq/2l9OkzDYd+fhwcTe
4Vm2mtlUyKWda32RfH2+VWzMFAgA9XxrBnyWww/c0gJO0tUsnNviw2fFHsF0+YJ+
kjZPCSXZZIyOcWMlTMSuXFCvFsgxg7ebk6yEX52afT7nTcFdl4EIDCqPmgR5bpT+
ATNhLBrE6lg1OWS2TMltihyBA1UDZz0BdStJFAJdqppjO0Tvh4MD3jjfILkvFGLM
rA2fm56UgcupSCFaGWzEcyOPXnnyL9H8EqKYuwpLH2U5NCu08oLo5prle5UpTosM
wmCAOJx+vQ2m9G6h1NIzE912uLBTCU7xQOjweHilzxb34RNT6j6+wfd1zzRRyX4K
haM85senOa/oK/04trLdLZmhyDNDsH9ryhH6njY/4OjgAmG6Y2r3x4A2wiAwcnWI
9Y8JSZXlqOVABzzgJBPCvIk2PJf2hinnpA9qhdHkinViw3NUIvXHCu2/34aE2vbb
OqJi2iYRFf58lzglG20oKB/f6agPS+IqpAdRAkVqaLszDFi/U6i1CuQ9IIbW6dJl
1drs1wL14SnwvKtncvy9sy/AOGxi5qJHqXjRi/lDf7pGp6I3V7kraAJEEunVpC9+
txwdbe4lsd2nX5j7/+7unsURufiXXn0/ubRJHn68lqvCW5WnpVUoz8U5SneEHUxV
wvfQvjJOoG1qQRvMWkKxfgbQ45Dk0JWO57uzElrVz5EB/RpSYOsJlJRpyjZxg8E2
g5c67CSY2v9/MRyOs1TgcEGyWIoL4RZpjqiKiUuT2zZQuBopMWXWG3UtSFt1drmU
fKl03ied2pFKHTfSl/H74bDPqqBaYisjqrCeuIn8IbaIW4gjvapyHSvaUI6Q6/iX
WaNggo0k+NlHvqbCBIfReoaWKq+juyrlcw9O4X8hGIPfQNPIzKD5GU98WJjLgaL+
IffBYpF0R5nH+HwrINsZn9tQnearwn1GckJ7/0rkz/D+3voLH+D78HBMhpsaAM9j
rMCXV0inlfzcjBYUcg0i+IQzUr9smQliuw2Q0aDSotlOeQG3k468Kp0wxYIbnPN5
A3grxcAk1OyPxcKWnsWcl+SnQjBNtE2XSBY+9RoqPd7wYI9+VQbYRdRYXbD93/tC
G2vqkV1cR4WiLt3AgveOSSMp2hNZMmSUNvjx2zzNU03hbbiiRejbCYJohN04rUwu
J8OI0EyJyzKwSYNrnBMfZeol4hY9YwWvIc71Vi4k6rsYeehxu77Xff0cq5r0aCwy
aMOJ7zehQLNX4XsQvoN58iwZSMMLkEQMNTBe3ytmVrZDudj6DSkIZgWQMmvZs/uQ
E1sNU6hz010MbI/TQcVKaF0yhvNo4erYpeDguI4DH/yREidpg7l0eQztpNcFw+kx
yo9sQFvxiP/pgLCxXTf3mvicvUIIYBzA45N+F5/droktti7c3KDd6mNup2Hw7BkW
Yu+rYiu6dycTcLhP0ThBnnxBEhmq+DKC1WRLqIbywz25Nv5fG1pXPxdalLAQrGjL
xmHRpdbv+tc5hHTJlzc02lUYr/exOLE4CdPzypUnEwjEpXylr2H95/Hc8sRJ8gDF
3KE4doPR8c6OU01iWOUw00fHUVs1DbhAjGtkLj2gg5qSaqzfslMGte5WaKdE2gig
+oY702iVZFKKPePFQBDQPs0Ez2QcqofGbUu3EbGu8Erg1/SDunfm+UvG3GxUNaCR
lpUBRWpLXjXY/Vt7Blq1E5ntX10UT7czlyYXLnTWeN1TA6xiOo1YivwiwM26+Jti
BmlkYO+E4tsH2lET9gG/5WIz29nBdHc5y2FuDbG9AfZXORRyFxwnNWfnblAdCE31
BGxNoryDIoaT5+Anl3TLa7rveHLSgNbTv12aKKrROmosIabbO039VFkCSZ30cv7O
QFGjJzTF2Psw0Y8Kh7butjxVy/gSjJ4wnHBLG4GSBk+sbHXlem5X7oTyHZSdWXkw
9blOwVbu1FU3qOXaUSp6PTKTDmkp/aj6cb68RanKP8tA1g0eevCu9lmQn+4lOBTs
DhZnTsCAHzhx3B1D/aU5oNYjLewg/5bh/jGeF3OEGtjSyqVqDwqVqu22w56bqSJj
+e8ngz91dvHE8uwEezxu8SMi7LSoeYbb7ruzi91ullG61vapDPAFlx8F4UDl+dNV
idO7pkjIAuFPU/htAc56shBBEITcv5ccviMv4cn78i5xmEGCYpGe6E1sOOq7Bnm0
ZyDtq6TSdCwzD4zNaivlKO8TM5GZqKSjpmlPNUf1jhwbZZ7h0goNIJSdp+n1qCXM
h0luMMy9KsrjUeyWItQQH7rpSmi4RNFidSLlb4/A6hVr/oua8bolDP2nOgtAhaNs
EMTeUqgL1rIFjMZJ9CUsCyoG3BsIjAZz6ZxGQBEgslaIo3Pev5RPm+0fu4nepMhf
V41ayO4zMuOQxiEE4Gme/At22kWbhm+VCC9nr/OwraypA+7+eH/sLlu1xQWGs0aC
ZRnVZf5Jv05VwIX2KrnGh7XZJbj8Vdln6VRXOHlEGYOvxk2GrXdI5ugpBk359Ady
nBz/a4REUyBCgi4wI3Sv2jyyRQ1xMx1TH0+R0vBVDR2EkEqbLb59O0rVGscy12E/
5lbZjlML8XzqZ7NOQrsxHRxyjcD6lIWT89g7y12V9A4Xa/3pbabc+yIa3ShF8ARS
a3216a/oe9FN8G3Ar49B9lW9G3ZHCexMd5/jpkCe86l8wUsJdUfP84dhpMAdizCJ
AZhMq9KDr3TvHToHot/1DWXO3nZZXzFY0HeGDbnF6w8jkewyBZFM26wWkj5JAW3y
HlysZAz5pGrR8d6/nqzEvj1ibbzapP6lT4MnMaYT/fh1JxGH6xRD3uLoPi0PxMc8
MpAkYOdJ4/G7bpghAswNQHLmwWMe5nUV1lHEZ2Vi/SGvV5aVeQ2vQU9dL4S3J6QN
8X0ssaXA2kqflZseSHQG+wlpJMUZBR0mLkgJM7uugp1O9get55uVd0z1Fz/+MzqE
3jc5bi4vut0xmVsQPFXTV7zP5z37ssEbnDb9HKVsw9PjDRn4UEchzTjozJeGS0Wr
cpCz9YNnf7ZQJ/ivDs2VslrBz0FDsLY68HHqFMkzLoE02rI3FzsO3HQuFxPi7FZW
lG8H6c4Njr718DaohknEDBmeBotZKqpo4XLTd+KAqBQy3oSwfUh9u2YLod4UikKg
/Z5AmXXA8S3vArmG3Kt/BvUC/LD5ltNlTnpVxpAPf9Rkf9srqXrjVOeG9AufJzAf
4qvy4XWOB6KZZpvY37qVFC8flsNS0By/0PTlf6tiXljUmnCQLqmwlvyo0NWkMuwm
NcdXIcFt4GMOfNBu8qJ4tClxKrkc6jfsD+kHYgUTW1D9Rcpeu/I3QrmzvtRx7jG3
S9jKnnyk9UaeBJIEpvrIhJqYpeN0vc/xwGJicHNk5HYZCmmVIcNjUs1pKVcusz3x
pxwRqxFpULKOQwZA/j9fX+9gqVK66rcoVdASyxFPk8NK4lLQoTtxUlwMl1Ggbi42
oByGdxtdjGd/wrg33pqFdf2Y2L2PHZ1yCYMJaB0dZUl4T7A842wtuae+FEVh/+VA
lsSUbiZmT3c8VwEaJwZUXldiIQcgFR/BopYANY2jf2ig/5/YdJ/bKpK42EReGxOK
ia3oTUnwehPIy316YnAubWWXxSO7TUCp5oyH0T10Uno8DjFDLdrbf6wT7CKPaxc8
zaE8QI2aG+PkNilE6N9at+LKTcWvMe7EDrHJX8HIyszxmb5FqYHJhqOaupCNebh9
HArgFDm/UL8ooB2Jb9pP0ZLP/Ga9IZJ1lVZWLsspzVILd3LVXiI5bpj6BoqXMMbI
iLy6+eilSIS8KT2kklqkqw3qIXMsG41E1k2zD1cJQAJRxU1VLGomgP+k1HqHwRF8
I5ZJpN16mYJ4cf8fH29Q9T3Hl0jqpbqX9TEicAF2B/IdVo46EQL+LxS2GUZKbfw3
3Z7Uem0MzTIgO7yiVAryS0qyjtAWFVTq7Cv8cJHUWsqNxp7fud21Xx6w8nzHkYhg
Lg90NVeOaSK6MhiPbbEHSEqHbRUuK+/RmVAKny6q5VF6sxhNfMq4LZ8sECK4wvht
pQwkdDGI0XzdtRnUxfPtt+VFd1z0tnOounJs8pyw1Lj4N57Qwtx2n1M0Gau8PAaa
ju+fwpY1Cq1jZFqBplfM94fthrKgg0DCROsiEc+NAhfxwgvOaQq+zoEuH/An7Yt8
vu2HC3ibXoCIcOMILecemGXld1YeQYLrqmahG6AInlMv83v1kaF51dz/EFzwRXz/
KEmprl36d3Kpaed+4kXVA4dY4s9bK5MwO/+csVGI8htu8VhefsVILX/0RGnLsLWs
BKGlFLPGRmC/sWQnhBenubGY5WX0QiCX6/xtVCHF0JfqczlYctXj401KkPtmTjUi
xFBEn1vi4SwuZi/sMT5X3YLjy8+HEFK+XCnY7wh1/lszDYSuiPfvuSzp7pobfPmS
8jRSSn4PSz6ugshPGnsVnOBaMWt03GkBXs5gTektYW9jm7XIEmAx2NHUyoa1hKJj
KEiXJJc2OrWVqsWHqSAltHxMRvfic1UZg5A1H1oWhPuxcOe2sr+PJdhjSOqN4IK0
5rqBfxvaEnjMgLbeC3xuq1H5RjbLazecGmVUZwvbTOjCNNQVVnEuzzol6bnlrHcu
Y8PgMcqboO1g8dmMsK0BbWJtRCXq0TZpelVMffS8WqBtXn1FJf/oygHzgOuCJLqw
/BQ6Vkb9j9wCvwmhnA16bwuwtWnxjXBpyt/nPXJReEdl8M7omgRGVyIQQO4R3YvL
cRQtAvCt2Dp9tsP0MlAs32PbzFZG3jP3N5gkQvOZapT1yp6UV216hi4T5IiLaIS/
gdAZwEUpZJkMd22ZiB3B2B5psstz7lne0BOAYPnZrkePT5x7CkvLi24k1mlRqGN2
G5c0ad2fuJ7D//KH8aTueGe7FNb/AQGi61kswZ/qUZfJIxwawYpiVpuklTONWLDz
1e/JdEMTuRpr1Bt2QG4J2xXYkIgqaYxGn1zHrivOz6BZJYl+Embxco+91T2BQ7/3
fk26yu5Wx4URRZ28ONzPDsdoZAkA2Qm+9AKjRiIstYaEyA5xdLubFHvcKG2RcCw4
Hhs7K1dueOiBkv4dtfg7v5zhOfIKmbLVc6CEQHUy2AjaChDxopWk0/gzE5MLl27a
SvDXnyII+Pvb4/l26FmqwQTl5oOvzu4n8D5gq9OUx+7pfbLtCiUOLTj0CPy2iYSc
uXBbXK9TPMwPVO9Hvjumy+B2tYep5pFtptyuayszjXsPWnyh5V7GPP2zCaS5G+HM
spfpkFuOh13A1cu7Iz5+XiE3P3x5YvrVHQG1RuROGGuze7an4WCnWSX4OtgqMxWi
9O7+wShmYx665WLCSNyEf2/1D25nnI1uOelxZHVWK6U0IgYUzRLjZR4WrHvi6guN
+0KZiGb9An4FFmklMenMSA5BHJgHMPfuS8aZPbY8/yIkHwcWpUjI3ZLrgpjO0Iq2
cL9TX6JRxmTQ4UMP/wSNI2498mme838BTcYX8WEOusOhoklXp2r98fJcXQhJ8o9g
+FSHWDPYHNligjXvLIY+uQdPLkvtpaDocGQKVGlxbVRGrranoYgeferBzH4BazXQ
rRbsgxZ7G7o9DrGudRIrOwq6hAooGeqirW1/MFt4EFFyetU3hui1gyumwgSPk4YB
oRXpgzQdePO7ZkgElTzbSD1kJDi5NkCcQ1WPcwr7aHYJZYIT0TRcLfOVZHe++IeV
TpfI752q41WVIZ4yC/kNKwqZ8B8tcZH4lC/4o70UES/RQFiuLHZlQalmg9Sa4ePw
UkwndX2M7q16XNFcpoQn0TNwY4g4hc0Nc3Y7KTY4FaKLZQ87aJAjraOqZpODe4PV
YE2/wgxGkZjBbqNnKBbsTspqvlA8Xc9D9dSyvrApgWHXt/a8yQGztN7JokNo0kZM
ySEMGMQGRz1+0PA+/a3fII5Ky44gg/J4OgIstZGdoXPJFSpnog8OFM9X793BrcLn
MKR601uuLdpOUZUxsc2pstyFNR4L4ut2J9S+3Ngjr8MO9ASS+kZyGVYRaGYZOgb6
+ZCoSzHxn6t/jXUrbP74fqYzHQs+1OeQG/hW4/pQVuOHLHUa//Ga57+c3HV5x26x
WV1s2s8Lwsg+A5NE8k3Rs7DYLdA1hPS2ckqjXEWMhD4giu9nEaaNQCtgVJIGjbE0
1x3myJhdoz3aWR7DFkHP7Im3M8N7whYRZb1Y4KjFptmYLIWjpH4iHfrcZi0NEdt/
5mwTwgKzMeRXZUjwlvQ67lidOuJxp/rtuG4TquDdzESlJNUdX0mPFutLAvnkfElU
6dgu40PdP3Imo+Hy29/Fbp1g2Zm6l9KMAiBMcE8WLE7fILiBwJpHso+HHRbYv9Dr
93i92L8J8umqQchW9K5YIshj+AU1ZO17PlFB58Hc2n10GFkP2soDTDdUYe9BcRap
tfqg3fMUArTvjeyFNuAEMVTj+aWJG6LTbfS33v6AY+ri/d6LDT6d7EhonMIVu4LK
KbcT4P0MMrP7444tQlE4CQPKWm9SdztRhMkM6phKhTvcbVpvvMZD9zUkT4hWq/P1
yPVey6sftRAPD+kLj2BQyCbnUFK9nWhDyt86Oxdhve7E6yP54fpVFR5dSx5dXyOa
c7XXsNj6voHFL0UArS9tR5D2nN2NFq5hfh9266uYYVKw+mQdvRWlm8ExN16TWjLA
e6UYNGXB73YUgmZcjirqyEfl22R6owXSB+OkV2z5PUHjAitQAaqjhCz+mladWTOk
hWXi4qY+V1dWU86fvguOPtPHe1TeTYHbfJ5SMR/F/p4mHmTYSKsMDqC03D9G/J6+
hKdekxjT/yJCYU/Sz8lruv3CDBTLM6cZYaUDBgj83NFKXN0GQga0C/ap4dbkMsos
EsvOeI39/aeNzAPXvyfuCD9ZBf5czPyOs8qzA2roCN1L2/zt5k51RrE9wrpzfgxM
pL3z4yhSfB5uHHw1BCHz5fnqr9Qcb9Juh2UAaJJdM6P76nqVy+uvBTyZh3tf+d+R
Wgpg2O+hA7D53Xr0XITFWlwHXckLmeDikekosNh3kbva2brYagSKdujsir8udJQU
nekhe4kTG01lmWOIBbDKTc0vdeia32o5QYNyMCnf8yLEsyYMn8Dh2kZtkBpmNmYh
07OeL9h5/dT4/Knk+BAQJcHhwZgvaMTnVmEqhuhfJRz8oEblMlMQlyx2oSWfzSDc
G64y4boBMt0puDHarTfDLAifVjlc81mAo6hSMJfnzkaaWxfaIqzzH94kGF3hm7p4
vdpZ1AnultMYpxSKK+zy/T2GmRTttcsmhrDeXbdw15+PqLuIJN+wmZkkMek+5mvz
CivqAR2v1qLsa4Ag8sVwlBTVMU3OMTLWyE3UUA7rCkyJhqrPlWFKHeYDKdpPM9iP
xbbNeVv+/SsuP07W+eGJLSukbpJ4WBB+CXw96vXrwCeP3Y5WWo/C5Ilwaga/bPvN
XVfd7b1ssLn5qcgJT9z8mDo32hqqvsbH4FBTIlPfoxzw8lRvxGyk7pqaQNv5+Gp0
NfwALIMfunuWL4p3ByemmVTEF08ov8w0V3IUg3TZk5rN2AnQudEbsYlqXkAIJOMU
QvyUaQHlDjy8dC83Ct0UqjQBUsKQEnbDSNsAn5BwzwJXZSQZ6Vk2G9sJ9A8eR1lr
L2WP6YaPHSAgWNKuflXLEnBMPKFLUOGz43dI+LDJDsErcgQf+7A7SI4EBW3GaS6C
hLCDy3r5A70+KtrKhYlewi5XSWKPxZwmOrRftk/ojZfIX9cIgbBF912FB385+yxu
0Z2/S0cD4g7dXqEEXx1AmQ36oJZqimMhWGoF9en7QCTkGJ0GX2+Wik8hAxA/reEI
HXbGQGFHzaCmXntIhqy6WC2FM24O/S66cBVkHCBhF3J17UBEXiU08VyGH+hkXUkk
7EzBtSaNPm5EPEntLv0qVzFd5xWNQl79zz/xgK9R+JalT7xB1ARX9Q3UEG2TpWVL
N6H27/zz+E06yxr1tAijkG0SJBqSBM8tfvMgH1JgBP/MAId1t2hnn71ylxNzC9Bw
5QY7P4mK2RIcIgzsbp1ap4wBaNDYDr/v4Sv+pN63+oy3FDxgulMH2bceFsd8ctRX
Cj7xhvM2EX8xOtu23Fywm+rXvwG3IjYTyEA/ZlU9O/cZVDWIKy7jV6RvUyVTZdZD
7LmVqLWOP/jASBzWgSnOPlZuhQBMthnqMGyNE6AlVqOOVekCcLIr2uI+w6ubE9iD
+fR9mTvFDr42y9acRCjn3lVAFcskucQLtnV/fs7rt47geq4D9qbUiZ7FyvKf2kAw
0QPKDuoJu2tIbzsvWvaIhLioIXwxFf6QVFDttOIcdogv6O2rfkkiH27rxicMZrrg
3tzkC9ZW9EQ5zC8BQBL8WLdfrqy5VRGIYYgJU3dNuwEkdZrFKftPzGPMz8uA4XXw
9OUO2hiTgGY/oeAqc6caVoBDHcZAW7Yck55DB7qqFoe3+hUPZ6qnXMebpz22YtMH
Gf5Ts4KFYo53Yg+Y2WRSikK/ThLyTNoZjnH+GJxbyOPi/iKgX85DDbC2mKRHWLTL
UMAQ2pEpb7OR/HtkyIaWHsIN6MWMK6+ksZnsPyJGeZL05oq+YcW3O9gGpR3kTWuP
b/ucS6hJtvQUanBU6osoHE/WPhuydDGqld260wsNbApwcNlW83mfXGRvhdckkbDd
vhCLLHUYkhCeHF+8ZobrvC0YuQKQhhOKc6ybRfv9tChzpUnfxkHZvwtcWZE0e61w
nUeRi7HFM23Oaj9yBWCj1wVSQ69/oJ1V61PvCG1RVZxMdw6RgkjTh+pMAU0EM/C8
k2W9/FnhMJykKtxp54wN9FGG2p67MKwVGYPAcWdhPSo/uTooHtEs7sC1IgIQhQPk
68X7ZS/CgjI3yMyWF4RGsckdw8BD6qMMJXzWnRs5CCWG0SK4Z2cBch8yGnJVyeJ/
enNhg2AHOV7h8gQo8VlrT+xzLZI+Y0FDi1fSCJbSJHFXlW4HOqphmgp+S3Ltb5Sg
ClFBUKEp33/Tko3jjmT22qkEo8ulYyZEsrecSmluUXeSzcb2bBASWO9ovGTPfhO9
nZ8QCJfPI34cWk4dXWn6PlYuXJMjWqvLyR94yd6H5+MaPmhNSvNWLWvA95U96Pcm
CQFJpcSrDKRIwYhrCIrqd9/wvlILwwDfz2kPvYLCvGlNlZSFS9XA21QPsikgqakB
PJsgebbuEhfxy61ldvOmcbYWm6c/8cHBdkiudY4YpBZYnSdi5inPrg1BcgF4i2mQ
pkSCgeljgDSPGcmTtn5SOzZZwzntlVejcAXx6Dq7IDQVApfNWdZKGN6hFoaD2v6A
AdSbm3cvMtJmk5MRmrstSEQruOGAArp4KHfrLGOdN3otUueWcRifNsnrZhUPSkx2
Gs0u376rnBuNjozM1rQg5j4dujWD8y+S4ki9dLZmKUkgH+iw28xqINl29FrBiGms
X6KoGCTAOV9YTNcz30Rt2lRxHLlWww2UqtfNzppSWC8Z2O4c7v1eVQQ28zwp5AcG
El82yg5ylVjwJTJaJ79IulucR9oIxZsWNL3w9kgN+tQG/fJzqidHgWFVPzP+f+wJ
b1Io8BGYPZxF2v2snmg6yhhEMND3f5WOnNvob7I3DBZ6i7whI8UpZ3JhRjDO0FGB
OFuz+QN2CFHpUIbH5i1PG1U80K7j7Jg4/dyU/eZLmWFu3tPsTqILLkYKqUHeLkiq
Ezm88ey3TrG7khTbF8vHm00WjCTzgpr6fAoZWFIoVKszU7poC8T4sn1TRdD2GDc3
XYFY1StsDUOjTyRC1Ngou5ADCFwT+vP++S+SIngl2i/VhjbNXFlVvNufZnYRF1rM
rAHbhXxd0UtsRrKGAUEMpPkUlyZrjyTqTJMZtnjVmJVnLHBAhHYaBpL45khnQF0h
dHm5H0Xc/3kz7JORioXIcgQJjoEXgWPmWjrFThfiOQ/AXdE3MIttRp/CbtOYaxED
j3ZD8XFoiAsL313udzGYEyK9WZ7Eqc5DOl8x8itNCfAvPLiquvSieoSjiQe1dOA3
POqZdaTFsu5bSAtabUqsnWT328TFodFHkXISNkZBPA7jHRdd1y+MEqPg9SBwAzDl
a/dlPf1kiVKA+U5gSjsVeT9AznJRphsxAntYLXR+K298KS5fzw7cNqpuPp/wSTGq
9Fj2kM7MF9iptB6XlY3mO8FxtY8bUgdkmWgmmCBYHJq2fXiF0oFXEua4UbP4y1Ya
q+SJdtwnXrqdkIUX2OBE2bY86A/RPMvC1y4fD42Qqrr2n6MLFeeOB+lGaQlMooCx
ueL1FeQniunCAulZzznrMed8HOi7q7jB/TurOlYyvQuUtMK2vgOpHBNKVQvRdEjI
t/dHfCfLvkj5qKsBTJ5x8ZRUIQKO++6KVdDZdmcqHDXyDlR8jjVxbiuhwilq5IEf
sP2VEHC/V35Gc5A6SJpuOh6rwuyv6ccGPlcRYfcSymW6A1I8pfUqxM+gak5q4SnY
uymqXyeUAMq842kQGdROcc90hSX27eHLdUU4/+DeAhIPMit5KbWtWyd/1tRZAQ4t
pRLrCN4FKxl0Bvb93MQU1Mz8qLn+kwTF/KwNdP530kwCmD2ugAdQprNHUzxm/fGl
hgBXlfxkIffsD68Q6Xfileg3C3T79wLWZlNpz8Ie3BACXGFxpdY4r1r9uFheYk3s
HIBNvcX9k3O4odY95YjGerkUOckUEEdeOdvzbJo6aq2pdBM5N58LIR0hHERRDvUE
iBEoNg8MhvtDOYB9hewg0z3IV6rGlOdLEGCkt59Q6cwzT8hNAM4TPIbP7SVfONg4
vgwgoTXFHdc4PuXqmqZ+3Ghe8SIRX5Vc2wBjHUupZ63GzlCs1Pro/DpeaRq9U/3Y
9hWo7OTdGGO0uYI3QWkgZXj2ysPT4MUwAOrMPc5G+I7Jqrk/prcZuh+r2Y3x02Tw
5Gt01jfS1FYK7vaP04FEGi2z1yW7DCb5gUGuEqmXl2sTqL4t7mvLzy82Wc1It+G6
CmZAJYGZpUr6chVJMa1ywjztUOKGQQaFe8oP39f4a3F6HPNU/8+ObNJoZmM3ZgMS
8ZVl/dqJNnxb9Bj4Km1NPpdD/kcqjXguiMexMxPGSTa5IbjlFAphYIwH9zpZUaBa
U56XxKdm8n1QI/bVqzd+5mN800f/nYIy7gEG8GHFDeS3Mg04XYBQyL6twN5Do+ob
PKA4Vo7R+kOQp6Pggpo0YdbcCYFWmtp7U5t9/+xfgpNK07V/obWEcnL22QFWEp1d
tMC2kgC7hZVmge711ClPbRalmDjsDYuxyIGjekZJFXDFelxA4KaWQIfwJpTjtPfX
acmeLB+UNaTtqdECme7Yy40X15LVr/NCO2YOTGW5yNRJWSBl7SxDatE0wv+ZStAE
QHTgOpWE3R9RXI1zQmFf0+zE1vxHSBGB35zVVeuj8dqwWIlFzFZ9QN85zgDwVUZN
bJDYIuJxMLLcgv1NnyiigQ+pKA9voT/nU8V5dDY6/WJb4IRUxVjlckUbIvOa8xwG
9SXIBS0keKerThUqPWVCShlF3O1KojtLyv154DAtV8RN7Dk8DyTPuuqN8aqql7Q9
XLc1DaZCllT590Ce6aASpboB8dZpWxFtAIJoiGY5ZlRNOJg3oB/CC5qxDe2KDTbK
Zesi+VmrmIfIs2CLfjfZQ3WQU9uySFFkiYA/c03P7xrx4ftc2c/jDkKQpaxtZwS3
Xg0olRCZLHw3RIIbEmsMgX9QNKRkECFazcyNaaCs4W4ZVtG1YdBbJPCw2+CqippL
0f6Ccopq0omOnHZaRRR1K14ylO54UO4eWSeNFGJdfJKisfr+h3BJomor9SBoqjgK
abBwIo2zuqoicqhq2WsyIBwXsiRJF40j+0gZiatQYWOViUHxYXXfAA44LZyPVx8c
3Qqy3lGRLO2PREaJjhMOMg23DBYaut6psfuEWOiuS8QapAXyvYUUvMgq1UWmYUkw
kqUwIPYoG4DoDCKkE2g9T/Go6vx7m9jWcT3uqb93no1VEwYPbSCfNcPleUkAxHBZ
HKBRVgOr5NlDBmNdHkz1Fu1fofhqg2lNmLH3UcLcA905OBkSHQ0XnztZZiu4xmQH
z99O2PWNhAWzgEwwkPumZaq4jQvEkGTL16l0eQ9JCUddfQ2zFn15rCch86nISHOS
+nXA/nla0XZWepq2iMRK/QNY1PP2wl/Y392diNF4RE5sB/JYA8pnJ3QagbFP78aW
s22VmW++Pe8qSw4J2LP7c+MJfbI5sQHqhzxE2kMPryXmyDQTXgGT1dxtYtdIRVnl
Ey69WGQrDXNHm/taCCj09POl+UWyJ2vI5aWwWwyf0Og0AB4M+TWiWqWADnxYORC3
/9fp57mAGRxjdRF51PkkEeSNlJIHh9EpqR5UYhAppMKUu0y8y1m7Z8SyXarHAU+6
2yx+lTJUfWjmyKQiw2LCnPM9WQBtkCO8Z8Z2KOhbEVPXbs/5e2mfIx6oEVFK+poN
1yW8TBS6BW1KOiT0yQ1J4hwTlsWRj5Le+RHHvZF9pe6YdYqjoXFLt6O2TRVdr6Rn
6YSoGuv7IEp9mrJWP+u9gmOqGyN+RneTqnx1KIefmWpSgkfU2afZ6QxnNfGM1Tf7
PHzqnzDSwRj65/nEgrv4ttYyUs7DoDSLR88oU/HMbtwP+rpzumtRnHRlodSi/N+s
VdW5wd+jXBIDc30VQ+kmKoEqTnGKtKX1o15Yu9x9PGDIPKJmlAh86a/Hu68aSkmt
Zsk7/i9kUP4/4qpdWRJSCc/+EiA6VoBTKlVd3FUyFnNywQtwP9sf9b7Vkh5E/9LJ
pDEzKa+ugEoQLmSng5PLh8BySVDSx6o14mrB34BlUcYRKRgbdSiQ2ljytcVoG5xY
eI8T4RnL4Tp2XhHUtzgVAvpjSlailxfHzhawyNBBThb02JHhJGNz9QwlpxXQfQap
84uPpdhMghSF4jFQaHuh5gCB0CirRBhOA9jxsZ7NHGcutlezsf76KLc932RleZaZ
vqMc/EPvt8Wpa82zP4KUgBEtGoHK/7NbNJrp2Z0xZDdhL+0AVjBlqy8YhB3F1FbE
T4Cge4vVbPcLQPpK9aQhskfwk1mpHoGZxdOIoQSsXAyVIaAJRbBwkQwQX91fQaM3
fUe5NYeHEmidf8KUUdrnr5wOEuLzcQFybSHOjGffN0DG5iQJWtDLO1m/FQqRdo3i
FkZqs3DSHJ1X0yDY1uxgZuUQrM2k722wz/f4AC38tfiV3m0mEBDTqddfv+pqJMXp
7W8iUya0/N0Nrx9D8f4S1cqmlwwL1vQYqMwz5UEq0+Q9UsMGmmfUTBJN0P7pUeiO
iqSef9RZKCfOkt+MZsR9077XjExXIIQKlezHUO1jD2/Fh9Nc8ZAacY22gmZapiVq
aL93bvAvzzrbjib+wV7CLjLjr/xKxnHlqIe2fsZULFwLQ45DyOO0pql1Ad/XdHpg
+rLTzTZ0YKL3/ghc5CcHNZSkd7E0A9h0IbxItzy4ch13kZgJH/8Zz9wBCPIAHiXQ
Q7YA4JZ1pp7DS1KjuVyvGukgfd2HLFcyMhdeac7+kykgOB8AgcyjP++i7IgXaCqe
5TRT2XTGqagpT+x+cTKepXrODJYi54iXvcX0PR7Xllq4Sf7t43fQDxDR/WyjG9t3
ZYG2grBeKqWKe/r9+2yBqnnU4M7bWKja3jdwJnZv5xCgwjseyMX+ve9U6akWcWwo
U3MPgrjhM5JbFzTEblfD846i3yvLuAgkdX8gq7PqMQZm64TP0H/tSC3YhfqXnhHr
Ve5TYiw6qhpx0+z+bhcUppIyAJq85eeTOzTuy3qAeQMGBDnUVXCs+HDROdZALHzb
620q3I7lGPJ3HkcObkXEpuAY6pyjLU0AMkCpo5WvDTplqnUkeiEyv/KVeYKXCNtn
s8owwAs+9E7Ej7C3RrA6ZZz+evDKMgtemwtXN6VHfjJSzG2l7p3OQu/w3syMapGl
PURJrbds4eCDGwWqLpjeEkMoB6w7YeKGbKWxi9XP4EMlWZUZV1vrodfehZ5iDydQ
bKQTCuDgzMeEeMtUjhSiXMgt0pQhfT1m9wyFMoDdF9iSYuL6EdloZseRGlZf8ymv
yaxNx7uxABOGzgTKE1n/Zj+cLIxn/h8PJydtuStVP7XRRx2fEYJNgLW07uT3G63K
tmBT5Hs6PV1b7q5mH5/Tqxv+V9Jd0QG5ElX5OCJJUZnc3fFOwvB9S9gkBetzp6Pi
fOc9KOinSFTCvH+Z8gHl7vIQR8rjBtrqS1ea2AnGH52TOsbMMysiwIyfntV88mXV
Y5pVaUil+2cDX34ter3EE7eCAlsTmx3K5bk/zBY3+kAGLQ7FF+1gdpgthQL5SWT8
+5i+QNsIi6R3f6eapxdfMI4F6mBU5+LHtVFFrRXI4PVvgXB+uceZo/sm/gc2uF3A
hWYCNAn61p7SxlGbQN+6KeohrlvmBoGm9DPs8WyhzN44wYCzvkWQGHF0HUZEwfvE
PdXyqRgcck7CCaXMcjTeNce+S/QypGQZvdo5mI6CMp61zxEj/F3XVc2XMOtMLP94
JXASzE13HNLvM1QXhnjyYQTyAxZW21pXeZdHqmz8pbWIaJeBwveGyijP6VFFwdXK
L5d6syU7b/DQs6Euf6DeljALOH3YpXqOyK8khaO/4p1WQ4ADL5NQKvSAr3c6e42B
jCGzte5mxAVi6juKVa4RmCZyp8pgWpIWfP8QdFthRhDtjN69+x2t378MuKMoXea6
vaHku0hgQJ/TEA99b1910G282qISmWWSyl7MfYSswAlbC7liHQH74Xqw6OUpqlq5
GBJgQjxDF1DjWh/QOfhB4PUhtUzQtNJoVnhQDN9OPbLl8/97NeTpBqAfZr0vb9QN
Jnhm4Ynd39k6emmz+S3xrGqqk0K20oI3s23pDf/tOyR+OHDGm8hOL8FyzQ0IGLxW
9k5KmPcv4m5k3EYrFfS6BIw5swlgrm/jN5kh5c2GjfzC+Gs8fFCe8enmPUjRsIst
LUPOiF4g/snrMsbya3Nr+AfGD1OOagggnPCy+KTNr/t1EF3ai7oyuoW1r7VG+aA/
zQ9NcfRjubed+BjJijJd7K+QU4M43/VzNP7/G1GM82IOS4IGxQd44V4MgMiGkQ3S
mEWxWId7vFSO0OLWRan8CSFu041J7hmd8YonfR4vHDwgW0K/oWN9+3msyQUs0cWT
lzd1TnqLsBpA2CgM4UXFjoZsWRZf0AvSw+jJYsZjXFcmMSj7X8Tf3WNo5zIMUnwD
uO/UkllGREdBNfr8XcNNDP7dIaIdrsrVsAbWgAHsC3+gRGikOQf3MelUKN+ZaCS6
aEVMTSTXoWyjdwnMLO4uO8SDpBa9zwBTQhFeE0kcNk6QHVA8/QcFExJbfyQ1OY1m
3rNFYYFlyuNJrC4yLsYd4qh+ysTh5x3m8J8Aa8lVcRLWay5y3i5ti7gSE91W6rKv
MtqPksuGNkOWx1NAkZ8T1va84louM9Rexfg+fFGSiboSmMN71pSIDi7Cz5bYrNi7
unw2ZSiYYXNCn0/9FeLfQZ+TlllBDNc2qHNNjaGMnGRNrGLQDLxMnI6fTEwABL0I
PvRGYottvP9L7tArjtPo2xbjudwSIUciI+chkrGuePRbHd9Ef9th/Qbf5U0wHhQw
VqgKyEf2tVto3XxNQSWeadLfyYMVE7ti+VXZAE5rKBQSEz6hJfNErC2x0GwjEPPQ
Az4DRrnUGJhWcWBBUnVQKsJjVSN9ibMH/DJKLe5oDBycOpms/uARN8JmbEztAAlb
eEmikjUHRLa0cb09yQYDSZBgN7dJsKR/F9CcvDVKMCwvEshmN3bHfNVqSNY10XOg
Zheso9NP7YF7OGovyEpu74SHRGrdMrzbmltgG3Yx6j9NAzPDZSj4oz4c1tIa08CH
/pk4QRnO7d1ZWAGZKBKeqAiGWuhx4qqMfYyqxb4V74/rnuyfac9faG1GS3wvC8AG
SFqdC19bKSUZWJRD78MnVZAfu9b4Ib4vrNf9NPDFZeteYJz0NpYl3RhpCQzNbUS1
hRMIiGgSYEYAYKe6Ai+T5joOmF89tjSSBkU2SlbCLZtwI++kTlUjWItNlV8KnVzj
+4QAa/c5WCDXBAkT0MHGKRDSwD9O+hYfkTMeO01/frPUidtb/xMmpGjbma8vV0Bz
ujAnrjqNEa7eeN9XLXCy49jm7zNVYvOp/b4sMrM9FNoKFXcjh2DHe0ZHocxnnRCc
ffGNPjlxwzXE8bsdMmnEzrlM/pIRbTsXSfjvoizSSJBNS4+KtWoUU6PrPQEQgqDl
goTgcSWYjPEa9aoPe8fu07gQHs/X40vH9zM3ktl7I3KrXcDc71+ip33GAHbys/ew
bM99lFrkZLQOCjJKENxbmPSErn9YZwosEYR3wyG+0OEqB41IJmWychGo44HeGVgJ
DIJbdLGfMa1KlrHIPDgjrsyJUPmV4Wwa09stpdFIxCZaCasVjd82GyieUXd/RN2P
YwfPLNPTRRnVY6KLodVOOvn1ZNKQAO2d/1SYGcW0te/npVzWe58WxYVWdCfIf9NU
K/EJGwWitA3GHPYxul4HumjNkWuohPnIeoqSYa63/YC+KDTl7RJZwTwTeKpMiguU
yQvTasZdcQxV4MMr8hAkWAPLLRHqr77b/hfGVa1/QmMDwTe+oU2JKdTecpOHidSr
u1oENPBWsLC90M2mGD2iyRumQhs7BB1nFtCtip5yAFxl24MDQkY2XyrIWljsuojE
ygH64rDfi4YKO/cPj3HdVEI75w8FFvr1RCmskhrtIX7LQjjJtmX6bU9rWvX/ZMqD
j05LfVr11xMIQXIVfy4kax8eBylWJSUUDdot+X67syyPiOVGCJENMGmIz/ToAQop
h/10VleFFccbKoz5z4vht1vLb4f2nXrEoeaxL6Shi9i+jbecW5nU7nhwo9Jrj6mV
q4ySzl2te8wWJgEOdbgBs2DDaryj6cb4PPPSeGOZ+wdHjya1g0g4Dgb3V6fbKcXb
UaG+k8F+NeKarzwfTQlIZ5js4IwYuv+pz6xjSfahI/6X5xpOj0pLXRpLxw5/X7Dn
wUpXugL6LKlXexoOzJar5OTEGvXNhQXaInUasXquvr2+wWsmdYn8Lov8HtVRsRJv
1wScWjZfwj2t8ERM04UEbP5XfZwDi6KVFEBmpumZq1UKpYy2eUvnyVIuXGkAXsU5
fi6w/WRovwRkybmf0Tfdlp+EXgGkZ64aqa8oqlBCaKBH66rhCMn2SaxfYcNCCIEs
fIqwO9aPkuY8RHgI/qBYLrr6FrIslbMuWsW0KYGFVjkDFy06dCgVEn3AgC4F/5az
7eeaCv+7Q+9QvUwUAbqBDpuqMGMRauPQQnCC4Z2iLqx066y6C17oFS0p1hj0+bkQ
grPT2yScoZaW6ujk1lWDeC9PgoEvaV3CoS21KQV6i6e2VI2n6sWWRiDh7DKyaC7w
fRyLuWnCtn6L5By2PviMfEplu14vQqqkl/nTFGKUSOg1i2wTbTrsHOooQPRVH6bB
youo7otaVfIGjzz2LCS0pmYRRflq1xxvxuh0GphOa+Tc4aEIv8a2DhLEf3Skfanb
EhFDSDcHo87nG5VLnSR573JusBqZ8lFbKIwMuIGXqctb65jXZBZlciMKS6B4RZSB
VHSlvgh1KXOge1vEqRlDnJZzB4mALGO1s7NAwpvcyKtBqCFHxHCfWiis368RRGAk
AcHWOmIA+ZsTKipSUdGRFlrLuy2vMS7o8wg/gf1rarZRy/k/SEc7udyZXyeG2l5q
kkf39q4YeXhyqAOMpBq4VnbY1ZzjBwxop1S+jNPV2I6mXGN1cyz5iIIVwtaZCFZ0
we4PMlAdFc2ToWzppJ1e6dnDcaVrrAYhdFPUtvLVq6LrpGRSp2qR9N8RcmzjPyMO
dGxxjj/D5oyHGeZUD1HbuZ4ie1Kpq+8IZ01V3mu2RuL/TC2rH9PxnVHwqJwm3Bu+
VsFmZw4XLKZkkn7ukuJrYYQ1/uofOZbxBMW6XeXvEf+pqcIajXyW5a8u8TZOXOJd
585jPkgHNPi5pBSnPxmygNDiwpOQX8yOZJwuNk5wQyK34wPPLYABGET0U58lYihh
nkW0reyqVjUZyKAWzKqvmNfaeu41C8uFDRaeempcyWKRhkEIES0ylUcumSDMqcRm
dkVCjnuh8qBZXF0q6wNQ0pTUgcWuNFLKJinM3bXj03xC3FN19E69VrwsvvU8IGd0
0u+EbXDOHvCUZ2iFWLn07wbDh+aoVj4rg3I+bSpY/jV46+JaacRf1bLK57gH8uHQ
2Ggd3433bxSl/glzygO3BJGAa4hbcg7VhGumTmwZAi/ayFSsZMSGD4qht9o8UMrq
tMpLSIEJaCrtYivethcJs/mfUYFP2TFO3pvK/FhwG8v06kbU7hAbZNFNp5RgEZqd
JkTDZVf5rSnr4UKDhc0i2J6eJr/fbjVKPuXiBtZah/D/BehJ1wFEpa40UQV4rwZc
DDMO585X9pDZqcYcVTgHsjbCgYnz1af/1KR+MigXpsqeVrkeDr2syhisL+VekF/h
IOYdgXJJnIamPj7JkUSFf7B+g7KFnalX6y+UhUvlRzVuabSTwhpg74jfZn8Z4quw
3HwJlp3YJDR9DLaWUb5I8apIm2BFt2nQ0/sphQgSiVR01gYERfTyE5zaR+w2HZGa
wBTJlGZ7YqIZTLKsswc5R64I3w9KVd4QEn8OTX5V9TVKgmFTYeXv53eXRlU7sUib
TetkeEAX+TGvuBIMM/ZI+AL9k/HgYBOg5Iysh+6u0rm0/oqhx1vOQ5CkFIXfz59i
06j4oI2GDIepcBBss/JkLKltGACiIYw2BwEzHYRi9lSThaP1wt0opmUVIiqEpEBl
PlXXUEOLZuBVKVVRj5xGxol8ETe5WfJx3N1UD/OaxVlpaZlrcerJgneWEY3cgO7i
Jku00QpdsVXRVZnjtusZFJxO+qehOVAR6t3BZ0aES7V463ExU5tjEwBPF/FhIxup
PgbsIhPKAImNsVW78LYWb8E7qa9/rfPRxldjM2AuFRmMQE3yN5d663RvO9XUHASI
Feu0kekjrGBXoQlncj6A3bzzrWhg3HUUHlRMXiA1AShxwpRr0TeM4J37TZG0t8vx
R54hRj3xiG/BvI6K7j4p8206kh19MlxvXfEghAHf/a434CypF+0lZmoHozwFhYLG
BjPkKS8nLilmipKtJi1uswCE4lFQSblCf32HsYAktMcm23z/1NR3c59MCqowVCey
AZCX/6EklB1mwTZyD7Ht/3Rl2ppAMOJaqAo4ShQ6nwskYmR7+b7GcrEmDVKC0xhv
KVsZf8grtkvliLNQCagaEDYxEeoZFWOpKxQ8JKkHeGT84fT/mGmIj6ZtAETPJ/ci
GG0FXFtXldxcI/3w4YUR1JTyryUHtnWoWRwU60VMzoSXcOEtzupi57OG/WKn2UQA
1T26majPq7C8NjdH1vRNg5UjMSGVv2eCq88DBtjfMrH2hLzZY3HWqCcWBkmO7Ycv
TMXnaYltevX2/53J9oLM5PPQGi4tmWrqIBu3Y0T15JDl8T1X5SLqqeZXMEPuGizR
iVuOgTvBhfjDx/x0kcn3xGs3blTDbQ5qY9fwkmTvFMQvFlCtCzKjCSFaNXqC4BBR
p2+3y54b2bmUjTxjC4ALyK8us9/uPF+JMZGMhvp5HOy/ciV+ie9miNq52e5pxBnY
3rihMqBY0/xKjtC2KIvNA+o3N8tWsHeWYP3V0JFd6duTr0tE6SSgNGGW94ssDrN2
F1cfK99e/jHYBKvf4c4ihT2vh6Df9hJPm3e6om/dLOhEybP8qS6t+OdA3Yb4ZXvy
6dCq4WrooarlN0cya9CZ0SvHgshBIdy9iyUuvyHOChqL9H4rQqmQmPEYqBM4MJYx
3OcujeMBkvX7Wno5WY7yqiuHyr5HcSLL9OQyBJxc5xKjhhFZJc0zyOZGdDD7ZOp7
C5EkioqFxPhCxtCaLvv5+D28szY7RfIBYnNprkCzKdS0ZbeJqg3qKENe5JvcMtid
XeQch5pLc45X73Gh9e4JwcwpsdoKu8z2jJuXM8nBuUOYsh1dyEfv47pJp/BbzkuZ
fPfbMDvoKh0vrWpUjLGZd3OZZdoL5K1QDDv3XZJ3Qv5PblmtnZwMnSyBL1Ka2J2a
+DT4G+5yCbmuP/PNQOWEoxjzIDQXlnzXhwh6Q52x/iztgssbOUPz4giq8CHMS+ZI
80MGabyn9Ck1GuiZma2lyxmAPvOCseR+uU0Z8JrnwAsHToe32tJr3yTHSexQkQAX
sqnmr2axnQYHD7RwP94kyr1/7yU5xgOk/7hety5m9cRAr+KBlyZG9lScRM4LT5Z/
A0t6Iz/kAsOwXBm1wXhrjiAUVLTWv0gaPTipcUcXM0vIF7e/aL/616NZ/e1vxa1z
WvMnFemF4OLO9fd+3z+RBPrI9M/jsB5ZcPSNBz7Poas+NErUTDFFdSm4ukjIlGHm
uQfl5QHJe7r8eOFsiUFYi7gg0EI5CNrY1tTVRq5S/MyougetI9OBX20xeKeSWHX7
wDm/BlZpl9tLZZfVUwnHcmRwvx7qrLFOc2xMhedao4IuOPvYKe/leNX/x9+TOpdC
z+vqw38z24m18ZD8UNYek5zXrsY3aAUjheoXzrH5Bt3+6ZeSN/W+lQAIuWgnY7XG
7mAJf2DlYNgUD90zD7UcH2hwGyKzO2bq3fCYa0EJ+I762yGGtauKFW2EZ5Zul9Qb
fiUIdp3tF4LqKOfVfwTCkT5VKEDgkh3OaCWwI8zEr5+LR9knHLP9GUTzpFCQ1gIL
//K7PjWHMzYbqM/k9AWXMSW/KwGbeD2zrGqkpTJqKY4L6zW0vakox6zFY9NUZ43c
X7u5BhdiJMNHg82MjmHWn0pkSrhmJGWYftj0lwSPCOtQEDEJL/ZTGTGgBCgq4nDr
atyIDEV85cItp9eb/3QbHUS5oGOl2PgquHe4zRUQCSGM0rP7Fj6JQMmGL8tmnH9G
o8eB7VH3Uvu90p9wdeJqWyaKN6TppI+KhaT+FqMe7a1IwpMtSw2fGY2sDSWQerdb
yeI3Vu9hG2oLcwQZVfhsg9wMF78n18ooqRoNlX4q7RSw4GoA7fc6A2/V+kPHcFDJ
/f9rLWEEzMQ5hXUmStNKHmwwRY+Vlfv+0fG3ehdIQETqIL+wy+NIVcBWUCt3hQI/
vJFqN93SgcUojEIZrDn2jqEy+inPGDHCs/h6QvZT9o60CC1JVJvS3tA1YEtl8G2l
g5R0Ufw5pQ1yQrwv2zhBi85qlyAaE74b8ZFw9o2Dt9fL0lW0fPINCakJe0Hvo/VD
NP9wU6IVUDTz7zz2Hs/XEtJS3GcbbBnnV/UqpKNFSFleCMDO/MZNKgpxRfUQDdRG
BqhmUuPbVqcduGmOL8o9OdH/17L1RU/Vw9kOENUGT97rsG27GPypv67SpKIkXFJW
Tv8YdAL/ylXfrVq/wVy6a0BUBp8k0xs1isekQ/N9gjmtt5uf897kMNSHfZ+p4GWZ
a+OK0mEs76E5vADxCAHy3FWamzT207gYkbhy4Jwl6KUc05wdDbQxD5rQet0pcF9a
APuxFxsJJuIyUMDDtwbzNC5p9xMoyB1JT7ZQHDZvZfzCEQ868/Qi4BLmymlzntJU
m5kDPSQ9EBcTMISYBct6ud47mqj4/X+eaFI/z2ZjeGw7O+RzPQao26D2jIZXJ21q
7sLdOepu2K/aUdkl4AFUXPR6pM3MzoJEiv7ELR56KO7Fywm63dMs14vYnnLgH9Td
P8ROcim0eLE8eLYCIZerHKX1LveCUM4N7kQludPN9lUEp+dmUOjijK+aOVxuoHjJ
MN8IIk/vas4YkJIkBZmvSefOqhxlL9m+oldVJhGhxsd9HfKrEcZjgJajYQl912MT
hK5BletpXwHJR4GyEdNMEGwV3W+A9YN/Za01v6rT/FRHtYjXx1NwULHqEw18O4B+
NA/WksIhZcyCP49JNOt5bUxufw0jc9gFfCwPPFA2mXh9VUfXkgDOvju5W7Hm7biq
pDN9FsNLR1gj1aP5WJEMMg+opz12H/1CddkiLfHhzFtesP1eRLOyc5qvKMaGX8Nx
N+nEbtNhZwNSd4H8ujulgYJEjCTbGWRswH/eeE2GS8x3qFBauQkjKOX9fZ5pXKfh
vC8EeKXuZ9pOo0C1zuIm7UOl6M7l8elRwQQEAoDzNJZRjaRmt3RovNlCtpL1e+Dz
ARQWYNwUwMp7RS6vPFWI8H1HsN0A9cB8cyv+KtiSMHGQBUw0MJyTjy3s5Hei5e4r
XG4KE+KDRn2KjxkbiY0OL5oZP7j/ITNe9wU8wXbzBUMOzK9l8RjjywCl/AvQpXph
DcdS1ujV1n28K2AN+m3IXgUbTVlbHX149Cxx9kLStNDUWqSOpV1lczIpeBL3GGuL
M69czu0NHww+Z0gycTcftXAX33DVR/T2oDE19eeShj75VD/GzrNRXuThEnkwO1IL
OCOgiAvmKyOrfyHGuh/15h9YQjRW/re09Gg29zmlBBVmE9YtN68BkejZw80zXPze
FQqx3iNGSN6yHk1GMivdEB9NVuy3QA2BG20EiHmKIRHx1Qlpy/e/jxyinTdH0p2P
3aCOAYd9DTgFwny53llnuM65FsVLu1T+l7AA5JN4HIiWaPWq7N0dQ89zkleBXKcg
nHiITNLI7m8pBjbYEtOaR/ldFw16AD0QgRyqB5J2AZzsD0cvfgUFgC6vP29K1NU8
foOS5x9xQlZcVCvJ3AuPUuDsN7Se15HvZHMUwNONQ/THEI/uxHlSaUM9Pyc090CL
6bDhfsHw40udbUqxnM+wgaKnQvcBnsAN+GNdJ8Fe1G7wwEBzVDNFnmyzjGwKuaQ4
/gfotxftOua8C9GVUwDkrSgzewUeJuRk7CvdWAoLQGOlJhdIAoZ8xWnk3Y+R49oB
4zq6+D+z/lXSDIoNnoDqF2Q3Q8tJ/dTdKW9RnlktV4A4+W+6kzddI0LXZCvev23s
AvdT+8z+tW3bLYJTnMsAxm5Yz+4kF1nt0NI1sMwLvyXMqI/bwxWaROqScJFzInE3
NvvYpfV+yfPnhvuGexQZGzFJcsy3xLBAtiZbLfBy0ldQskuXyjGOk1YOHWk35MZ2
ExxKQruQjxlK4Z5mG1PZN7SvlKawfEzpZfQVjQ5TNP4UNZwYy3nDLm7QSmVEBoMu
OHTZgd13wVdTrlmVHOVKOBasxQ1AUIh+cglhK748gBGgjglM0nru+/8bEkDUGJdT
8I2ewCN7Ufnk/3DUE5f/8PIoeKSF1ELM2QeYDDsx+cQ5ThLF8xFUX8zwwmsLOy5K
9iSTIMdV8LCh4z0li+Dlt6G2gijK9vUmbnaVLN4KqZpWqRL1Mk7YstTMSbHraqdZ
WXi4tuNrNLV5XpnFkHmIcnJix9EO1GYZhhwyJZHzQY85VpvlwVYMX1AMmIOKDkgF
ir825BN7lnB+aTY9Myggiz19V6cyJoIaf6f+Olo92u+f2wUCwn6rfBfYicanPSD0
39H33Qmv5c6xt5cqiU6CDYDjqFxY41HbQD4XwjfL4AIwMuuJX/fZ0Qg2DOVEwjNq
fsfLk+XBtax4PxhGaR2OB/0nLGMID/Sz4ZHYZy5DZDYmPNvVXPdgssJigmpurZs/
3Qm/N6GvVD30HY/x3aPL6wHX2mjttQ1ibfCAL4dZHpvCGsTuaHhej6YfEkKpKjur
agajjHdZm8PoAgwWaSmULkH0nYK8I8GkCeZzF61/t77S+sYKLGCkTH1WUnQoY4Ty
QvJRWGr7i4upY0h1VbViY5gZliiWB1EaS8gdMcPPjjH4s8M4r5KPZrK5rn2XckFf
6+CQIkaETOz7/T8XXbZXXgX7YCoeSNXoGAD0P7olxfQ7mZKarlPquHyW7o8jVum5
sG0tbgu/PsQ9uvmwvuEjperGYjWrwVwPsjaM1QJFsFptgxQDEA2okx3BCGJCcDaM
oYaKhFJFv+jvg+Sk8Nt/QYn49jPyNn8BI1pFTWsj/fRoN4Y1BHKlap764g3pVmMk
ORYYvvQ+89VLHjqbCcr45Jetc/VBO3Q5mc8xpEVVcvpHlXnC/xHLycUtC3Yb8Z0x
fCmMfATfJpBCJ7S2DEbROhj5zRJ9HqAttKsu2jMOrWebcHw/DJp9iR/bbZT/b1Ry
FPURQ9g5fcJe4gY13jos721BS3WnHjwrUPVp0mGn16kMMjzJ1OVjN2dbj8U7HB7n
ktMKYSS+sDVUCx40/nuIRIlbZUbxY+wN9rFApAqGFDcb+EhR0EpCTC4OT7YyeK+8
Dnq93wSOcLP1XznQTkKB2uEmtGv21IIz0M42hIGphmy+4fyzqzrsITJQxiEubf7W
pUFVde3t9M5vYSWxIpROLd2+p5YGzcDE6PmtkQlE16EcymSyWYimIP5HULAofloy
w/27m9482R3crvUAWlg2Bf3/CznvfsVOxH4CJNTYRab5tiCAsI2vXxJdsNPfKfGD
uh/EeITQ4wC6rq6p2jhfSPnCYbkvkHeB67ozou4eSrR+AyWFBM+VWKxNKPTqn1Un
VH2ABufDF1HhsPsQ4gTf7PMNEBsJEIQH5+HHbx8jMYdwQwu9Br/zC/HUYaACXdWU
Ti3GD2DtJPxYrzt4K87rEL6zmDhwlWywIVpUwPecdWlGQsAw8scoWE77HDMzH90j
nrrm8d2qKhrJKkTRRn8zvzKdpc/1xOT9DZYEUmrZbyyzxd3goUYXEiHg8WLZZ2Ts
TQhP1/SDgqWmiX+Qbx41JigXfzBOjf76JhgfkiVxJVB0CaZQla/c21WGkaSOm1Oq
MVTxlTulf957dSf5Gi1qob1HCD8AJ+IdPriyDpIpFX4USLyfxXE6O1W+rEkJUq7n
FqD1RITek0YNGHnGOcDnTJDFuDJh4gF3VGTMFsQA8ZqQ4iAphGXChA5X87gSaMfN
sNCjKQ76XbosWsSEv1jV294Bhk5OS1oZQDKnCq+tMcgGvT1PvTXEWxW7KkrjAWPw
ZAX29kJZQHiZqGElJ+s3F65vGh5IA3Pc1MjdVau7vg+C2VmSORcphOUmg4fBW0Sq
TP4Po04nrPEthZ4wdDs8u6XBs7eANzefd5dyYVmn+fq9YXapaKAUdr0Xj1aRYJUG
H/XjBFWc82fCyyw/TSFp+3VWVP76995ySlh/Olf3CemGlWjFpR4ziBrqDrJjegL+
HkK3k5exwebHBgsGJvAlcalXEU+kx8HnnT0tG+BJ06rkMmkwVA6xDQouqJUcd6yf
MWWvV72Gxh8aTn9I6/rZ1GXUpoHOJ1+oPQsVfgKo1EOaxOhF/R4VFzFRNtg0XOoy
3GOjO90KzgIHrBN2wtvFefCOA32EhBdmnPIpKV+2Xa1SP0Oux1rjRuW1crSfb+C+
qq430d9TZ9ELr2Qi9j+oSS5QjZfzlg1T14uVKyjp051LIAzLZLgEXkODqTUEp3so
/+B5TYuVyC1aZSURpTKmUSHKZLet6ditTwVYcqiXT1Khv7bi0UDCYxNh8Edh/3nd
kiXYlbwHvxHjQYJn+SCTv8BT3se9XRYUlM6wXO6T4ngEb9P4DXuiTKP5yS64pp0S
8BSI4CBBsybo1q46Z7cNFfFoWU+4bvJ93DC+H38VwjdMFnnG6k55PSc1uXoLfQFv
zIngAw4PM7wF24ciekiaVXIz0ZUr9CSnL1ecPXJUYdhK9pxQS0D0xymBiNojSPBB
6VGVa5+fA5cnivC+Z+8/dotCNF7zATEJFJm4TZ2PdN91a8Kb6MtqOK9Kqt41HsfT
R8omfDZHle8SOLA4zFbBHXKgVgfu17VqFrsX6RwEgeHv9ZaMY2XW8+YnRjr0FKN6
w93WLx4KSsiQ1psA13N0eFeqRk8VyMaczVkrXgEfs6N0I4F90weamJ/aKYQJcEW5
Hfvyf9VGxM5QusrYGV6x0aaCxegNTxdKfUbw6q7sdtt/GPbmPKKtGhHVNaB0apwT
7pmy2j5VnEDGRO2r91tgaJ22FtpX20DVYSY86S29SyDMic9H9ABa2VTLjy1tG8c4
RkgaTAhF5CKV+cTtc8EspMJ0Tf3o2v9hldBlHXy/CjC+mAHhU7n5VL/xIs97sioh
pGIjNVQF8Bm4qGQuOpaf0kxkzxgk6YfLwhW3JDRsI9kefrWbEdBtm4wIKRX8o5YL
K7MsWLz/HmU6bWz8WZO2/PPye1Rxfa+g4jDKWd7PmTWGNTiNimW1JGKE/tGEATqg
mq+DDCSe2cbf/Fv3WP3xmnpP4podSXPHSuuUTAcz2POhp3rAEeN699KfzErP1Caw
E2KVMGZYCArST4ZIfnGPQaVKdnoKeX5Vpp/fKDg9jz9l2jMYakrI+CbEi7c3jfSh
VHIHg7/invyK+fvSBwwp0x1nasAg+w0TRnXIIE0boC51xWIhsqHpexwIeWerzCIv
pPb2OqzxgbmpcNMG5oO2l8AgtDl48+n9UIbbnis6m1Kr1me43QWC5WBvEP2j2qDC
1+rnywx4/ijwrpqrrGK5/1XFqd9GJj0RUkQ5QjEXKr/VbOiG3ANLTkMdU3FK5NDX
8fdAzSZx0Wx8fyMOjREuohbkDBZP9WB78Mprb61IdmFLW9klYqt0PBZsbHTgiZum
wXRw0fxlPBKHCGu0Htn5t6PlXPQjd15aM5j6BRwyXF5DwWgM9DJJg/Y+4P/vhuj0
Lmc26kXcUbpWtiwyQkzYCy+fSm+OPzg+E/5kbjAOjmhRUAxsDwMWSQLrojaFJkzk
vaiVqNZUnFs3pcSYWjqUWEKTQa1dF1U0GorZ3ClaVVokHmB+SP609fgS/mFO7Ae7
MLFsl/7yXjBB2AdmDnqoJOrFm4OiQCobENZyVjb5FThROtKC0g0lvuhzNo+ouG6j
03VmCDqCsjQHSRZQ2VQmL0XXlZ70DDLHIQEpX+qL7m/VqN21VUxQxamDWNYMzCDZ
ucXsEYpXlJCmucq5dwAv2mr5fl6H5lIMpnbGEEkR3R42gg6MEpXCdavBfPacWEqL
BIwUs6H+tF1qoRGlVSgGKtcAauCGk/6gm2yJQZ1WEOIy9OPoi1FfDFcIfZrBgLka
wqVz6daokVDTlmmB2FvOKrfW1e/yjG9iGpefRC0J2x1WcmNN+/TxVHaSuL1bNhBh
uSg7jTYexpZl+zyRo2toYGnU7DBvzhR9DQL9Nt5TrfTYbm8QMr3w85wew49Ubm8c
MBmrnxCGpzYy9y2cKcxbOsKLguuO6Tt+A3aY8angUJ5iFdICR3T6UQ2SVv80/u3O
rk705JmZkm7eVFRgXdV4lNHuXlpPlQhKf2Jzys603vpCrPmTDBQuuW5GUezOiF3G
1y2N+yFxknsGe1OZpa1g0Y0sgo7lj5VIInIYQAweJpoGK5HJCw3es1/AemZ6TD9S
E87JkThpRszx1iMP9JY4KAaeeAi8a931O3uwlkf12E2UG8IWfJF/QjXnBSky2hV4
9e6uhRSrZ2oSmx+NwDjsElmEfBICyVbaulN9ee1DLDRcK6tBU1GX2KLIMLk5DL5N
/qCL3pq+ksYSMM4HWGyPTIumJ9Xk2KNnQUrbGCKBh+T95ebc4Php6oOBC57/Lc7V
86W8xQLOYOPmDd9Ri8B3H4NYixKjtRb0y+6kQk7exqoG8lNsErlc/6YpX4SaGS5R
y8QLOLm65E2v/rjq/gmMVFkRLWkFNjCi4JGGNTV1PAMSdYrJwno9tT5DGC8cCnf2
/vvK9/JQQzwyIq74sI5KWwl3vLfUFa6NmLie+sT1dmi3N7eCgGPlelcuPTQ+V47K
+rtFmzlsO3d9P+ksr5TfM6lcxH471Zfs+L6AuvaId3psK6GvAEWKo6RzQg9IDNmJ
M7m7QkVKKsR+KHKyZJ+SVQ9C14e8Gz5xrLVcY/37ZEQ5MMiFUZDj1zLBRDpXSdjY
pDKxMa0q6hsyxxIOXlRGdWXW4E5ZjG41Gxn1qUook3aTj8g+IaZ5rtSe/4Sdjrb8
x6QcTQRzmDPmefPvo0SjCqvn4FX0Ne2cOK3hwrUfX2hZdDm5r82bCJil70wLVjoJ
EnXbgFMXvyZpgMurNQJJE2wv8RG6eug4i47sr5qxHa5VX75vbazPE0ZojsmJKvdK
revC741r1KR8AEukcTiga+gr/sk7YCC4i3HQnIzMJe5M2cK1e7buN5AuBmrWJtR8
rqDDNiHZO2bHagyDIrxAinf5mKwtw4Z8ssUZ+N+k87GTsCsFn6OhkDbpfcIKHcp4
l22TmaZxA37vyuO2eC99WgZrCRM+dLq8bgNnN/rxu4D2ZgDZbxz4LHDMtL480DqK
iHIPaH9OWgdA2O9bw/QOpIvJdhB9kzmofrFprVi/ZzRlZWU7xhFKNAbo5AXaxcVs
L7CCtXxbXXehsaWvR6LpCdfWtGTiNQv0gTd4+7Rr9cEiaMa0/O3UyPMs9q1t3X2M
cPWElr1SjRptKPQI9pFM0S6iLtpEV/292HxHd1XE4wt1b+0sWOK8hopKNkNSaPvK
dViBXzGhfgqmC9p/4zCwwTQCp8tBYFcY0aSR+gjADG14pTW1m5gVnQgp0YvPQ5o9
Mb2uLQYyWCdLKAudgpnRMpdjM916sPzpG9XMgUZ+9HSorhRChXqpPPqO7/SPc1pI
S/7ad+FwKrUvt0mSkFb8QeEWRZQ7taAHJ3HfWotI39TgoYW6RCwC+h4+arECeU7m
YvA1LaZ64DLXS+lPnVU+QDcPeJe/Zt31ViFjEobOE45Wojddtt798aHEOBxyYt41
PUu0QCZt6jQRfmH9H4YGRr2Q/4qArlicaoWUP03078iinDOI5qVH+1oIk7xJigIr
iT6oS90Fo5S/Nif5YPszGSaQJiQPQyGbQHPwACxT1610Ty0W9h8S/gVlB5q31AqU
IQpdHzSSZroMfHMcj5KmqlHIhU7lJrGs54cjk1IFtFGZMITPk+mAlydTs7llFUBs
mh7TUPk8CqnwIhmafaB1eDCrZRq5Rgv/7vQOFWKuuTt4rrKHPTYnbG3VNjGFAyyZ
QqcLaD2dCAUR4oxeIrcd/XphwGHV6dVK69MSSADW8BuG86C342ovFV/2TO2lnUwy
jC+3LXI/zh7VLMlxxsBeO1M2Gnoo1hy2gjFRDWU8po2ZOkABbi5CTf41gLXXa5N0
hEo4mavfiYE6aTkLiVWc2mejphO1ZegiP8CXxAmDzuPVul9jWfxzbv5hNIAfLWc5
yKu2bOks6fi7Mqj0TFCaoRev9fK73h00WZ7KJ1fItiWPl6+6qvxhRMdQTBoHRIv4
mSqWtCgNs0IGJa+YOvp9hPW8xO1VBPjangFSpjMEbGwLT06BkWY5xsrXYpEKJunX
vKbaMqSeta4oULVxWy3wjFXXJWJ/yfm8l62gniTvYybJ3M0e49ZkW3N2OSKdj/iX
seytX3n1PAhYPg1C51p2+cc35y60lDeujcVxNwVZTdeM3TS8F+Pq9QNEHFEP4ndK
yV5cDsYEHpscxRYuxjCNxAmkxj3Xdh2qY6wiOg48YBOP9thAumvHZQgv9CGk8Ii2
Q8WDCvrMGkGqjq3qET9ninByVU6ykblVP7kPAHt3iT2Id484urtW8MmH4zC/dsS2
t3bH2bdFwEjW0uluJ9XzVsQdhKqmW7yKKMD6rrTJd8p+VP+KulrHk+teuI1gUTKB
cnFCgOJRgEiYJXPbF8Jp+m4WfzlxCeDINZ5vY8LxMhW42TWXHlgPg7W1N9eoFJBC
Xf79asbG/uElb/ntK6nm7CPC4eB/3i0DfcA6du9ToHgtbfrvlrroZgs1AFVXe3oz
uogY+M9f3S6/2HV8FafUMIxohe8Zqxl+2RklOVoP6SF9xifF3pXc1CKZRV3fg8dp
WbtGySQcu1dZhiwtxkqpGWWbcsXPmugBQ00vjsB7NAgG6yk5Q2wYBfnmlptkf7ZC
aDZHi/TNAfXsNPsW6BfGB17hptMgi3whNdIljgaOLxsQgaTZWhXX3qgydVwpvnMs
QJS+Hmmtc0amZChViSRKwuodINnKTWs/aXaou9WizjsqchdZC/9NGarl1p7NnD5/
QvlEFdaZ0qmL989U2k1HWBCyQSNd1D54liRNHmHiLhcLDbOBoBQI87yFKMpMnzS6
Mt9xplgr3+SE81lh/WwOHnh1oYeP1N+gY3z80F9rGRjUpS7qNBY7MgqA9J788WcO
2rbwlIrKfHZsEhTsQ4xzafdd+s3jyNQmE2oKGvbuwqEZNrsJ5u9xlcxXxo+Iakc0
0tPuwF/66rNyGBqcm9vcAYvxWzdid4zF3olozm/t24GRkhLPoOUnWAHSkWnN+sEl
ynJKYRwSEofnZTB0oD/cuAUsTyKIyS9IYgMIyrQoA5OWzPrfhhzHRaFH9KMM1/7Q
4ARfTogihDo6R4ovDmejqk7r7aN7JnTNXKVdgPpRfUykiNjc/iz+/ZjaierM7/JQ
TmNnmXciZfj+V3bjHBU5Zi6D2yQl3Wi7aXIy9uYoQT9NloldNvV+yBEDkF/abnYY
eFtLFIEWYXUrQaLA/KGyRHCAx2bDa7FcG8DmjHGmoTVhYkhhDh1bX9MqinLDA1oQ
btdSXAJeuFOn5DKkrvawhLB5HdMxbpiTNAwFwdXCJyiSK2K/A/A5CFREPge+Dh9j
QWMj1ISLkoROSteAIEUH+CHVvbtzIDlb1Dqe0M40Nh4Gpu7IUmxlHSSZ48ThWcjC
+zGidp2W56Y16cOrJB0XaOx0RZMGLM5M26zUbK3tcdHr4xuztToTjHB4ThaP72OL
kDCnD5h1q8wcM5lvC+eAdMlvf3RTayRLHxcAKtTicociuIsqdkon6U6jN9lpeiM7
zDmFUo2hu7nA04h6w/273VTAtLPuxURNsIBvFhadR35GFAtEwgqZEX3FZfXOGxVv
MhoN+s2lS6SXEuBKb/6Gq5F4wjZvpLx3llxTkccZ9hDLzjxi6Ck1VaoM/xNah7ra
K2XhiIglgewzHQPrJzw0QBKSwdkD3WWhBFRhsJC5itOWBOloYQ1TPa/qslqws8Bo
7ZH/qB7ElXPCpyPO+2wfO2k26UtF/0n7suNPnOxYangS8z3FmFHTtjggWt0YfEUE
oWuk8tpALfqYcTzcFR0mirgxzDStq1Ds3YD/ZeGcMAQyFRzB3OIo6fvAylc7TbwQ
bK/6CnNRMGjrHlApAmHv4i6Tu+Fn2Z8kK97qaZWd+eY0CIxO0uB9G8T/AbUVuWGQ
9H8/YlyzfN4W/z71NaMqnlXzldfRBSJdDlBtzFsKJi2nZws/zBtE7yXHMD7Q1DIS
Xa29P1jnU26cfy4EszN2UoYekZCPkLadk3sB0YHaOhTU7oGhM5QrwTiVBxCNCMpf
gdyicMro2Ju0E/+7FUmCj69ea//Twm1e9iCqJTddBDDU9xMODuT/3fXR2jpYTBVZ
zbTh/zwIeEqVq6PdP5/wCdH6RjjV+F4sCBEnoU27H61IEzWWp3EGjXsmGEcreBws
svPXbhomOsxjLHDMGREVdizFrEyWs/ofpFS8YcxKGfiXv687RgQpG5fHi6sDYKiq
8st2GKUWLpF3ONaeGUS+XZMQIi24dYhjq1bmv4+YVE+DzQCXFuXCpD8r+L6bxqsW
UDwFpV+MSmil6eONXmh7aNaOUNwHDlxJkRYieiHd6XAmH8fMrmVWOnbcD5C39f08
SWr8sVSS16Z8cVANmySBwfp59jW3aVVGf1zdbmjRdsVH2EuYDcp5comBG0DKAGoU
CfI/M7XVkXZhWwjXCjhP9RCtTPkkFwkcb1lNuPwuE0Ic3Z82Y/im3w0E8rDA2jA5
qg6QSZQLJsOjjT5BApSCE7qD/l4VuB3T+EirxEmBdz1bDYL5y97ZhLXW2e5W10go
7GHWS4jE08KrE+NsWT0iEWApPHwAY0cnH+MRr3anDVHrkw7TgEKoBCQe46DpqeIc
78j89BO8UxuKVuqHsCY3oS5JeiDmICgpJqUnDopH3GuzfhqHq413lMooxdwt34wE
PBC8LGEqxcAf3HN3HanSGydCsPctHszhBzQEDG2m5/q4pwL3D4Jsv2+YUlJN48Dt
kP4i+6L9ZU5MIo6QyZfO7pTnaDRT13KCHIEKArjVWXfSbS5YGr2c75VPRqAP0gE+
BcM1sJxEQq/74onHX6B+wvF4fnnQSEju0YznZ35FzPSUDzDwMXTyEY3oBTEdM21E
GxRgsw7L531nM23+ISXpmkEP40xKZfr50sh7hnPkd7Dh4xJOooYhjyGCxUKtx/3w
r/9z4FeTRhjYdKbGvWH4ZPC5elwo9OQQBqENQFLrNbQfyamjygU+uVJMvGQYtMqZ
ZQ2EOn1CtTnWwv/BiHktfaQpRkV81Aplx3kFzuyI8vhUbqYhyJ0tcMFM6Ih3qA2V
7PUAoVUMtB/LZA+zGFcbGl/v2FPaTkglWEjRwjycglaBrA6+a55AftO7Mkn00BL7
QLkbDJoNZboe8BhX7qXnjp3VIc0JfIli1BFHRm3Qewpui7bYJhuotwpkfuzs1XE6
LIqy11n6oQKUoz9+LMVyE4FSdSNdTZgSyHv11YjwEgUPPbIDWYTXdagRapjl6g0V
Fbh6ObPB+OCUNmtjsmbFjI7V3jw2G35gQKnwzGZZOImVKRxeQsFLhpph0Hh41W/O
e58FURVVSswVZ1kV8vidMUA7b7KWZ6DTKwSxiN2V7VIdzGYI9uDZjpMmMUGWP+/E
abE9k4Zss7g4dPojBlt1jIyZ1MbB4yuGtMlkfK0EbtBO2MfQjHgCi8So65q8yeb4
4Fz2Pown6A8aJFV54nUKomWsyR0uZ4fNFXC6lhUGslqCcXrdIXblS5Oea12dSPs0
KRnoyXyh5XhtLvjStrX9urEX7rTMsYXZuVFO2DnkX5wreDWJUd77zH+WcYmBCM4N
74kFy4AISq/a8dQzCVJ7u2Be25T5i0QIYaNaU1H1SS2n9zDnUFHFtqyWagfyu0P2
rBVwvlskLq6oLzR8xVy4rP32Vk0ZTylLqar/xgBGRdthMy4miBkPTQQ4fhX/sOL1
lo8PNgM5SverQm0j1JnKzLGWV72L9PNlvlLmgt9weTD018VoSSBsIwBPRh4m03m7
7LMjzVzVajy2uZt676T//OFpTFmrZfWg7zC3M2Cu2CJCe6waZySQUh7rQtYkYl5E
OLF9+waJZUkPbiVct5jrWxOCo/4TpAZ/M9xV9/kXW6R7JPn2ttd3fGUIOYavFpCj
J/1fblvuxZOV4TAOLr5aFdmZUJvhhWjw7GxWjTDaYF8DHnoQ5yJSyzMx3paddVQ3
lNsYYvIIV7v0fLeLxQaGJlmeVfrBXPKZPk+Y0FgvgVh5C3D3k1Y10axRXKcGBULF
WPSFoWoJvf8qN10hqjjqfkrCrcefrYmpcnzxjjFWCm7uYKQmHVmGbAc56jz/nltb
splApRZtly9B7Sma7ctBLsPkq/n5KKhiLIviwKvJuV4ZxYk5dCFVs08945Pubk3v
lrLEtwXhlfb1DGR0LXvAwrrvbolPmdtR9rzxsfAhVvnxBVSXHyrO9bcj+M6ihdCN
BdIgTZiA990Gt0SuCuwnfqtkN8CVK99mv4bZIYzfh8Tn+OwlDzDBLqnov9J1Ycx7
FJuXG0IIkJ6dcaWME3r5/zN8SD7GUuT5s/0jq+b4EqesvTC2IW+htYT7fwKwq7cx
hJjERLZ7mS1wDOCNbJlCGfrUVh/Sjbt/pAEYJjeYwHNtqAt1l//HiR/pjJqWa0Uq
NKazzJns3gLcuvXK4NwY6VJKj9DLZeFqa57T5O64vEIHNhtFvTkqd4rWBDIya0Oy
/bV2JehE1szS3RClpTm4Qkb6QdJTFTl3lAycCxur5M75lxfSR2KGynKDZKkW63oO
YAr7IccT/RHCTcgfAsvrucFxcmfqZvt3pwlCDxj7Z1Cv6bOba6qbCliOavLi9F+B
uh3iEIfsH0ayKpsen7cMeMKhjbAzgFzCdYJClefg6cvhRw6go/IyIkGvcxNzTKDi
55HycOQqHgl/159cqcJmDtK4goN0FZrP5+7j96QNqwWr1lAbVOvfKqKZyIYlUbx5
h6WADACiTnjtzNxZPVFmsfPLq6P3E/sIg93mENNPQzYGJLSw8W24wnPjuE2LwvSK
ScEYKLxcGYtKFy2mqEZE22J1WpUGK+WEAhbwjGLgMm9nq5KWFRGvFyjOvlwKb2bJ
F0mM5D8hikfUcF48bLd3ILZCpPHNHKkCdR97jRg/iXKGwFYuLslXNWe3ePVx0XhI
x/K+tMWDXil0oQqZhrCrn7IR833O7jbD3Y6Iz0PyKb7CPKbq6vN4Ar7xfgdDXyuy
lsknw00oneVMy0XagJZOuNxj1AaiKNUyggYPbIRj+1oJPIJ3dTAOoH/txmGXmFmn
D5eVJtsoj1MwwFkjpq2rdnAs3J7xudmBZzGu+hk5CokIJouf8RGIyxWv6uLgdUha
EA/enC5kro0ozKDB7tFV3BCvUZhJMObmYb9hdfQFT+A1VqRCD1rxxw5zEiN9a4aY
0ytOYlkDlHlMJMkZaZ6D2NGZpXuOYmULW4goUoXb1WXdquyFgQ2dR5F9Z4Ep+6Ed
vQcvRaSSFDiajBg84KeyxqgfIsyS8uGKrX9Zgh2LpXpkhnDDUuqI+NYyEzhsGN2Z
SbKIA35143fHPenshmjQrHf3QmJ1DRCo9SthY9xXnsLTY09lBxNAAMn9HhopyQBD
k0hqTY3zbeYDI3RyVDefF2fXEjPQ6vwhu1jRK3UmurZ8mfRXj8V9Q/xwvPjcVOMY
2SBlRAx3L3LLLS8YZZ6VlV7I9zMEfv/4y/UMqXAvOdkirn5zVPTGc5j4trzDuq6C
hSqHbOpefh1vJwerve8cMPqrzfgQb1XEmUmDvsr4I5DCMrkaOou2WGKMvwrHb1qR
VSl2ZKJ3bpNo9jarQwRKeT9kECsUmdK45vGPE6oIPmEim4UID3o8qIPaYDWi1ANk
orxBRmtV3liYxnU118ukw8o4KZiv+xR+PTwE6+In+5ylhmiBAGOVDJOAj8o75RJL
xE/SGzDrjhp3PjFWds1+FGUdGyusLq82W5Pq+J/pnYCyFbdHhI2WU0OKcEsOXTpI
mDMhHYCkWX9qjf+lHNbYAt10Z3xkfS+Nvrta9fc7urlfwzzdLETGOYTOZ4gd/0aS
LUzl9VZ8BXfGsvJHLSNjC0SeswbDtbQjdhM3yLryNtt3IKrx45NFIYQDFaKrx0zD
BeLV5UVWn7VVQlRqL0p/HnxuHX52cZ6Pl46d2d7eTglRWjzYATj7cRrs/H+xvcrz
89vBSDDWp/7ZlyPr5glfUqKezjA2e57f/hxib8dP3hlY0PMXbLTAEXjnN+pjhyhm
5+Z9wCsIqgjiy87JMxmarl7BM4BCOaajzKaM+rTxpGT10LZkiyRJNSWREsR7IKss
IvKmF/rfpmTR3m/Fty2scqaZROuZMefVH3hxpejF2sTG4R22rnO9eOnMxeJhRDDG
TLFsGW9cuwmMIlAXEoHM2SsDus5qJkBJZ1RTKhkzDiXCBU/frTSt5qEyHjAyNVUj
MwPc+hEvZfrHKArmfi8T3ZsajSYdUtJDSHhPi6VpU9m3bFEh+aOhB/RTFNF+HFXJ
tFgFK67MxWiSMkqDplUCN85P2WYaTs2FxG+vs7MkiYBHbIhnGI4giqxMeXrXGVBC
ds0S1/No4OG4g+rihn/3V+ZQQrpKyQ7tT9oHZ0PyxsrUokjRCLoiwoljSdTG6BuY
UXVUZUAh2QPDWqfT13xpByXCuYQ3+AK6CSDzmsJ9comfNhy4A6UagyYeIkG/LBWg
tjxg9qjb2/J1Ta+IRSM/TVdkv3BFPWNS6yGNjtYnkNkkWQa6zbOGmOMul1p68QuE
mkT9HvDJPCZrwRmvksICHCVTPMnm9sc5eKSDHo51nVSiOjfIOHa1soIp36UlbFPq
x4K7S5xnttKMNsZZwEJw2Ax5aaTfBdRLRVcMeTOD0Qt0ygcjBfPvRM3MulYTLhv4
IngbxmP3V24n1jqXcPzYhrkRVMFulCXxpuBfGiCx70qL+5Rv5lHnvu6tJKIeS8kb
Ti95eBcbW84kJZn2qQVK3M/qKpaPQx8ZFwtoW3rv69Par27nr+ToGux274QYGqYI
MJD/N6hurFo0X0QdRR0ZD/mE9KzqS3AUqwaa1zEhJaJs7ItIRZ9T8wV5vqNftMea
Am7pvzcvPdAv3ByxS9/exwLrRmB2UVI1yqhKoDsw0ILse5WTq+5Zp26OGgE0vPRd
XTGzwwUCIdBrSGk+fdCyM94y/BhmVfRQ3J31SNWlPSCJrW87yg2pEJFJunOuAu4+
wrDGGWXUsMddlbvaUBtQM/4EYFQFl/aonlHSTT4unIj15rFFBpiXm1P9RszjOmSZ
pyyCElMKBWiGLCQLPEQJBXkiBtbNkN3XzbCYBYXMgiN/nb65dfajbXkFFxZbSTQS
CHmZbQUIgmc17wZazjWC4H9o7H7u3FGtUGYZ722wkwjevJGHeEQBumu2mMMgTCsI
3gyUxcHR+y0jHsiO2Mg6uPt8ogypvwx60i/72zy/yjk2WNovM3Lapi/16migvFTt
wnUFu0he0GfP398i9wpFgrlOCCx4dNau8FrU3xINNfqgzKiJz1rkhD30XuDvPLy1
P6zWmAOdEdHy3YR/YnuLeMfySBZy9tnpvOlgJpBGYZO6KW7Xfa4hCjZOYHLGKR3i
YEOmeLP1+o5i5fhryvDgp828mnwwpoYfjmDvcjbA0z0kY2xfFtGSluHwm+j5ncM6
pZo15wJRUriNsNjjxyjFWw4kzZgPX/x5VYo0yUH6IHDs9PcsrR7X6FJOpcdUkm4o
T7eI54qlcq3J9X8pM2umZVWUXOOSQAxfZ3uHVAfFu2WjJm7/VRaUml5EhGlIXvT1
FjVKZ0oMPj3Tdz5kpIvbCfeC9tQPMGl/VZogI6LqJo+7VF37d/wIEYmIaPv9J+Sb
OdBtUOcVNcetW+JbCG4/Zu28LgjL9nxuCnU9TlY8kzehrToxcqWe/nYichg+8ssc
KPE+rpDcdLcWF+a1qbRfBTiQrvg9iU7pRSzrWweRXrgeSVBTvUg1g6w4nWhrzPv7
PD1lwEtt01oD5CVOvWUMoog8StWjki2UM6e0iK6O91Btcl6fVx6S6rAvwe1OUdj9
IJGeJmAU4AdzI/zcTrxn0EvBMxI+vtk8cr7UIcK7NmV6zSqYKOtrFummmQxE93UR
lDSvfOkZ47GGJxgJSbQw+Y2ORSgMxPRWxOXh26yclFdsUDojuAHv0083tvro/1tD
r1/0FKcS1BNqMTy4bZsZHYjZTGYpzw+KbjlSCEg08WiYT+BPRketqscoppiFSXhC
vp8E33LT2PMNFD3iy/qgCPiKdy++0EZKy7HLiPQtumHk4he8UE6vSSvkp+ZhnkKv
X4/lCfHUB9HNyFAw+qMaOm6ig6Ym7IcBI/KBRdN5wtcTEBXIV9G1XpKCjKExT00H
jkJ9dlg9aulexVnWLIBMSTfJg1Db1Bpm/lqPUWtrcrKRsDTbvUkMpUGgsA+zayBc
rncseWCfuPAD0XZoZr1XzKLzY9+FJ8pljyHo+OG/QRUYGsxGdUUR/aNeJLjNy8dy
8sN1qNIhHoFJ8cYl2OVdzvD2Lwpga+NHBIdqWp3GAaagEvKSR3XCCgveWFVV6R3U
rHEOsAQ2TCz8GaWwQyCzDe9DE44/IGsVVn+fQD0cs2z+QRPAbNjBnD8CRIrFXg4U
X7WmVL5ok0Ba+/L+tRpXorOPsUg+Qmu9s/FoFFAnLfYOXT0G3gNr+z7wCPoRG5T6
JLKeeWY+EfPdt5Delz11VD1gj8UQjiqwQ1VjHCctLDqISKG3qTtq+0ZYIBhT+wC+
+fTAdztb4kPLIaoBRa7926luSHF3uTfU/wm0bTyz8BA/Mc1GexGWW3Wt6nbydk9b
5DUS7SLyjpJDrczkNLvZjoErqntRgN1l6DFXmQRqz+S4BmU+HksUBo44fd6KqWdN
WUuM1apZeVq0q4up6POhaVlD8MFJEvvRWi/ILVx/BkRfUEhjidGCXLY2pLi3Ijxy
XtKV/k09Ks3Q0QVHl+avYjEFOjIOUnTR5gul6WsaAGqVFIYOLwJx4NAhmm8ry1Nr
TlQsz1JlrNWfKC6IG/qnk5ZYrH7LM47a5xqK11AF3caxu5kH5iZ4HEbktH3dORvu
mhsHWG7rTzZh3R9KSbC0L5g/whR9dxl5V1Ke+mS8NLMm5oE2/vOckMK6MowZmJ3C
kVQB9vxpE92h8C/FyuV4Ops6UJbz6010HWD2aE3ALzU4lWtx+WMfTeoofEvLDOjG
z3MW9KElI1jw6tUAbGPE7sxaSNQkEilGCmRk2yK+C/8rJg8xhWe4KUSt2e3lPWDJ
coke40+/dQwL6PmXJ5EmfnINNM9l8Rcp6YxOvjXGflx6kAYjoGoQ3ldpAiBgyHGw
lvJeARKRvPmyaHOG+mqMdKkyT5IrmgFbJCKFGBDC59lPFc7cMbDNEgQSyWsdWPk9
yIPrYrFbKrdhpOSR5mL3GG+DtBimfWBHtKvVWHVwhEbeujK7rDCaj5KNfVOO3EPi
hpne5+88cgzS3Wq5XVISck7TAmYDQcqeo0IZnXfKrEVyQy+jO9WDQeD1VVqNxzLx
Ddx0e0swtM2PQQuWONgVnv1BXh2kOlWf4JVUv/311T8H1GJ4oE4PJnbuNony71MU
2MmmWRqkeAw0gHM74KoolF9zV9LkwD3jZ+88ik0j91CV1POg9m402KXI44do2DnH
q9RY3YKj6ZU7dle7bqyGt0b5osZh0FAqyJ/Y5pVQ/ucFI/ZToRUg5G16en/+SgUW
5u8fLx+WA9E6t5qMbUx4NN5RFh8BDSMBGv0K1Q2zlznZA3YOn/wMFKWo31bA/s+Q
BvGx1NAaEBri2WYmFTmzv4xFNuCcdQxjwcuISERs/B+UTxIUA48XnPBvdEatgPdI
McDHJRxRAA5IubQkjTHTcw4BbSTNq7yMIJ1aNT9Fw1O3G62ly2RsMFQRFDWYwpSC
J/6Igq8C9FmUeTY1kDu11Xmm5bTTlHo/ZooYK8OeLQt04+PVBTkfT+9xQ4nflwrr
XEjbZA+NuTaoAUVP7FzaEcxnrIVBByW/Xc9sTnv9hcfVQ0Oil1eaAenhFxhSgvIx
USMD4ifoGVDj86WAoz4jlRFoP2+SNmUZ7R1Com88rxpKs3bc2cxWHUl2NPKAzavO
V3ZufF6mBeM5SAOaeuyx3B44MN7PixoBi1LMC5VQ3crmGH7qF0bqZElZ3oGxDswV
Wjl6NMf2ODY+1NQsZM553ZNphDqVKwMHq/7DUd1H9rQj8zeV0XsqVhTYNCigp171
9mIEIxfD9MCdm0lvgBnXAa7EbNa/4xohg0FP3Q+Okcx+UjWTnZzymeH2Si3gWBJ8
L1xNhtxFPfs43WOKeT+scspGi0RPC2+2VANKOuwYlSE2Ic8ankJ0B4I2lX8HiSLI
9YCr7wngIi6IpFCP2WYJ8LuE0eG1qqwlndB1JBMdimBmO7OoBFWv6wqmqQuuWOCc
3QSI+GmMYTwdtSTKoxMRRFqNm2/PAKymUECtNafBBDjA/i1dGAuJ3o3sWI4YaTp/
4t70bzEiKUk52OGprl9IHItwHrtR9k7UWxTBVtp0xenhT9NveaQqkpgcwFF0KI4N
OkazxdngBUDuXoZcX+o9Nfl59I/U4KD7GAdTPlcWn0RvCnlUMHHxLEjrp1DMZINF
srVd8oYjCuznRkFfl3uEDpmtp+UEu8kKO7PH6qN89DzFFc56v1fBHHl9sdzmh0cH
FHMUP7GGl1ZF1NholUtP+uykFA1ddWkiM47t1KTVHEun5HEsLupOGJcu6kPlwee3
CX8ZpeaOH267h/uAZs8rIyvR0nFRAutp2iMF2sUm++ojT8ak3gPhfZgKYeRBHmQ0
DXe3AX3FjqGNSdMQ1OdSIVYhJgINUS2VIsAsNP0AYmH+GBu98hHHC5sXri8hfulx
kVpxa/7bLn5gOmVovn0lm2WesowNC2KdSiATZi9rUl3pwchr3HetS/0F3gmqNdnT
jx13eqnbKWj5UCc8h6SyVusAttbC7Ir3TSdpqPYCR63Takl1hTuOqGpUVLb+Jlks
FTRcn3goxZj0UxEHkME/R8r+iP4/IdZlkv6keRorLKnRvGjliOYVd5EcuFqLg7zq
BsWexDqOn0KIxVWhYe69ys1eUOcX27KBiuFO08I3EsxkLfVQAD3MFwBFfs/MKpw2
IwEqgDgFq/d2TrYZtPVOWVCd5NpGqqCZddPwOB0nVlEZNH9MUJ3pHwsumnqlqVOz
vMHqeKKT7oXOnuLLi8I7EncFZynRGYvxXHmNE9jLDaK0zuajHCViw1/hlOVWujZi
x9RHL32Ir8W9x4UTpimi93xHQ1IRXaBp6eejixGidja5j3AGYJ2nr0r4BQdwBgPh
OO/H0NjibMEjPKXhOyu9945ljqDIs1upnhy7a+GL+1gwBKZBAwiWcdXi87r1Codf
OQ2cv7GenZPMn0hiwefSPWhyOzinqJJQB8eg+LrrorLPGq2ZDUXKOQYDcSlLu1jl
Av7jYvjMHjcOW1BbOUt8+G84HAl7BwmkAm+3wbSVDnK0lozNLZvlxbX+IMnUHB/W
ZjMzs5zMKHUO5kRdlJInoFu+SgbehznscchzTJc7LINArWnJaqKyL/Bdq/r8IaAy
EatxdKakeQSKHMV8NVAjHd9nL+O3QubOr0x7Hr64bqq9jQexsifXP9cTe4yVJI+D
+nq+4Z13Rrf8S5IHHuFAM87/FKdDXEQBnc/ncSsp33z5igrjK+MrfSVVWOHS+nyt
hF6TWbmOt6OmLNPSOcY+Ijw+zG+sOsGxbRqPjJm/TUqYXL4xJvJcQMejU7atTmE6
ntvFv/yvOUIZFSwn6ZGSoXKZ++qeNwpDS3X+NrM4Opu/6//otMst9ElnVYV4yI0K
0Aw+jshxWE9fL/qN1UmiKphN0sdNlaIVIC72Mvn+BdRoB6fN+mrq0BCVqHeSxmz4
OdN8/pROth7EdeqwRPzjFHkPj8efrNQMuEpAu8IrqPl2FQjDU1N+Lgp4wtCWaYEV
t6sleew7l4LqtErwpqTRtmhzP75hro447WWLUUBllAYbaRExU6a8WN87MEizRc03
NuFpezj3jnEKKMX1Ep2C7KJJKZtzFHdVJ7Eqe+B1XeuD+w1ghETMpKl4QUs4ZBtI
LtyCw2SX/aJi0LyudmI2y0XJs8DhihZZaLQ+H0GVuoxNpsnwuagABEeTn9L/seBl
iAzRuX/TdwWzd1vaxSyZ8CeTDoi7PQo6PzjL+K4eZR71F9vsI2vmjaINxVf7C5DE
HryWHGcGnk88+so+CsSfD+GK7d5laDpXceD6/pRVf7TI8s2OFiSB6TEQ2XJhsFeO
qkMXiaxv8lJroZV/V2GtfwJrr0/70gouGuTDueG6l7PeLa+3kNCi5luE6TuGYK85
ce2EpNuc4vGQYCQGOZxznN10x2h7Sdmvj5LawZVpgs1/cLeGmZWbiOU4qWYfa5I1
pauwaMb2jJNbEDNSxbsd1+lFyzX1vtcEedghzsFO0tDzWWO+lw7HVSVAeKqBoTsU
nBg2FsSEdJakhYHhvBODoi7W4QJecKKZSClFA09kZtz/FuNclbKDyCN7WieG2tZL
ZCchkrqfJmv6wuWzjllam4ZXzhiuBpnD7B7t5drJbBQqdZDwXrCJClibwAXnZbPB
NUC9r5bU3HjiiCOl3PLnLp4Y2mjeMvAevv3babemr9t6DUr6V4ZC+DlGJhh3p50X
mSL8c81dz9WQmxLeakdl0TvYjNmurH78lh9gVAYlXThtRpnxl6hfUx1ShWCi6B4k
2spfwFXFwvPaobNTL5h4pzprXapKk4rUVVPNYV/4H6Yrs3uwUVBXkqZKyhFaaMCZ
kLH77a13YMV0lA7kfrXgBfAAu/kU+L3yBSv6BZciepwdJitWSQvqrQ8f/95oBoh0
xUIt2VO+ZuVj+47kjLbZD1aqAZbwBSbIKNYgPDTGbeCgP8E6VcmyCsupEeK89MgP
kJ1omwp/Vi/bNLUeJ4GI1KabJmIDQVL5+WCWVn0qhlhpGBjQq84Teco0hWLI6cHO
B/cHNshQsq18QQ+BQ9e/WaEmyUbslrrbNtXxNWov6mlSeENcykHk96DlzyOeypl3
wAuahvymDRH971NuZAdbs4ceOqKfZ81OhgfXohz21axBjloovcosGRE26qtzOEoU
drdsE8+IQNufuD9j/NIK+ry++tNWz7O5BPQCus0ZcUhqLCEqEzePKF7HyGod1jzO
WLuq3DTqVunE07hitkoQQYhEDet9GeHJY2iX3CNi2Z1qyyR7ISJaiGiHeiQb6TPm
3JpOUu9xQY98nrTknjk3g7J2nxEjdDGMGtcFD3rnLXBtACcufMsRFEx2icZnCz4q
qUsi/KPxuzmSh2H+NoZJuBit2puTi+ya/XQXooMj5yx1LgX7ES96OtjWD4DYtKug
Epw4qJMFjD8LuglVP+D0D74XEGr+J5S23MhzzI8X6TvBToys/OLUJxJR3H0BzUoE
FVxRn2JZpWaKJz9agVN5xbbZaL44pRzbMQXwbZ+uf8nOfMMaLejFuRq3B/FEzJrO
91WGnAgendCdZwPh2iWXWCBFuuPL6e1uJCVItah01v0sGlt9OaAwalhm96gEfE+L
cja3XToCKJwwlK2mIji21+9VXgAB/Sr+yn9gnS8WbbUkot1HkhaixHoXdYtomJRN
qpkvnZcsQ/BkcZgRIr46jz9mYFgqJq7I01jr3XjNmK1ZS7Qnqb0lFjHSs8mYbVUA
fOfJo5QhJywFoUWEYFMGb1IUtILlAscP2r8FjcSIXywcQGX7YN57ESVacy49rpsB
fKubYix1PuUrY3w8k8KJQIfcNe7eimQmVjy2ZvskKuHLfqEb+wMkfLCpQZRVbRKB
GqppGKzV04HCLMDX8DZBdknsmsBHC7880dB4K8a3ekYw7sWejREK79hxV9FQZtOY
AbebVD5D9D4f5BXLiRWIip+ggnrr9Hz6+Ep0zalfU85PLSMch5jPnfklWzcKyb+R
iqnCQ6CaRMJsECs14168xYyzGA1Eth3tPgqNzX7hy4BT90YTndtR1nqhn5gy17xu
oRIfxQ7CoM9BSdgx7H/2BdPy+nvtEbqCBWaObFJf5RzY+CoPp48bhAkp5TyoLn2Y
L+WRpAWebBMU7TqZHCo8ethXRCNHZZl7WM2Wab9KJkmaPCkBdIhFdyHbKNemjmVX
D0u6HXVQiMRpGGB0nmvDO8WPnhIDLFBhlJgAN92pQ+RHbp+OcYIh33FRy0L/VajI
Lcg2FugxzKH82rjoob7eULvWcj1zs7MUdcK8NRfTn9ewmSAyfXMTVCuVwta2hOVy
+ZIyHn615JNCLdELHc9vj4NMTebD1z7c0j42WVWQAUCnrltSk5ioZjZw9NujTHBi
XTURUKM81TfE86DLzQdKgo1YREumGXjJ3k5ZrZ+LrlMSnnOOP4kdjrsYtiP2SKuw
RD3r29cD/vHM9Ak5ZftDWLhP6S2d427VE/SgPI0/L7Ix+4z0VjYdtbvGWupqTYqs
zcq4L0vBXHNMm8MkVdkwMj+J9+tiUVq/syI0C7YJvVxrVvBkt/0gTKGWJLYfDwoP
wyf1r+J9Vm5Gnn7srczhn4FhLxq+5GVuKxBHR0PDyrWbPAEDSi7TxzYtMEtejvCm
ixk0kSgTdPM2eQQktrawTXB8glXnk+kI9Byb/gf0FLn37ptDkoERZjzaLjXwt32H
qonUBzPOnCYzlircVeToDXLGFv4n9RPMMmBBwAmq8DKv3uDhNCFWKRGpl0byeebX
d0dhGyBmixyud74NuyoKc2g/4C0i63oG1WkYi5hpONQ4CninoHZofze3laQ/+Zpr
NP8Zd7WIjR0vo15go29DAWFj151QK3iDH8s3zewoq0ZmQGlqDc7QVjVCk9YhL21A
2MhMVpfFwrGOJ4Dz6EHNUkj5+pbTl1m0KIyOtQ0GfjvuoCxlN2XXYhCP2c9VlmKl
1Y9TIyZHkqf0KRLtBqUWwzqQFDyaPYJvIsNEJ5rM6XAl4LVnh0u4qH/x+rNBEmoC
tOJmykChbBdjmIDPCo/rfF3m7J2RljGb6Ngqu4a2kdwGYKiln+Qkd7TJAd1cWjOr
uc8c2GTsuREwxD3ToUe8/c3iXhBRHq8FGV5+auJH6BrdmzeUhzLBPvZvBik5DAzR
hCFgcr5YoXZRYuaL/6I1eXeD24tNigZ7HbeH0XMjX+5uWHzJ4sBmCnBlLXs3MtF2
7HOVT2G05GJMEBugIg/7DZtDrrNjMfptTJbJ2BJxf4UyK4U9Nlhx9im+cW9zq/Gg
YWlNIxc9E/PdilVU0T13TTJwt7smU/h3YHKaEmxgwtKbzck6BMQZvm97pAWlM76F
7kN9WzdNl4K0qXTQMYmAw18FQb3wyXiGaC7FXHbjJDdsDYybUJKeEnmQ/HwMlvFw
MgJMcjLa4XLRfz9NU07u7qTATlqvYRcbsrp86vknIpQ7755+xyAw3fQkM2xfiPTn
VuopoGOCxFjl40SQZv83Wt9Rj6d3QsF5ie2g9g21q7GvqbCf5I6hkq9HoQvoxvyx
bBdLmQT78s2ZGQMVP3QwFXP/41lNsq/lqaeSEfwgjARAU+L3E2s9rhl3A/hZdVIv
xdPelNjjt+aNMunHWWQ1UWPe5cQvMcnMbT5Rd4BCoET1A91ot3ZVil4XWHzaEE7q
xjLYIKcwGRrDWCh4kvyvHIkD1cXAMmbxchUlyBzUhIVre6niKP0c9BM8rpbxg9HX
ICkqwl83LP2EnF3zsAMTMb/34HKpKqL710E2Dp0OciFeb4kY541jfgSRYyqjyf3y
FFcB7VBLg8bTwfVIlLW9YFs6MFcCh20Tf7jGom1ellQzAsO8xR8RZ6dNx3XHXLwX
Zvx87Br3YAkymZGoSBnfVOf9Cn8osstNtMUCCHTKWf8crnlhJ56GKz9TQ+Fb+KQx
Q72COgSwfELGJioadGS1KooVjFw2CZl10/KbTJHrAl6gkEZGezpSXmujS+kEj1Rq
XJR4hiGBFI5brTlGhBI88yq7Vf0oVvYVHicg8DdEjosUSlwI/AR59morZxrdjPgd
pxdyKMR8e9UnOkKxyVR6jkMD7njuILojg141DoNKuC8uArvn/XwGRCHNh1NPkCHM
H5nvgHMt4nj1QHBimYw6MJEWjfeSTNenkPAUEVLgacRhimTdr0fZIpP+m85Cloju
6zmO/LDiKZmcXILzcae8JBppPmJk8lB2PqLcULZWDOYHOSnfm1knLjh1PvQTePxu
Jb2pGQkDbohBStpbUcfAYiW1BpFcBv7yhFzGJ+oqYjaE3Z3HljWo3lYX8yET918+
Ab+cpqDzkLi6MX4BFhPTpDfmzAyCOglAIY9DrsnfEF5I/3gGI148C/AeDBO1SHa3
9XQHRAgdsu2suZnYNwN0nom1DZLJbTTcbtGDIP44YhILAgdwrkHohwdvkbvybz4A
+npYTvvpG0bWCmxCLEwSve6rISDPGcj+nnMSXcmKFmleJoZ+0ondUP/XAiQ9LA24
60GKYPhzGvf1SC+mcS+3W0nG3ISQpMcuZJ/4ERb21WDBT/n6RIeJeFaV1Q46GE4j
3tX1eR85mD3FZ57lRVnIfqjgfRWuCE42pEUKOba+X4eKLSrQXA+TqJbB/jjdDibU
XXrLVgvJoFcikIUJhcnETZjTtKh7FieptJWOxuPGyokFJdWp9qJmbiH+s3fHQyDi
T6IP254LtU/Oo+IK0SiW3zkVQhIBcO03+SnbqGX9MDayAFxc42gzHOdnPfCuN+vs
HG52JkjiO9CnP52+zYHkuueSYA9RpwY5B4RDdSx8U2fXDCWhqPfMbzINhGKMqGjn
b7r1SnRWifUIw93yo+wVFfVsQxp2voryck7dhg3b6eE5pjkoc1jv5ptqgtahRgWa
WhR1pWClhwRLIa/A+3CXAPhqRy56JKWi3apmza9pQvwsXGE6OaJahxfbU4lNo4Rk
LvpWgO7mWvAlsilcfHS9Eqj5Z6Zpsshi+teax8QzN5x2/CTF3tZTAGA4Jq2Vy3Ye
JXSZKbIjQifZgQIYThGJRobrUba75aOogYMsMblIVOeBXlCaCy3CPdXQuJuQHEcP
c/WI0B904u3054RibZg9iFFQ5nR1n4jrIwvl2jQgh9/KX6dCumqc9bE+5T04j8bL
W89liMbILG346KDyGo0iVTj7+HFXYTzOA81QkLX392+mQa5QVuEKIseRHf0Dm2PC
oewQsTyTBe4LI3WTVVPatp7qXmYotwj58LgvXTlDGrNP87aMr0UDDdFBoowfkj9A
qDXARD1fnG8oF398P7I7Vl6yDpXnGg4NvRjKqeIX2/qvwMc+unPqpAd/J+LED6PB
BD/oyzkTdTDqPt52IBYG0kh6sJEvhHZibtO3d173BtLmjmo+PdHAGyzcttd5ASrT
mUqQgHPBDBZ8UzV+hm823E7TGlaIVQ7GkAbFoQD4ZtEXeM2zGxvTHFg2BPI6QrcJ
7F/hSPPL/IfspYFOWVo1eI5opTuhXOasM8N40TEWloqxd0zIPPTYmL7R25hnnNk+
lW+xIwFRItQ4MhF1nco2BaOV1RpxJ6VU+6mIXunqU6CQG2SR+gepB+edXL5nCQM3
kQhVzsl8kR2SPa2YaIvm7+1dpkgfRucfBttuVqlos8whYlXk6DauvHJNoad/OK+A
0bazirYqgSD7PKE7NqNvUgXJCVRJS7MtRtL0Xy0D/IdfrbbP+IMErx5+jLns3sUy
5d1is5L7PNwjGJn/UvTPlyEER/Qrz3U6iUwrFvAJUgyhjLoq4Qv6H1328IYHuNmZ
zQlVBg4lmdWzyt58NvPYuxxqCv0idhejx0SxBYvSF2eM19yX4Mni0HgTsFfdfslW
bm5RG24PhO6VJnDjnnFWuMQ4a/VDsawZQ6SkhDb9f9GXFbS6rbBP5EYvF19DbcWO
4sy88d0b9Ygf1tKr0AKez7htId+2AArCirX4/9Ao1gzLRQNJi8BliDhLaoZZoX2b
SUcSTd0t21Zspbjrc0q4iJSSiE+5sO4tikiNsHSm4zU7fHQcCnziMRzz3s0NhaNz
oiI6FBP1bMkMN5a+DuPj0/mVNKeOi1rUb5NvNrkRB43tyrvEpmvqo/dO96QdWseK
Pxg/A+pbHC+IvIZDM+Hafn+G/d4UmF5VVviHp5YqAyydQ9FFo2Dy1i4f2H3E4oyH
ccQQAjsZqaL+SzzyvDta/HCdG1Cugfe2wQQrWh2i27evXtvcDO4AAHaJf8TwMCU1
v1iR8oZHIUVUD+An4OpnCBFwUdkAQxyFxyi3yGsTxTzZ0fk06VxznPGlnVfq1vMZ
Ht797aemXQmmf7FHNQZACkivBl+PYCPzvtDq3ImAPoRKry+jk2i+GZqb25utcmif
GlPuiISofAOKA74nJIgrA0tpstM9Qdw4PjEV863BzEegTCB1mP9mRaMMUc25lNVU
/TojfTmVMH6MH+b0nguUKmTJ/UYAtjbr1D+FuGiZrQFLXSSpTE3HBK9BbE2QG6Yd
AqwNhBKYK0uXvq1c6B+mlUs6aWujqSmI+dq0/tO9j3LSnH3ja7M87XoHNFsvgXyx
cFI7xmUB43+UHrJ27bfmulK/rJ1jMQyMnXZ11S+TDZSBiNoLNWHc9e6snDwdHJHT
K9QDSaoAo7HEHJxc0RdZUGKPZs11S6AkEJTN3ZUtkSuF7kHtISzth2Ev/gqme0gF
oU/ykhu8nOf2pfuyjG7D6HCoXhJRsxHZNofX9pJJeBW/mzGAl1CsBUdjxuaw+PHC
MVMiyX0uYd9+y4xXG1fsK8NcyvkrtO/rPHDHaVPsjtUBlCtQPohbdDThAWI86Zva
RRs3OccLVzOtlA4D3ieyW7Hkdm9kHLrVVZZgTA+L49Wn/9y+XJfSVbheFcViOLFT
8MT/unO22d41aR6mvtvjiNatb3XYcYKGj0SPKrN8xxoONIpLiacgmsyQQF9BMq6y
WMzH1OOZsUifiyT+7odjhbFouuqORUVZ+sm0Tbw5MVuyN8j4C6PbaHvaJHXii5b3
AbOzixCkIhdr2V7kYwYqo9dMkcPM5KqSNFZ+jy8jWd5IUKQGr4SfwPFixfQySuAt
n5x2YwxWtY9jHj9QtWg23j0lVAzM11k1djKXaHOiI6SBCU92QAdpiO5QryOGoT0J
nKFZgJpiUzYzCwGkcGLvZw4odTrtCUuAMeF4sipMZEHS+MKaCSZX/81z6CELvIV0
0jRCKQJn0mdBYDWdzj3Y7L74QDhInKkzPdzORYmgdhCij4Jt5ntlAqAk37Sppobz
SVBB2meACUOqyddedk+vsxf3n7tX1c+Fa6GnGenwzrCa9xpPRYKkXkH1pi6wix/U
J14mHmTyopl0CpxkaouFX6LHlFIqnsanugGBQ84DQvc1ntdidSpPML7T2CzOZR/J
Qi8XWrMytu7SIsdF+W+pDF/ms7KX47AzZGoSoxnEPnohHGA61WobXdRtMjNDZODl
r2usO06Izceuowa3o3HT3pWfifU/2iSK2Jlo3hPTL8WS8bL4AOYu9Vx9zHuT2nAr
+pLxg1N9swW8MsrHbpHrIXDOoisScULyqfNE0mgzxJr+gzZA03hoJckxXIpm5G1B
5EWklP62T1R8KM7i7mLTC65TMVFb8Xpnt08LX1xFVhQx8arq1kAGX7+jqfqWW04Y
2QXrUmaQww8yq2s0tGVkllZKhXtPsZ5NCecgt0rQNxO0l3LH7K4u8v5LBVVijD5z
J7YBVv+3t8CZ9+D1r/w64ZOtd26fZrUUfmn4Bdsxn6hTqrlyAJmF8jLlLMsiCH5n
cnKXwp2C9rHD2bjHkmbtQNjyAY4ozCHsXgpIXG5321o54YIUsUFjmGMLcqU5b7bi
IxrGDosKwy67zjVbPJLFAQAgR2K6xL88z3oWeF5ae8qAcPcPsboZV0DSVy3HSvLU
nkB8AxanUvDLNfyIHTkN2FBSUyQPhZ7lra2PXE3M9xNsdZqRGme6rZtz7ij/+KZI
aDbsGpx+Pk13lq/nImM3KpygAcxwSdy5bV/qH+hkLorX04auMzX5FzC4qbwWyCpS
rrBMuaRPg56J7/DXh04AMnlHPUu6gnzofyxB1+kiQEZFGRSwXdtdjbH/LhJx3mBH
vMrKFFblWbNw0dWWRt2UuhksbjDPav4jzj229X5Qjj/iZBgZVHUeITw7JeN8HhA7
agkhgVSGxsh5sApgcQuYsXLWH7VDBw4ZaxS5UYgfnSTG3kuAzLATUnX71jKL13PF
UB0ppwk7L775W0YtnIDc/KJj1zDw4aRqASQTROpl6KCRe9WlD0NbgwIeF/pBNby9
Nd5lT2XV8uRr0ED5s2o/Msvv1/K3zWMU6Ry613xc8omESHdI08HVARPwSiOnfHTK
pourqhkeVbfsQ+fVp8ydodHKknYrKB/1s5qdYpuwsNg9p+PjUGYkiEUxJIinz8LC
hLyX/aHYIU8iTfihBBBcgthyJerTqn6LCPYDN70zDeTYU1iH4BNmruIcyL4jlyhj
jbzc/761v9RtqMSmKiAiGYa6jXRs6o9kiriiGhZK4CVE1xzBejdFu0M6HyLJa0G7
dLcVKI02Ky0AEh/YKTCfhlGifKXlg8azcDIq/IJD5T5NMIO6vnveIxE/+Fit9ZNF
Gk4rpBA7J/q01LzEEPbo/CqswKJzQch0WoTQ5FyCcvwgG1r67U32gLvHXxa1tgW2
taugyXE9F78A4P2s7j505mHJ6qZoWoD57tQGRDJUOpB8XVusQlX1Bz9hhmP+Op2o
bkfObVn7WV90Cl0dqYzCIE0gD+gUPYU40bH2XA9lvRdGyfiOpLImguEIwfSEhvQ4
NM8YIjWoMj4lg+NxbjnXcyW9xbQj2ZYwtQcPYj5uONs9ZwLk2dxtZd7gE9fjIrzY
BeIkTqYLXh6n+37hJhC0noiLyV4hLhwa97M5q9mJFG5BoS3DZnaSs+Zxbv16FWFo
YxMbC9xWIOXqqQcfKBcEc5HXhoeC7wMF1C4M2QiuJtHvIDVt2MZ/IM3xYFz+PtS0
0G2/M7pvIkxkXZeNuIylmnRwM5su3k8KxCVo9poomWRmhbjHMSp6x/awixEeYser
hamcwEez7sDhd1MYDsQNJgMtnwjypFxSoJDHKweiu2Yt4eGctKXmzfp3nE7t0iKl
XInJkEEpyvXw7pjXD1cDBrmWKp9tvKfRBfA0isbOYDq9nGoiaUFWTINU1V3BBRM/
PLgSr/Uzc/mAl5rd2fZDQ5hQSbZdMuqjOTIIvbLRET74DwSwEQ6j8HrxikowGz9l
3kR00dILzDrdv+C/ru5gko2MYD6vZR8wwJBcZJWct8fNqUA0WZlLPl2phd6pSVIx
I37FFrU/VL7D87+3Ui6f9OYbuN2uLEjpmikCPjab913FfcJgm+oimD6ErgbmKU5t
bag2L9B7PkcAybf42J3ZQ+aoPbCXnq7avZtTBvyR8HUInkI9Aedht2aagvdSHq6D
szwUZNusilokpI7IJqQKrxtexYg7Z34O5LghicwUirTitQ8kwnXLS2MaOiRsFRIT
oWWmaHpp93JMFTOQ1HOCe0CZmT5fIoZfLqU1+y+tooPk3+KkpeSp+DIX0vt80eRH
uYTAJ+swndldhHJzkkrv8JEXbIArn4tb31BPhWU4H2HkXJv3FYjPGi3s68lfATT0
tL9lUnvu6AM63ywvw0UWcYJX2J9kMShS7PU4+u4BQtPvvIpKuWyKe7YmZ06Lgn1Y
rUdaxavvgBEk9mw5ABRn4+Rd9/tlRVsMit6OmfTAOjFyzmpxR/SYCwvyPoyrjMad
VKvA5+M8OnEZ2NyZq6Asl+BUY0sd/cPhA1GM0Mhh82vDvoPlmfhnyqSQkUm/WYSN
rYq1TomBsE5GxgeYLI+lIbFzMCr3AAFi88h+1KwR7j9j8KO2pafjHAn+NeaLLo7v
Xg/gr5gbG0ua7seKwZV5cs2Is/xf92weLkLXXEI2cFhBmHo1COevPQG/OQBWEEb6
bniKcUuoQmZVixoyKFquauNqTO6fWyqk8xA/Bc1uuBeEGYpx0Ryc4/jVC7J4YVvt
s8L++E7SfFlXCeouJNTrKC97EIIj2ZJoFdXrPOSDPwwEL8vgv4irpWIxLkCA4hkq
ydkTogLK3sHba+7sgQGN3LyUZV3BJb5MRSdEb5f88egvA0/7vgC6ZC0qJk0YTkT1
VrBmvpU8oXnTQKCBLSlxyovzKKdwnSf2prwdIcUSMGNm789JiCQkcOcqzUbRxK7X
21+LbwITpY+Qaal4pGxaZjivbmeMnmE8runJUHQZb3gwj3Jt6InC6GPzY5oXCol0
1X/VSNnViwRTvZvyrkkBNC/lVW65gTtU67IBKuMpQnwfHG2FAsgx4mzEo4MFDk7R
2MdyjtHlh4BwmnSEMhs4dQ3dvhuVoL+FHx2Q4xLVlqZZIRHXfyDoLLGlQnr8U36O
QlggPlOm+ybTJ/6l7jE5yuhe6llB92TVoIjzwbKE/z6k/o2lppjp2v5W+BgK8iqI
RMAJpYKJsGq3OLnX6B2y4ls2uIqYD5xGJHwOZMKHLyICXWyjL11d0VqB3u+Z5jdC
MqHpNEneVRaZWp22W2of7M5vqHPC6FUMRpak2BveOMjXVQlefy8rBJk2fIB66uf6
ErvW9R9GwuXzfolATItW7ZW1EquhDx/DYvqy0w3Km8a+LVH4T2hPomKaPSNjot8G
QMCQPMSrYSzXinqMKfIzKFOC87Xo2ckqgWU5aot7ihxmGxWtVfuVYU3Rv/GY2K1U
nxjpO7KABvPK4tA45sZw1O18lgHKlyW14INumBMu5S6QoZ5bQLMBS86QcwtG4+ps
d6Sft6brBON/yTdDuPcrmLVNm2IuCaDJXvwD5X7Kc0are3m3RgwUoU8UbXkImU7A
BtAalQNiT+fav6XA8LHZxbLz0AwG/01TX8dZwAvJxSHN+JnhO5wBzQJPcWVL5Vty
lS18dw3CVf3IjDwZ83JqlupSxO6DFKIjaWyxG/pL2JMJSMhzHMvXIB8H3MwECsjq
tL8UT7g3BBdswPfg2u71j4UExP7/hW/jMzYbZqRZx/Jxa+S2Hv9VreWc/6iAWY2P
umzOXApJbUKcm4bLEmBdtle2rPBI+dJYHgrP8fICrgDkP9g8ECu40oqS7ZHUD7ip
sLGoce68HXb+fXKvjT6ItAU3EhuRRy3E8eL47YfCXIcSLIdtZnFNQ1/hLdD2T19p
VHEKR7/BiQDOGxRFdL5lSo7fqBReVS9Zysn9Ht115Kfg4dvlfUSvPqR8e2P6mYzg
EVCKWuRPopVYiPvMymQjkzWbVR5CbXMX1sFUDwuhd3rRkKeF9RxzFv9g11sDAbmr
qdmB61y/k9cPLT8Pk49GGsJP8tCdg7tA7QTWI4V8wAsC10mDjA/jXWpjAK2I3cBK
2n5cUlW7GWo8LfwKueYkyirEuT7hyJVSH7Do01O+64gFjX5mJl0VbbrluN8kvQB5
A7jEgR6Bw8YnAxQh+7rrV273Sr13P3v7pLZBOxKbUTtyA5TKlF0WhA7ZFeKskJqs
9EwpAxGYq4mQGQt8RWYn/hLiWb3IWRr4zt6391NB8/g1Cl8Xk+C6zzMFiWT1MxDd
NStg7nockJ6GWmTPMtP9oifJPcbZnaGY6QHaJgc6iM7svnFbyfjsi8dGn3kgWsT3
USGEzWPhSjiigN+EAX/xc6Au+xZ2tnp0YjDtbj68wuJTcN+qjsMONmVwxkff3YlM
SyX7hdo/qHssGRtAm2FUF8objlCWp1to8Q6mgmeMeSm8aCKs393rDXAqoezll8Ck
6XjGhohrDDWPNHtLXKZwaXvSmR+WEkpnVbQQyhLmno6WuUanJffWaAHV/c5Ux8HV
Q2CgUnfQnvK4VfeFkjp4i02R/Z+kFM5S8pKW/LTcH4jZ/xC54SDvpvBU39weowkt
aOmLW6K34q84PDRm0J7BcR6DMZd3BAD+YPSLeL+hFYTZyZNyM0stjj/aoalBayqR
Ox9r6ecQk9yCPhtryjyWB8BGNpcPsoo/ScSqzKaBhS5fotSQrMbM4LNjd0j46Fyp
MQFgXTbrmttNUL7VykQEGIiHJBPp4M4lGDQIMxBzgAiwlbpCJoB6cd6PR6EQIfwX
I3WyBFm32MH/R/YMk8Tnb0wRnYg8PXQC9BM++QGOsseAAZSLvnX/2fMsjPeBZG8H
IliNPOemItsyvysOQwIlgb1REJDCzC+aI3wRgJsT/SB9hSFS31wpWnlKCEqPS7DV
rZCfPoH4EDKLp3aWQ5RBN9MUGTEtKjGhIiW/bgrWkJh80DRfrVIhd8Cqc8IdthwQ
GadZEWDcj6APhhFV+cXhPq219K6mMx15NSnixoazomDt3Yl7icMc06J0MofASSLT
MLrXmVJKOEuy1ZFACc2NeLdg4Xa9ay5a0vAWMUYfBoy/FAKELfLsGzOk2HqDeBjK
KnTSCJJVZr1W6gSVd0Q0R22M7faQk7qtgEovo5uD/CFYnqnG3dJmdmn4syKVjelZ
IOz0lPA0/W7sy0GkudG4EP17ysonuetzGWR/TLV0TtqgCWEvfxGGxdigg72p327B
gd0H6Ves8urRsOfiq5vk+FstOmTUHjJ7zin0TnprpeV9muwDsiaxLTSH7Tz68gYS
X531OYjUMTCz6WbJMfr9/xP2RD+NLAWsu2GDRgGi/i5CZPLHXqhxbktI7yHWykn9
DUq4uwtS2YHPDgEkUrIJDCGNBvxzHGOzvhZv/3KZkRebKgj72cfkPQPtVaMEGcM2
EQzwI22/X42c5Zx5+n6r2fqwwsHRbNjUw8GFJx32iCRl/sA0+bSAYdgli/RmowCN
eqSFJvR1jldA8BsqnJQfko9vpYpffSDYyUu7MSAGJmJIDzh8r0ZJKKqAf6i/Djkp
9OD25SjOR/jaxPzvYudVNRwkEpBsOHaWuU9YquJsMOdyx2KWWwPv4aM1pmIqBXDK
b1ooFjjBftxW/yc37lrLepYjBDzALLNWVsKhR58dugcyYRvchm/lSaSPCPioxTKB
BA7CIl/DfPhufnbA99Z0ZUgFjv6XhEtdXd9uu8fOiCv43wEqlLmniIPDObi8/a8i
wLzitu25GIEiJK6uq7D+G93R6h9wdBdyNSN2d6dDc9LBIwbqg56V56BGhIOrY0S4
5noLYCYVGMdRk56SB5siA6qa2QYFnnM0TsrM4Czo12qO2moWFRzgTsc90tWyZL5q
ndkiURiukgobyzGpI7/K11MdzXhI0BV9a0tQfmx71QQc/OxispUwh/ycIjVHv7yr
3JHpwMGJnqMWblWWxVCVbrNwBoGpgUQ9AkRbNpWPcrb6pPbvD+d6sPfYiZqlq5t7
Pj1egFKccNiYc10zScu7Tamtdmgx/EmRvmA5Eg94Wpqm0N/fTcs/TgpWbD3R0GXi
HmPYiWjeE34T4XCi2OD8PeIbr3b9iPwglqCijBu6t7Rvy3lRELdWOY4LdR3Em4nh
dYZy1g9RhG63iwKdZ2y+OkET7a5d4sBK5uqpYj5ugEcJcPWZan0yubO5oYCSpNt6
De1Ca4E5JFKWccg/kxVILmZ2l1AAwIHyyblePtnRM8BoRmQHHZ3PsFKwyi5fR4To
nt1GOySZw9fImIShAJQcpyYtB5+MxZTL/70N/28K1lMzBroKO9ZMemEYIxBBhfIu
SLZ0a/lHI0GI4dLm1sxjXvlsN0elzLZsbt6O8dfDB6pqvF64T+d7yyIPp0ZBq/KO
XaXp3hl+dg00hRNDzvbkbxBsIBw4mmlZDSFv2ZApsaaPhux7tmojXacTg7p9+88X
+bc9sdaDulJMUdDeK1RUmn63RL0HoPLhC1w+BB1MJNwfbm4ZBfLCEWWkswb9udGY
5pc0/xX6Cde2Fw3tKBSJIJCSOInJP7fx6kUyVsE2PGYVEssgYsr3bSUc5sUq9l7m
ZbDm2O3XmT9wv7eXFE5R+2ERN6O7vUh7DkvtQ2mQxFn5N6xdwpqn3OZ7wHOpVwql
wco8UG3Xx4cY7nrCUOyEjPoFcpwWo18jqW2WSMy9TrD6Tk8ShjE1ZLte5YPd7y8w
y6ebwmctuUrHPc9bKXj2L/yfSwQ2M+nVVxbOCyG3mwuhPN5YWtY2G+M4M+fHC4kl
JQEmkjeYp9P5uCFexWrQkl6XjjueWUOhObByYHOMYxy9zEg85QIHMK1X/md4XwYP
96r/JHj//2Le94yy30h7QZXf7JTSpDpUfwhbPqCFQdT7sU587Xh2bJmKEpTQ7t/C
E/EdVrPsQ77pM82rsWfm3ByULrWBsaYCCPEInknfoUISlDtkSodozWnPO7QSNX9k
I5uhYGI3hh9TMYOP7na1B7emd4SW+hYh+mP+C3oUvAF3j0YaybWWmMd1vpPtK5hx
2O4Fd22UYX6NEa1J9PD3dpqajjRh0Th93t9+dCf6pGhPSxPwdmRd9ybZnsUTwBOn
GU+Da2mn+hHIdNjevm32K4dRHU7qpMA2JFDk5MVo3aXWmIm7U3TMlyO0lmMBOA4w
rYHWj4iPFxBVXZMOCsYIEOY9F+ZBA3IZ+ZLpLCisKXX7/fD6ggwEGXw9u0GTMBZ4
D7XgG0gQ5Vp6OF1eX8dazXSwgYRh0BgVz1A5YYjzwtGX+lUs3+UiB7Or1KpIoNyj
aW8DYuH2gFFrVcrpaqD/8lK1SnqJaUL/dKShEft86RwfJsmnAa4OOqd1rStL1kMa
UHXJDOER19Tg3PVeRkLNOrIzzWvspir2ofDVAIF7znVEAtpUiGHRvv1lMJ6i3uZT
4WsymzBxdo3qMDkWsk2CI9pqxFQ6/2tWtUj1nLhQbBubI4UP2f1uv8bpFes1+Iv4
u896qRU4JRYS7p1AAS84ovF1eXQ5gafsbm8NtflloyOHfzHTF+Shgo2obiaYokIq
SzeIQFZNOkJc10s9oCVbgww8sZJlP7Byc957ZnOHMcPMUK2IonRvWng7X25z/tI8
7e4qrF3JN9BsGCunWBI6Dxqv5NzOn0e+G3Ip6hkeDK0aaplDss5h+wUyoQzjqTZd
W0CdRswlD7V1YDUDDN4mtshj/kpExOzCaEnUCOu60zvJD01/hbslskfDCennBfF2
sB1HBr3pwiTjy9n+alESzVBWjb+gj5xXQh+yDjPMpVyWlo4z0VvS8poOirRsdawy
2vuv++a3k6r8/mTp9Nq2ewyFdGmY+/glxK4a9F23D7LKhCVK5du52BSBTpBHAwIf
T7WTDKvV7RQ9GbcolXTDFZpNjjEUfqOKqCnn2KhrnBcfN5QH+pR3q1cgxGj57Rd4
+l0sIwrBtFhz693L+ooIMWInIMDNPN9KD9VGwMHrbnkTxMT4DeKUYobSASy5f9aY
OdIN4iTd0EvcGhx3FutxfsMYlV1AfapAzlfoiUbJBgzwS0xL1UfW5ocHG2PRRS1Q
z3opOsmpXKca088+tK8E20O0ggQ7zE6T6QwJrbL67JoIkYty7BrLN3TXjEof7J5d
RCZecy3ZdoUPu8Ks+zMqwEVWyPkaXbrAtgtBzRtbLkSwcjIDT5w3nJ7+wSzmqGsG
vCwhryWtfo/vk41kNvWH+5eFHR7Y4kBO8bzmYEG1LkII2EF/+SSWcNAkyHA4CzA8
3h83Ffwa9GC/ps3achSL/qGrd0HE9xbrwo9gExwpZ/+XRhKQuqtK/vF8wzfPZ9+r
6/Y8TRS6LzJ/9Yet9qiLq80zK+FENoMrbq6UZVF/0EAi1qPVtUiVcQM93mBogzVI
Xiii0N9aD71KllJ3nDIZktWAv1BiSk0UMliH2aPWpyOLOOK5Myt/RSbiRg3UGWr7
gXsyUGKd5ass7bOxg93iRC34VSgXR6yLsKGSLhzUdtipzuYmygRD8Gz92v5lBmJ7
HreQBsIzC04khJ4RcZnvKDvIxWZoJT6Vo6sOGPoa2M0omY1HLj5v076TIdTGsKYu
Yy/AKRvCWQBoNUJ2Qf1rsPItrFSlwcB3H1j4iRNoYda5eaQxP22xkZ5OIXIHT8sk
Q/iqpugiX6FH5xvWPySwO7uSzYaIm3IvNst7zvuEebpVX6KpEABhuCSD//ZoFyzQ
+5EMs0Y8S4F4AK7AjGuA2n8EcTuqZHRTSLHBC7pb74C5s3rZek/FfW+SKoQtubmr
HPYDhIOSWgN4caO/fgRjeV7c8SehLTDH7vHsaPFD+aeNDdfUfyJT8yX/8I6bbxfq
eoG//WpIm3S7fSgF6bOphQIUDoXCn03QdwAt14T3URZMYITQi8TyWUoGDUM5oVws
stUepVmE9EXFoDn4IPUmD43fsTkiFWrlgkNwBebx28iKoFqHIR2cLpNZv6lMEHdk
mvuOyR94Tx1NntD1GZW8J7xZLu0qGRnCCJQpg4A8Ipa8V6s3/BTaI0DjASK6h710
hWEDxs0s6hqKPB1HyFm+wYA+Cb0wFTAOLvoxCqnqzpU9/I4+lutwHZ+b90CJrjwX
646h4vniFi3Xz7mCezx+aHOcJ44sfncSqpElg78a8TF0O+jwCs/1+5A7UKKtSz76
FINr+9G9Z23lnQzpFp7ETJzdqr47ZJnbGEAnh5j+DAMHqkc6sThXzHSi5G2mgTbv
WrpBxdpzlIgNrjEv4dDmiXUz4Carjtjd6dM+ylMJtxT++XNvMhz1NGT71qXqWiGi
zffHg4GzfzwpfcBQc7UmL/J+GGSTYX3lb/l1kpLT1m6CmHH2geNiZUmBWKb3z8wA
NX7xYwRSK6PxTOcHa4Nj8gyU34CqGXICCrETspDA1rwwWalBZeCSElryd/oDD70h
PlnPfNYB/ihMzZ7WbfG6Qq+tDDN61B08bJAuTnKLh5LZ+//6jf669MaFkb/7BFbZ
0IMxUhfbe3v+KSZLG3c+QcFGDPpU4Wz6YKXHmKf3c9e+jzb85/JxgOQmvMkkyr6r
AC/PzU4eLmA50EX729i41mK+i0VIZPq8dsRj8TwWacWo1apXph5YDj4aZjf5SvPw
XBL8F9p/Zzr8eHlhzEpo2bxouBcXqbG2AUBJbhnzuD3we3dzcR7xqBtdn3wvwZc9
3thLfaehjATv9Uo28jMUTY59W5ckxFpZpQfER5X71+Ci7wZtOANA62DnMp0hRcix
wT9zoLdpuD3fHoZ2Tc60lManqHfqZ7EmiJAJVvFGgVk46h5oqryIUynu8W/ddJUD
LraoqTDTaKmt90ZSWswFFRmPq6Pi9R61a8V39iRnw3KcaGtOEqNkf2SHYm6g++g/
KP5LYDQtm5dKImzOYeyOxmW1xW+YMUvE/I/a7O/8Tc8sXhliaw2YFFl2oqe4irG6
BQcnjqC4b+lQWq+PbcwhK8tuIBV+sGdCaTynACKIIVBgHKlR4WsD0E6Ogn44OXxO
uJVQkW+wi4DVrc50/NkyRZxH0ZWEZRio8t/J6hV03O4j+hQt3Ai0seImdkZ6YgCH
fAv6m8aXiFKlUM1OY2IFkSt2F/ldhx1bdnQ6A3fcw3lNmcxCwEN0zCKu+QmUnQr/
8gaVdAVW8H2G+N38kGwPRAigt+mRjAJoP6ipWhDSekZscXlqGI1WYkXqLT91o4OA
7VI/NXgeL8ofRygBddJdiUU6d58omVjRXUc5imWqlxS/AOuGUzSYL5PzuCyPrVOk
R5t0iKEyrkOnC36c6PowU+yw8KvQrWLvpX0j4JFh8NiM5ZqJRQ1x3Tx+GveqDQfJ
q7eG+2qdmg/oR/iYPU9WbwKsnKQVoqhv3Qcl+cBcxMGxIrKBb/xe1EJyRpUYXl2d
r3x2YR3B4LpRtMVyWNM7j6ziglf2B1yh8xpSlCJyvDPTXxbOVbnSuD0o2+Yutp33
W0BYEFmnDbFPTjilmMuBzeG0cMtEqNw7PyAR1oMetX5pWH3aLUxEEEVr9EGEmNXM
XaYXgcWPmFFcjovrzjoGzhwjbXP6Vj8XOHQuri5spZZxqK6zm12/yhmCpZNbg26/
W5HOg/JehKp7HsuSKO0JrUfTCPGtYVBEPOXyh6H1ulsZ4ellTSXRkdQr4f0bVnze
to97NOT4gfYXL9tjj7KUb6kqh65NrfItBEQMGo7CrS+KL1aTkzakzW3rehn1HQAq
rTWp0SnanvF4sPGRnWaPHlifqIITZR7uF1X+8OZ3ILRajxp7Tkzr4+DIY4RSdCqN
Do22kI/QN93Ch6WsnRB2QPffhnMxztNAnVMlNrWYGRmudoxZ8mjQpqDcyBudO98I
2Qi43RS/DolXix/Ce76FWIs7AemYpEmpUXhrAkG+d87OnvShV8s7cGAw5NldnmeP
/iJusfBWkSTdDxR9Pj5agAd+6DxONx0qZokAi3zpFOaQGi6430SRfTH8wDnN+4al
eU40lbH59b42wCtKvsnb9DFh1NeSUjT6jcxHxzg6K+5hkAKdfdwuW31ea2spbTPI
tDIFS3lwJq936JP/+3I5jmse84aeumCEvUKUTWkTr/5TE/bJrF00bRWnkSRaDzv5
zZhSzhV1/w6wz5DaE3nHcmbX76ffHCHMv2L9QNelPV0vbOCwZ8N3gk9KZ5gaVPom
NEf+BpzlKysNCJsdkvEN51spFn1AsqpcRrdEt6nRN8UZoSJE2qnrBhAtjM4laZYL
3ydl7EdKe7VZkoPHCKeKj2FP9zzPTWT2YYeaL/K895un1lR/IvHqd6DgaBIdlTsS
cxQbr5QtxH1etUBjiOxtw43VU2ZzKBz7ht42HopWrY/+WzgBYZ5u39zp/xRh/uzw
SFMxNp86uiWF7+NUutWTeFRb4gGB4ngKDGMO0mF5wbi5da3p7KZkGZb4QawxMEbM
cepXRbIZMRhooad/qlIviwFq4ROarfgW05I4cwSqXAkWLW4Xy9kbvgTaEdEClvFP
GI41uhPQ0GlE94nUGcsaI1/TYnsoQUFojdSWR1T5wT5i91J25RyYWsb3mQ/dIbLY
2lhN1GhrQ3EvT0q8+s39BKtPtgwu8Pb+trx8MrlOdjilkZ5TsNb3PHuzCGAtG2I9
euXv/1H9U8ACaaJto/a1lQI0iB2LS7HW5Y33oRoYYzybpSfj5PQ0UHTRVUdKvAOH
O89xos8iH0ofaF4WJzpjd3BRzsplbLp3nXOzzuxorKu7cfFdE8ih1QuBM/6MOElA
NKgeKS5PF1aVqUVG4U18TClaH7jJXTlWOxTqDAIE8WwdtivHwsnFJLmrsRK4sbWg
bau9GU67y+aQkuoCublRAHp2qoAcWZY4KfdsAZsgVuNlRZe2dBbIPh69+tTeOxuq
ofs3TsaoTj8UIYUDOk6vPB+esC46/O6KwSW5L+5BB7Y0mnjOo8jigYs4p56h71RX
JGv92O2RcdV4ReNthZQdd5OVp+lHR0ScsJji28F2EmJSoP+ZhdvXAzXDbjij63pa
3e4FyBx8bMhLOLtyI/l2XlSj5FyBFlZM7MPVhMe5rqcTWA5VwKw9HZNsOVVWUAhK
G+UZFjiHguO/yTDOAtYF7whXd2+TUxbiq49A5QrSSKyGt6flcz8wiNovBEXWz6ry
G4IzBAqPnQwfs7f5McEEDvhgQmPZgkG/fq+i7QHcZ8ZxfYIzvb5WT52eVhvyxHDG
FztihbYi9dNIFcMh7CryY2VMZMI8DVs5MEqHs1R87g8tsrO19tA7+3kkMaUX+ZAz
tpRWxjlRihej/fAglMcTRpdBZuqNM4m7rDgseWej6P5wAB8q99lYik3fbwmfDQUB
bsr6QTay6dym/XUr7EukdWjs45ZbuAM8fWnjcCITgAq0/a+qH2YhPxAtWsA9rHUJ
O6/NCMVaqhriLrXOJBb1c967tkZYYi3gKZOil3h+W6EDPHPvt/Vcw2G1uZtBc7Sy
q3VUEC750j7SvZ3bpyH1LDtnTb7MUJLdFwm7+wJNnGcfsQ/i4Xf3GCDPKRgHb3AK
wAWOJfrVJAK+P1jMKiOxyY4ZY201XDytvKHwcyzlv46MaJvFQMM4/6LwTr2odxuR
V0bFTepKvVJluKfIkoLvgqvJAswcyUGEZZL4Sx2H8mOh3Zcbu+C1jjIr4+lxvff7
qIswNxruC+vQC1QN1w013KA2LhkghOQWoo7tFbvfOyyqX645QU1YzkuLOGq5I3Bj
tsJKEU/kQKCF63Nhkq0eiLMfeXOPA7stx9TxgLRpl3/ppl9NG6k2Thhm/vfLPCDP
6QP5YMKoZAIY3vks0TDmAVxodyC9AV6ou1UWVYh7g+QOl/V1Hhehu9jRreGVufRB
MdLOeYpMyubS8UAxhMNjS4Q7fa5lNbZJYMUK8zz0+tfdeFuc10PxrgEUhGJp/+N4
w3bEgOpd0czOGZ9zbfBo23lolQZcPBmLFegZ1cqffQaXtn8tAAY22hwh3kEyAW7U
q/DXY+f9eg9wLTVVU6j2SxYSoAAs+a54NUxNwOygtRRiRXG42RzsRlOsrLi5HTIg
BPJv/dc59Nl+xeBuBBhH/1rN7nFfS9alvU+D1+/VJB0K5nDMsKEz956qlc8sghF6
/XYh9Cm+CpQjMl3GP0yzHtuTrloE4GM94YbMfCivn1In00wZRCPwT488xlQ7RIR4
9VZQnp0GEUgr147HA73YvXBefZ13S14V6b4wmahch1vgtAIeRj2ywK9Vl4aBFUGc
8G3eMLLPOd4F6auvHdZ2ePBpwLe2Cds0E49cgWbXIM+WgGezuu2pN8z4THUGGElW
L2kbtJY7xAKxpYfg7huRSWhPrhIIJU3EyHoL9BvotuYXe3zeUsnaSus7QUGWAQQR
dzBnHeFEzSv7ENO78sZvLTz0CSsz+L7iRgLbgFnfvpsDV0Lje1eYq5g0HSVXlrSh
jK+aJX8AW+wO6rwh6EJzoeWgGnalNoEBa3m/bQcL9hY1qwIwlXrgw/3H2lSMxzEK
daidpGNQbGnGkyR7dnQpK/2G8GewY8KZM68qD/bOJ6BOWebKGnW8VpohQoqwnlj2
qN7TIhWZYtWEEIHnYqkOE1D6RY7lkXU/hc8kJDRtn2A4cCplvRfTU7QBZtQ2myKi
q8CYQJrZ9FiQU9T8WkVywTpW+LCsj1itJMWUpqiLOAaJSra1wsSN7Bl6z5lHvZE6
YfCt82zL/t1SGwkCAx0QDkULTuc46+J71WIEZH+6ghYbRNbZdMfXYBQgKQcLxkuv
0WwPIJmvhiNm6iGsYVmDfINUgUjSXGmws/9kLiXgIHjYW+1PnNX4N62WMoSQGZhe
WUNkgychiW4DryM3i51SR5lY+Gu38YKUvf1Svqi0R58nrHdKwtcWuHOhE1wmqocK
qSMqxBQGpzbxcV8r8NLB/hVA/UBI69D15WPXp9K8vZunWtTZn7LotfoKq97pDGmh
w/fzKCcotXzyj3DagtR/9SXT8Ps327om7bsEySzNngeyNkrX0eQdQoaBDnn1enRl
86AuLczqvamO+nwGZ4fpA5ocPKrVgvfQURYHsYb/bJ2ABz0sLDcg6/fwFxcMXd3W
zDWVLJyEq0hk3ccMSBhbYT5AfdJxThKiF/L7L6aum0d4Y0DNp3f/1iFcwfyQp2ug
wMma4wJX3V6Fs8SapyRQwK5UMKu8zouk/zrvQscpfjfVDrdcWwjC/0v+bjMtAWJa
pjYcrtdOPk7wGANY49iVSurAteVmZGarOmBEF8tbKJKo2ckC1n30BEsUrixzqmMr
c6S6y7P4xrkLad3roBbunl9yHEwrSmNwuE8uz+6qGz4OrljeNNzKwZBhlsQAgbYT
WN+mW5c9QbVwT8WOLWjhijh9RolycsR96wpZilGn1kh9ieryP1yFtDQ+aEVxc+UT
tQrbWiYeVbuYpM4Yz8Zf23tpceiD4v9JqDsV2lQRn3tl61kNOSjEbQHbWV5wjS23
Bzrs/grydmphRk3y5XdhUqKTHdXzmqBBri+BYFsyt6bBcjg/tKIJ42dxsM70gf27
oQmgO8yHU1QTPYG2OwWYGLDA/2Loxo74xh2hOA4TNWZfANq/1JWxrSWPdXQfLoQ5
MPcJHrtgJLOE8SBOuwpU/NOmaxomazJ0HaAnC0hTKmFTFVkwG7JVFtpZzRwHDPqc
y+0Al4PMndacC6pcaLS0LwSH5tbb3peUsGT/oQ460k5exmnPV2bpep7/OTk+BtOE
8zD0S+E6GzAVsf12WLS6O+eeEbGAtLw5L7P9DAJnZ++UjoxH3xkRoQ0gWzKViHGy
LbAucmGgy6oG20+lgLvWVanELYMS/jXa437cFYud2gTgVvMjCdWifRkBdQxNMPM/
VYXgYnwLykgl8PhVYZ8RwLUoBP8F7D787nCdntNmshhy/4+B8dzJZ3kuQF2iIuTW
zUQCyCdFwoYjHwHBNWL6xCM+Kan5FBvvjGYERX4Hh+3xUd1Ma+ED/GwnnumdDqgS
UTCOoKw5HDCjgm5FeIqdkQRAZQ0/Obl4nAjujSCvUagVgZQG0QEx32isbklWKNz5
nsnsBD3Ft9mniFUCXC9+cfnQypQLRvzP5uK9tra7eg6LXqPyXraK42FAjMNtYCsS
+xl46NBDq7QdMO1B31JqCy5/wWkM/aN4ulOk/3N+pEb+CChVmMc+tG93AetfVafZ
f8a9ZToPUT5xxQmE9yYwvnccStTv/q3MTu52Tmtg111ZTgvVR/gpa/+2s+9MGf08
wy4fAqTcT25a0txdXGjNBXQ3+1Sv1yWZImy8tEyM1gWPrgoYC/MlteZhW49gVdsM
w3n1dTCXQ4YE7VRhCLGuw0Ars89jQJcQ/AJQ+h2Djl6QoidrcDibbrrIHyQlcL1A
kqcJWVOSJ2lYS8exj85BGUdWQkS6BeZSqqFW0qQpmWc0Z9a/yStI54P/3wTVJjU0
qK1KY7Om7PTBTAaHrKCV0IsZYdPNCSUz1kK++A7AUXHttVjp2tA5AkNyjLTlftAI
9m/T1DS2CW85zBzpZcxobGIWbrOL8imdjiyvOhnkWtdo+3Lap7+2wslaIdFVU2oB
SpiISt/rKqft6UdMldLRd2UBLvXPhkNcPSXVFFZOlFJcaw1I9gTC7KAEtLnCY9yO
t0jCHFBirGOlOLV0D0n6GUNwYRxkCqLVQTYXb6Gd8LkVi+glL2mSnte3cS7r/6Mj
ygi5yPtKWLJzvNq00yGCzq20U0ESF6d1rkA5PMrGyRFp0jokR7sLCvoD7NaQDUc7
uXpDAxQxxQo+LQqTfYf8crbPSBUv1iuTOE9J5hGVYQDw8dGpQHDUIbnh0hsc3Mo0
FvsgXunjlYofC4lZED4mXmr05dA7LE+40OcjpxfSOOF27JKQo1jQw3WrZILTyTJU
3R0O7lCo2RQXzpFGB9NqqzgM6OC01jI2gedebefzFuh0k9MIO3wQdHH/iWhMbNCc
madbMkEWqArqFwtLYDzYyEbUAXLDvORoY6sH4sL1nf9kfRiDj59qxWGCpPqCFJyw
UdhkQtlJ/yEX3x2deQeWccLxaCE9f6tbwWdMGwtL4DcZfr+UC71P1GPy1O5hLpJ8
isc1xvhM0dvyUWuwFiKnzqGtnn33+XmRVon7woPzvzUHR7RfMUpla51QsRgdFcZz
N1c9i7z3P0NiMic55kbezOe5E0w+PQ/4/8XH0Xyi188IAbDBmulEbbvsN4buofnz
CDTfmOCs1SSQt/GthcPA/kHBAFC3DX7FwZs2DkIcipJrcM63Sqz+WXwveJMISxO2
krslePF9sm6LGK2pw4Gj24tQlMuHqVIZ2TayyUrfKZnQ8lu/gPZ+2HK9R50ERb3d
nEb7ikGDCNJInLgQ3W9tRWJke0qA3kaqplD/3AWGnilGfW3O2s/brYlVUF539Nch
ymJ/WgW5G/U8sXfvJAEZSrd7vC18jdElCD4rDTNs0IWwe2F5fHmibhHalPVolYRo
v5zEyerQGlwK2U7qBOgV0M8K603N4t0kgN2/QYbO+3IXDHd2dtQVWcO14HuaZa1a
VebE0Tf049NUgnvQdQTRKQMo6t55iiZPXOXr+hHe0pSqST5tA+PIhwVcl9if1Iks
4Mdga5yHIqCWhPHBToY14QxMtsl9YMyLVJN6iJV/5nTFHd0W6HQb+A4q6Nh3vGDC
Kr43SCTOpX/pEk595PeHA1AgVgGk7b+4x5zBzGU9eGRX2QC7JFLMWG9iEcPR2T04
E6epphOlR3ArAdFX1mPqQ3GpwxopNECCgaEX8QpXr+RNB8tk1OROSF3Bp6lakgih
zxx7NAYJSGt2p3Sn8mnLBENrlaCZER+oCwNJ2mODfm0zjfCkBd3Lu2+NCkLxObVm
kZOq20z+mvC8PO9eKsKObITwehlWrFENrTmlrozPaTEcqEX1vQ0BCmM0nf8ndsTQ
9G/dRasB8kajj1SeeoiMaQTEtSXAeLb72avVJncFqtq2DzClro6U3xOiYNFFYKQ8
E126xS3M+4FnclvRtjLNw6/mHIvNSiyw3ci2FV8/1PcMb+8v485D2b/T1FfHmyrp
RZifoGvNTp07B2/4hxXP6oA75p2DLSn0Lr9HdIjwb8QVV6gsl0tdu7heF0tywzlF
iNiEW3h7oXCjHBjSxzWdgfJaVtZlV4UX8HYQPsmrzwTkn3yCI7TYii4HMyOfZ8uF
KYHkGBBhsm2wnyM3rtqRaoya9gp4RU1yP9xPAUcgLoJ3FiVV8rMGpRyjAPKxZ/5G
IHj6LybIWzz7Dbkwcb43KpK3s3rwpUWokFJ8eqlfrOUxwwTvEGOfOjsRXmtBJyc/
j6DIQ2Y9Axfp+SRnWOPxaw6AAqdbcyMNn1wHyjAhI9Ghkl58ELPrwiKWo560i5RZ
xHV0v8NZdvCIqgJ5nJ0l8GgVkadBkgd80bbCesYo3KUPlDd6qIZw6FEwzksTKylQ
zxX3oTK9Z+PQOvPM/B8BxsRt9bsW0D0S1NSw+p0LbJSF/D1pjoxICGYQYI7dCOMR
UMh+vHigTkMDtIMI1DcNIjTCvm6JVz18CTOOiS+QrxHIJM79r9SfhVjquloZsI+U
2Re3vP7qCcBJ2OXGi1BGysm6ZRYbDF+LIfJgr/Pl3b94GKZ1ATHtFK8Myxx511wF
vXFwCF/vYIq4MFiWsG9HFkoYo1O+B1vSp92Rr2qwjksTrkmCMlFWfkfjo5HplcGe
Y32P9+JbYQnJGyDD4QLawlZ2MYki6GVVg+rq+7yz9W8bYQwK+WZNmh4uPZiFqWGO
u6r2akEE3YX6U3seARc6X97MOudTrvoFE11kjFiQlX084wfMtSrp6jO3cBjuCpL6
jt+oUfTBnZ8eogjVrHFXWvjg/jqKJHfJ3chAf6Pud4299KJ4vFwHNlQmCPE62eWN
1jLmbjayHB6j5IJy7YdXSASbThhER+Bf3gldgGldtMsPg0o2nYYPcn+BzkPxApmP
56cuci46+FmvJHoONZQtljFB3fikKMKxP+FTiMuZ1ISfGKVXJZkaE18Ivh5QVKjI
Tqhe1PArrgX0VFljVdZPXIpxAfDRUwbDhonVbM8vKM77/8sLtQCEU8Fg+SONMxL9
h2E4opAJqNR8QSlxKGwtdhFQMQHNjfsOajvU9eMhox0ld58aiHwTotpU4xXpwXnb
zKQF6e0uA6EeIcw0DfTLcnnz7d3P1X9l7jmZQhBuyvspEbzCBq/NTN0R3AqWtCU5
zTguCCj2tvLLfLS1Q2D8KybOlit/huRaFhr7ICnTF0Fo9dzPGaIHsL1ehy9oBUWe
/K5u2gWpXLLTZX/gFFJXe3ZKTcAl8Ti9AvGhzaeY3Cd6f+4w0hkgQ+0BawAofxBO
cHoyzDdP7W73vlBxuF/Mg67nPraimYosxJxqqmE0Ob1cGwJUVIAYUU4dUqajnp+K
MfNL2eSXkKRLDnGU8WHV7fgahkq/RYOmL0dAe+mpcfw43d+XV1Yz4bTbRtl4xka5
3WYmiHfEgvR8846pbXQqXBIyBOOEKtC+HqJt1rAau7bnNAkNmcXKFisA1rQxZLBY
Q4FV15mSqggzo7dg2nhijrejBMvxL/V2G+CqzALph22gFROkIDZIT0BC8oogw6Ku
hPzhH6nhwgLQtMZ1b7AiP26sCT5DBqTNc9UVfNoVjLhIEcpcYNGY5HzQ/1Vg3nSn
HZ5GhOz4PhSqV/EFvLHqZCfOpbe8pKhQV8Nrsm0LgDrEQmxqWGO2m/aZUVt7eGTc
XXRnSxHUyxfsvDR8eAIwTeuGbSqvVdgNzaqMP5Di1aS2fT3AFYRpOkn2lvG4NB3E
Svvf+ArY32KkH+0t5Vf4VkhUI+KbUs2Hd/ftgb4iBPCGoX+o0CqhZE7sLjuaGQLX
CmHlXRw29ZKOBf840HSOabg6+jmU1lIZhblONrnjnKSS13Ia9MEaFVjh0bkno7uy
BlHDd86PajkbXoqp3G3uBOgblwo5aBM1qnt26myDSa0RZOu8P8NqUKn7dw0fHNQP
Nve+Ge57Qg1F3aGjnxn7R0xLwuc7xgba1bjyb7agz5AcpGKJsmdJmJdpuQ+cgVLg
gpsiZKatmQKXU8j/80ZkuYBksItQWde8bjm2iOI6i8lK99PoaDTfAAyRh2kxER6p
O/FcpW+TOPuc2zwtZQRkqVxcgqEKLQShvfV6v0breoFjNjKiHAuGKP9uaKQXyYa6
Gv+6DPAa8v/f9GuAn80LcmgGK1d8xT4xzFDtF22iP2vnEceWGZ5vVBpTAOJv8H8j
WKrpdcuHS66AwBehff3rqZdbexPdAJQJY90726wy7gH16vJ8o+t/1zpR6cFvhOso
vYVvBhJXoQWWu8ADbtBlDfb4sPEiuVfk1t0TwuzVnj+GLf+oJjUquQtsYCQhaGOX
xeEBME1ydgRvqWGkGT3zS9UVa7lHbmFZ1SYL7tHebP8ucB5chY1iSLSj6tdm8FrR
o2bpwygFf8lIz106gdpAWkbJTKssp2uoSN6up0K2d7YiSUrg2zO5f3/8QwiKWUaI
4B92ubeANU3ZP2rlm+pco1Y4zXzlWfZoZ2xNGuPdIhBm4HEZg2aeDLByayJMqzH1
aVVzBk/eziZOZOxznGeQ17b1UZa+sPc1uKe8EqjKD48YRXxGKRE1FLhWit5qkmQ7
920MvcpzrCTPaeRJCXVIKZt6uQSzlttwfcUh5C0D9Q8KRSQmY7IYlluxDkY04kOp
m3YfMq+cAkS4snpPJ3G5Xg5Gyv9k056faE0d5p6TEOH0RlIHewM5c+b2Ee8KB5NS
ScrjvOEjFTsSNvrdkEoYDg5Yw8Y+d0tKKPzBnEHta/s3c9AsYiyyI/OJJl80FIbx
Uk70jl7omf2L/TocuGz+MwH61AG+Jc/ZS7GjNZqaGGMVurpB4qlnobbZLkkankVb
HDEs+/ay1PMYCo1iKHIs9RkLaxHTaciw7wxeqdOboES9BdfT+vaTDgtHxVaWRZ6+
p0l03+ksOgqCSEcBNuMYqsnVeSbFf5Hj+pOXOPfr2drQi4sIui1aLrtGyxqnts0k
kOJcPmjFJiBxkqK6GN2sEbI5jKjAQ5QyZ4P02dD5Vu6SnkFaw3VUf8rXvwKX/L4a
ItC6RctczSDDVSeVlEHM+170bL1RbTPRGS4aAtRfxp083hXEPULykihOKCWjt21/
XYy/lOJAxHMHZ3KmDXzq5BLy2hMMXT7m3nOTDtyWDGypkqMIs+oOoN8cEf/eeXaw
K8pnRLU60Uwn92YtHzv4i4b5Man7sdOHF+tpW9WwW/njlNDdceMrBkkMU1p+1epN
hHy/9FzUiEtwLy0nmWUsuvvmExc/jtjMNM2QQxc1PM660p/EvPVdI8kT64EaAHX7
MIHrZWE1GUtJ/SgOArZKTMTB1owjanjF2wIzlqvrf/hW5DlDlL1v0VZthe0r7K+Y
rLHFTRLUys2g1pf76k8FXufIun6h+mj2DPWSx7beBKHY76wgmZ1m3bgDRJk4CxyG
1b98giMZHD0l85n2yctcFuDK3/f46tCigieBGp4ivWEtwuN9GcdvjH6tNSg9bvEv
ahIQAcKfBMeuJt7WdH6ohi2NNYsbdGjLe62/nrvTfI+gkkE6iacAN2b4HnxJn3Pn
pnugWdiVbZC8Jcs+fRRCvb6Hm7Uy4ok/8g9FVt/cTlXwpc5VUvA04cJITWhoq5qY
9dsu4V4hnJDLv8gDbl2T7EuoB3O2dVFgT1Jzm466qz09QC8EQibh1RODqAa06BTI
fopbHZEYj4U6x4KGDYtjpClwdG4KtBa7XIUrGToWDWEgBveNdrH8jPvarpdh8W2C
kFfYap/0Sqkq3eoe7XFZ6fIZ2qfvOn0r233nE+Md1fb8mUD3+cKtLGEYKJCYjhi4
n4V77vB0ZB4oxNXqzDFeFErMpToHQXpwDNzov2ApKWFz046MspBhJ3eIjap0g43s
uwWyWhRX59ZEAlSmqPVAtVNeVu6Q9y+AUm75Shk7T4SOjF7+V0rsaAJMeHaQQggw
dpFRpZb8Ar/GU6/6vo6hMth3pg+xqjLFN2yVfqwKu3qWrN97hHRq5D6yfoJW+W5k
dQK6K6gcv/+/J8v3UR6Feo+DvuxcSanm97QVb2HXGSJ0O+xq2OiYS+vah33RjwB2
6H3eVpazi+RhQ8fY9ShGbnKUrrAdO/kynv2Yi5fQ9csiDrbylVDoROeVqxC6QZRV
E88x7tfS/5+xVstC11DLucgcUaTuD58S8lWpc658cMc9xK6uMaD9/ZoMdnsZeZec
n9SG2+m7/3WP57kLpr3K4fZmJ1dd9K8KJTmmfAcua2i87wn9+tjGxi2dD3EaQ/js
cLqqXAD5eAwkH1+38TPURBNnsvb77Zz55/EZxTknguySjtdXTSfuJroLBbVY+4Ox
pRGReXkIsmXNEoClhase2TqWtF63utrk7wrEsPJYGL19yILReRd+m9mw1M5wk6Sa
XZEWKseiDzcAVQPvUsI2MaJr5Uh32QbgeVhJNlGS+dtttiLrqXoiDZVjzkmdGizs
moz49nQ2Rm06rnaeoBMFhQZ98J/liwZrdCejI0hR5ErbLtpD0ZReRyI1zkXoegnc
mKU7k4qktUfLF+lWIEBNucF2BomQdhtXRDDGi6HjizU4Pnndx2dZaxToCnKTr7pb
eOFurg0/vB6PEEKaw7VTY7L0Tf/Uwq+LHxJBQXNVPJSG43EO1oyoJTJVv1NHv/p7
WAbtDDTEwvJvYw/VTUry9Bz4JckoiEIVaOsZLFjZSrwfCM/Zwn48ryutLRsGv2Ug
i1IUgD7tJcGCRdKzvdRrxFuY4ytegX/ynLfyNVJlcPm6zFWGt73cdtOsH6oDQJE/
DEjZAaMlWN4rFOeYXB2Ck4j48prj5XxhOYH9e8hiYcWrVYGvlCxjBaGV/fdR5Zg+
I53CCCABTeZgJq1pAiKzsAVGh6/2oQehz5NiIXZbJTifciPhQRiqtevs7qIv0lYb
MCVmbCdFAqi088hlC4/Ph+1KjtysOA2dcIMC+5offyTpeE3k2s8pfSfYnR999zGD
SOiPPgXArh4t6KCO19zIWpI6t0u6YPU4lTzXPo14yfajb8ZPVGQF99DPCKpAosOf
V19C6BgkckvSXvvfEAybHptZYAx1WPRd9KKlr3ZJP+wjHW+Vvz41BBH8z+sW3FFN
Fu3xE4cYs9DrzjZopBz7pCVdAUMNmO6Dfww9edXudzUfDhtpOpEKNKF+x1UvlCTy
PRaR7tL8kU9KQKrDE7ckpVrbt3g2OgXAwEzsQhb44usP2DpjTUPnK7FUbrAs5N0m
iSotM5XGWDY2cVEMJbYB8Q4DZLQ0ZGVZnbCDUjNBHvci/Uc+ioTuKyk/eV3R3kVQ
JKKJ64PrdYV76BaZNo98UDCbl1ZUFwB2zsnsT7p0gWqEm54PXusS8bgWgmkbPAOd
+gUMI+Lw+f2JEEZpqXfFtEsc8Tvz6fbKwIdMWe/hES5ILoBqb2+1XWePNSGga3VO
ArRrBVKLCHWkvs3eano0EUD2RqQdncYTtLyPoM3cgqkehmVm8Kz5QpAjWd421u5k
ZFtygT01Dd7f7zVOwCRiLKVZXrtUayP9KTF7ew22UavabA/08cV3VDF6e+5gwTia
XDSXAALrc+QLBXENDop/Zn8Xks52LtaDBdraH5LXdwbDC0LrkyB4R9rLILPfbydK
bF2PO4OMAMiMkpGOBSVMkkPvI5Yts4lop6wzfrickegUg3em7YjiVdLANbMBOi2r
epXC0q1e29V5SYWrqb6UyUKSsezSrdN4acNCwObVNEMtUEQVZ6NpH+obX+lzBJ6k
6DAdNDu4RkOj1j6pDat8wdECA/gGii43R+7ynEXugye12X6npyGnh5H4cCdnTidD
ZKqp6h7rwP3zDKUghc34X8pM1PYdG0q98RkpRj4wa/9c+kMuzacCm1hDvaSQUCT5
5y3CaRr5sfJkKXcMYduRJ6Ce49W6wJYIXELDJCGna5C94Od1yj+NGExC5FLoFfFb
EkmGChmMkzy2czIrbXcVreJRUzXahnKoNGVgDGmxNBFweAl0cEEqtjrovjwKAjRg
asYWCaBD5d41wYL21erHz0hCHPIJpbQ9fHuOo7dnS1vh08bFxiqM8+aHwX7LnhML
QgnODjzFlvMrDXAZVpttzkb0Mfv/oFCA3AOT+MOCFxrCiXPEqdaVM77zlTJ5FmdZ
zeaGJYSlvvHGEbIG71VKdnwqWcyFs1GvPeDmejN2HG9iDvJwutK32sVXaB85bkV6
i/VcLZ1hpBwaIYt79yrOp+Mi1PQgjCUyDsPZu4LTxjq8qBvowk8UFwmgBLyiDvAt
/HGpcfiraSpUi23FrGWKKV/p0/sua/Qnk4Gnv4t/PRFw/SrDaWRNIWTOL2COOTm2
psxU4ycqzrHbauLsRqWhQbfVGwq/m0J20rO1blwgkSnOhuMF2c1KeutOU+SYThyN
4fUoNt3w3NYAp+x4cY0o/XirY4h3LBkrH8IfHj5YWLWJhrjODnzMmGeBhULDFHE7
vtYibOjMMZ5BJqKw0cdrSanMBks3PhViDE7cTIUOqvljF79REjH/b9yJevwLCEWa
wX56wYRMV33eIi4euA1wqFGYazln5YpnWuk8RoN9v6+/rcyy6prAxvuHNJHNWcjm
MTt/thWsUHHDhbUAEvkY1HySkoYgVYJWVA2OLPjkD4eeHSzaagxBjZTqQ0d76/L1
+U62nV9Cz+egVn0dqsEk2QK6WC+GzvRGhl+CilqdwTiIhH/3EfQ5+h5elWcntB57
2aOctOXaZ/5uhHZMdhBpR18RWBYNtH5EdCymxn6sznTn19EqAg/NHTZ5xA4RMBIa
PP/x+RI4IWtmXa92fJB3ujgC/BF3lOdHxn/zcOgOqLjHxPgn/N1xIHo4hpThmzL8
MG65n71fs3FaskV93g5QR1jYVO0UfVE8Wps600DyOmGioW7fPURVrhjYH9LVoXR3
qWAgsTMax9nbna3YaiO2sgvYA04C/nEfSeyYRsa4VhoCA3ayKiX67hDDEjKMOZW7
vS9ZcvsAadu+Qjq3+2UumhqPcWCj8M9NyUZVHM94AeRDVwgqDKKLE4zWO16Aq1s0
t0XpcekQHi6L45a88JfalYgiTjfxXwiatNidOhEjCL/UGBYgP2l2ru6IyQON89N0
3phdxPfrdTDCyhNbsA0aNBPzIPAOKs6GO+foH667POyu3phn1iBy0285YFqQFP9c
lU06VrPN69DxExMq0d9tslqbXasNnZ421gYxw40JIXIgvTMGA6vupp/u+TEe3MAq
EB7Y4/aS8KefJgE6V4zW1WSgucH90+OFLdYBDzw2RQccxzahDclmstUEg8axllyF
pKqn5Z1fStVPYEPtqt4WT5QHOcdlWPaBIlNWJtj4dygeR3P947r3jWUVfHcbmEYI
T36dhY3Y5QHtV7fLc6nzaGzeH58o9FN29bAwe6wA7r1BT9/uYZVa5QnlOtq7z3/k
ndPXrff9KS1ZEQvUsBXJbcDz2cTrhGkVNdLccOextxq1pikgplWQXX7CrpZiuJaf
v+LbEbsQ3YzjDeKjUTBxvQLiCGsbqk2mlghWh0O0cQgAHQXKxXJkRZOo9LUGCCNx
HuL1aYQxAq8nAfM7Vlj3jSWpEbxoBHJW91oterLG/KcR5CWQFStkmMlsC8I9rJIW
BmAnkq+pti4tpRVsNuWRO7Xkd5LAhhhID1LV/VIvGSPU+A9bMShftcv5GGhkKnin
pgcOWfINCUG5TCOb8U29n66r7zMXevTRcWp64jMTfTydd5+gO4Yg5SBgb0xqsO66
SnkYZxd/Ha1EZNwk71c0NXRmN+wIHp1EAyUs43fQjeDRtEFRSLgQGTe+4qBH+dz4
i9ke6QBH3JK7I1mPkEj9icZdcj1CXUavfi/81jJS6bWiFfBVFcDzqQTFlkJQ+XWA
bT0en5hx5Yf9zyheRNlvdoA7fUJz5joN2jCYnRTriwpBCch/JXYUxKWz1m6f/eCr
z8p1Og+T5FbbD0BcdeoOmf+YSvEL9aownt9Df4vn99wL9DVdXLpnIhdgrUP9Fkv7
aSsNDuo/G+aK6Rd5PSV0Xc/d7gQCpaJJxrdQS/EyanD8xdTrLbUgErui1qWNaXRz
MIchwWhDVB5x1NY4+TUQpf3vDvIMuP8Vbqw3OGqEiwIxyR+X+50I/Ve+FQWqslkG
M+6yaEAO1rkMNpzenvL9d72wO7c0/G08I3ooIWtJYD0WjQV0nNHmkWQBotHuUbJu
FKLmN7OaXjkdsUHgqJhiVZyt63o4uMDZTyomErxzLQkaXiPfGrsLU0f2GobL9ms7
4+HtnSJFIP/SMCw7GbODSgha/0hIr2jNmlPQKiwd+zlVaxxCzYLAm+bzwt4VOT6V
YWHv8IGPmS4uidzTHDl6HZa0fWvXigP9nBVCjlt5Hz7+Ccy+S6lzxZjm5z0nnFtw
hE77BzcTRE/403r1oGikMai4MSbLkWFYst87DR+LedWwmcDFW3e5gbWZS7Y6WbSg
hqA8JbMC9cO0nMgCkeJajkc32LmFiY8R/Fs3CA2/cXHjIXA05mySx3q/QhUgYGhg
+KA9TJl64/813qnhvr2MW/2jXfWcvk4GZRZn5eGActKc/o1pMPA/QXM/uDfMtvHo
5x/Rjpkw6nAjluBG+DhjPlnM9E5TxxeL9HghFW7qV76ScaCMEPiJGB4Cd9V29UZ0
p1PrKykwBHer/9lXoz3joUJwPlBGZjAwvavM6/sbrOJOYcedi/C9vKQQapQxbkvQ
YARMdKM7dXUxtMayX0JlLNm+pJ+yYIhmMwx1xqep7d5D/MC2SUPbMA+xX8eMJsJy
MmFmGA+x0EU/G4ci9WCNmBNA8V2ziNvwtaaw+H6ocW97VRqB4UoYjyz4COUq4TaK
RuZ/hiDSGkY38hY6cbEBnze+RtMjWhkzZaFtIWWy0mmX6+xc9/46PCon1MiwuujZ
bA45owelOhwiecMp80pbG1o2BqbK4qPxefIvp4qY+MPgXynMqouRmlxycAGb8ZnD
oBxwezKW1H8Y/xhoKBt0T4pPFd5ubqa4xoVjSaLEGwdqW9Kt9pbRYCvUycA+1QIc
D5XFlMK5gEQTK+7vq2ezk3fln04FGLH32xRpcYXkRK0grzJZPsVxODPFDJNcpKOJ
/QY5lx5w544wgi67EPwhbSwq6yLnGzlenvtHT4ia5Ex0dTDtp5TCjASZ7RJLgAwj
8rS6xRubuGVujyhdqvetACwzR4xy1UNtf9xWwYg89zoN+SNk4yO4NF7zhiDToSLM
uPezo8lXrO2CmD0mCkpvqHZOmmtboo0JjSacsk4rYAZNTBSdwoRG8wA/f5z6DS3W
HGqjzuBY/bKLtlrZyU68LYrDO0ANU+AT+evsKQmgnM+XXkddKBZHFFwCOrhl26DQ
/pa12XwfXuG56+9KExRn8Yd85Ygro8+E2ajur2aloTe4QTREolMpYNj3EsPcy083
OZpBiRtUui09Fs96TEkDNXlZWEuS43LAkq/uiYMj6gRI5BeYoWq6kkR0pfKoDXdx
cG01lt5JZdjNiwAsuWV5+GQP7PEgqwg7x7fctrNqWPlRc/sLwyAZYm0kiKcdPIjy
VZal5V/7wzM4kHHlKWQvU7sgO5CdzVhO9VGm9MEmn2vSD13lQNvditECgYsZUhhs
yEnaLv0SLNC3czn05XEonOrGHEIcvkWEIMixZ8hQnXS79NisHRN6tw9ERKciZK3e
p0XY088BWGsGYAUiLw1axiwsaeZVeAKV6ejqTYMTNONvOESdwyiHVzGXlJds/heo
Ju+UCSpH1IFydS/Dytgn8qWqItCdOGlkRLmvXoum/nGBjLOdbs0RMwMMLAe0ElEs
9i5DT00/Lq6KQ/jqHwtQNNq258J02RJX5Rx77fK+M9N2EFwtxLy9LDxX9Sy9LvJT
f5FrDYHYbTpjn8vnM7gF4ZjkTb94Y9jJ1mCo8k2I4RdtfCNy6u1N3uptA6Nwo0qf
Fovya54fV7hJGRaEUbLikSaivLd1aF+Gj5kAKK6WMVWSXTo2SOvj/bPLYupydajm
l7OvtyMJ/y5AhHCnQ+tbLsDdOj4HXgjBi25Mt2U2JfIId73vj8VgcunSg3mrsg8v
JVYEe8+qUoL0E+mPt1k6QXvC/w2072DaQh0GQdylvR/tASoMsoZT771Mz5kTJeVp
lkjX5UFTwOtXD+y9PfKb4UMHLxOEVC9/S9lYkFi2zXGZaQIuUCzgqYkJ3xcPjZYL
1IDCn+O2dgMvtJozQ1no72U/fvBXRY2l/7SnTV10bxOnEHHgt9UOxr8C3ZHvf07l
k8YGzem9gqazW/pPuxKq3ZEzlmQ0Litj9iv40kJvwxu1sG/eK6nYQ4gegzgSeziH
kaxFmWr1GXlfYWPU/J89PIz2LNoNmILf6HJN+Yube9na6fwXur7oXkAixLGanaSw
3db/+ZV+K2jPa/bd3LK2vObxogAcLxCQEoyiVA4PQhLsFGN7EE1IfxmT0G7DrBJc
phsLF94SbcyB556FZuUpA9WwdeF03NonGfbjHsGBbq2vs7cPv+DKCfc5tAqEfJU0
3sVPxn6vF6JJLir7vGZ5WqT5WfeTS5NQggWFmPOPgtp+Af45tQdquX6cJM+Wfbbn
/4y/BYK8l3GN6y6TJ09LOWAsg6kyhS296iCDXg0/78x1n37/50LWIOl6LrvgRAfI
Jhr4cLrA10Q0FNXxLN0YzBzFoiDmtF89Ja+UReDzkjOOgGvRcNgVq2EnPKYMqbMr
UXF/RhKVGXBvlPQJ5/diA+QP/+UoP3a8SS/OT8l76lDuvhIadaRiwa1mpCOeLjTD
RBaMBoZbIrrQPmHpi+h+Z+Dyd0N4Rfp9BLidajgK4pZiZjhih2gE9lTkSM9t7+RX
P9zktk28E/uRG5xatVRMqG2usbxJ1G4ocCUqGwuXRi9F9AsWk4cZP6f9LWnVPNXf
DsKK6jp1PQtndkfw0oTg8VdIA2tkoxg4WHDCKoMIgkY1g0AR5KBTHh53ho4EakW/
USlFWL9/85USyvHg9PdgFfeoyYQhFg4oMfwjBCrMNQTfDff+6oHcCuq5NOQqrryp
UCHdas8Q2x8Rz6vl2gcvM+GKGsE2Ysxla08obF6zu9ZDpxNa7+/Qaqpy+saCdYx8
jfI/AWvKc9vNPiyT94zdHHSnIBrlAvsAfDYJH/eEh6gVJ3+IbhxeaG8Vg848qEZE
LmAzSUZRT8w7vcshLQ0YcdGTNSTBNfMMKY7wRb4uBRA3+p8CCSAKyamCRn177O+0
6fT++eksqf1IhagDzFWVC0rGalWfo0vsP5eZB+tc7X31cuvUAYHAdfALNbJcqQc6
izB4YJOJtmdF7fbknX7IvKj5tVXN9tmNOpbJrv63WVtazCEiCWhUoreyauhhwc+y
6UmAErV23tCr5bjY1BxSQ8QBOXoQTmKz3tYF/yc1WbICwASaKDWy3Emq8Z8xH1cC
EdcrgcP5mBV4rm5Mgs7mO6N2Qze1PuLDTOquXW0G6rqDyldyeI9+Ngr8/653pG9z
Mx/x67/CKRCss+Xlq8CY2EngzA/lahRte+63cKPAsMymB2x13kFqUyc6UhCrOKE+
omHS69VZJ5ZZ58/cSWKItSyZHtUm3Kh+j8f+bGUxl2PCxzUdFTzQNrGDSLuxIwuQ
FRZkAP/x6TxDZxYNeNWz8XjpgEhrSniP3wLUH48l3JZTRVai3omI73+U30p+lYnV
l33ZKifg7c3C/WcN1bJWxB+0G0ALm7scLPdDJ78aBRAQ3eqnVLxycn+Y9F6M3gFo
FJ0O10eNcoaR5Bo9e8mOciVFGNqC7kTxIMOEZSPt+sGtjBFKI7f6Y9Novd40rqPw
HRgpqtlZ1N5rOu30/kWMh/9Zaq+be0S1He9XrKqMCIFh+K1JiXUoPFZsyIYQPsoO
2jADN19iHJ+xGjPoxC/Kss64YH1mZDcRQ7hwuWeLY1kMmHGL6Wt/ViC82OAoAMr5
wE04MtZ3U5bWeBKOhgoU5vEGGZl1L8D4ooyGK9WumWW00W2IC/5Hsi2KlEOVj+/s
O2f+6CTH2ayhQL0pRmsSDX4WNzIAXS5tg+0T80kBCpfGglJefYRxLdhW6bDgEm7b
7qxlYaHkeOnRHBm7dW3rlrtCdoKTUWQTO3BIy6n8TT8KxOZ/9jYEM638MgfI83vw
+e9AQyWlouvHJEqmbs6Oww3gB2F6i4lLd8BvwtAa1fviIKzqOGN4b9vGCezyVbux
IS57LYhc+W1ngmArE0s4jm1d0qwg5Am84DGye7MKePs9PITUa7ocNbsl51NB19d5
1qFu6dBxxeaPAoRa8BPiYsYtCp7c1mgcAQjimThxIkON06U9E5O/YjXkiYD2Dwcn
K+F/masTBa4BPpuyzPfxoUjeq/fvZm5quCCwR5BFvuB76DBufVzO1GAC8G0wq3yq
eQgRwGDjewRyEOziPNQe/lktxKQFoqXqpsCIdU5CXlrjGADUUDWtvxDE71O1Ws+U
0rZc0QN2O3grkrIgu3yVPzEEzlMnVGtJ9Vglwk6Msl7rtfl/3IOZTtDcC8ldCK+c
GoTtqvZWldT3zfeu44oH6SpemGd3D5pa5WdTNQtmzeWzG+3fzlBavSkJJrUJxRrq
w7zGNJnK2vC3u24s5Oh7TnXk1Za7wwDWxPl8ARd1JtxgHpPeXjMxN2Ge61O9LIed
7DkF/lTnEzjgPd3itFc/I96eQWXbGdFkeRehDt+KcmFAizxSLpah9VgC7qoD6XS0
6elEkQt+ubI/KRjIbnzTZXzOOg0RsxbC/N5oglYWslDxYsedE0hlCs3fHBl5Qmj6
+qyO0vZ4EC24LkdCq0yeyg1EDY7UK5u0rjTI3ffj+2ZI3IKx4qSgi0jiwarI4bdP
zU7InSHcg1Dq0lKr7qbYsJutdGZtu3FRHXh3mWz9bweGaylKVt7exJxfVy9e2dur
763mP+PyTVnjZeKMH7p5IQ505zSIGiJSZkfyNdNZKkceKjkOg6Igp5/KQC1GHKnX
LInHsRpA/+7Nk83F0Kosl0t4eFhTM0AAW6EizSk1BoHodMGMNULGh6E76rny1xR9
eil4OGM/xSm4t9WFY9rL8MXFfcLfsZuPcTN3GIprAgk68akutoSFabjhAKGGjC1O
hs7nHaVaHa1fvMhWmAxL7sig2UlhRxNE/w2rT3VZHOliDx8xSBjtALReTtdphG3Y
8hnboBAClE9NfhALgl3dS0OtvJ33ROkZCrJk2gXvyka2g3/uvqcH5B5s1I0ZXSNO
olsl5GR7Q2Kkek/vSZaiQk8GxQMBqt+WPsiW7iCvPPwglCgU06JpnCJNBnHqlIAr
i40ZXIo0YaCNX9KyzMHRzClWydEQU4tZkLtw+bY9ooO32d/hDQ8+e+m6mM+eOLpO
45/aO26UXK5CYwXvJcCJknjlC46o4w7PsmL2YAeyqotZWECHYNsN6Y1NmrmNvxSH
IBjHdPGDs76TRX636pe6u8HnxiKkhrApcahCxG/Nx3h69TJECJBphRTC8/8ou1P1
ZZ6PwNPfLKro09lwn1wPfHNYiJ1F89o9yyvLLupX6VrAo4nn+H4a8bHYwN1nJd+V
Hm5cjCri6dL4jBkWvmARyYRXmuJAlnBf+UEE2R0BQFZKCzjvvyJp2UYOXLtWiUzz
XshSVSKu/feu2dC+zDbuPvZHX3x7RurNYn63nm+EZ4ihE+24yKVSVdowTpHm2iqN
Svo9mmdZTBVCrdnt6XwwcBpQtD7gO3UQGIBpM6dswN3zZmoPFp2RioYTBzYWtxlX
rJ18sAqxUedBDJ1J/JPr51mU3MNrpQboeTx3iapSeTrNvZOzeTHhXqfUTOJMixZA
cY6Lo8dQ9bDJwrSP8Td6N0NTosPRlhKnWoE/syinOfJoJQ71C+CsgopKeIm+nSX5
kJcc5we5KKLzRF3XtG+PBpbeesFvFTIDj6L23LEY1X+6DeUBaeZeXog1OPtT11RW
uxPkr8JATH7ahZDxSoHctoJCGqkgkrXWLtqeXpsb99Z/nuhXuhobmIL/R6BeNtOo
pEcZ4Rrwi/8RPppmEpWJtbW5l2bLxJ6kNczmZdozXw/3XzomWjf/6ecOOAle36HP
B0LbZmiGUM+oB/VfMdNPi2px1gEs2Z5vMvw4lOxhAdGza0LrV2GiEQuBaV7AxgYi
y2pQ7WcIL5ZKbFB3slfhsurEQTLSK6BKp3qlacEN2ZldgjjmIi2RZ7O8j1vp702l
yt+nDEVT8GbfDmJhUzf9orgFOqNOMTJXWXrAv2+BxHc60Q6ZYYL97/hez3uap4nX
8cWSmGpP1+b+vSV90tl/hU5OX8kDihjmpnC8SGwZVqNdYcp96fyJnEMD95uiNmUe
LejECaDtj7k65CHk9RsEPMyk9KCuhYaTLoUpkpSDFhYtdHtWAWsjrAw2E2cTHDAK
1+XnKwkRqmTUy9TjqQJ9IYXTMMc9wGmmAF8jCFwhtTwI7uFJj4PPmA5EoQ+UygjL
2Tdws+srQMVxHsjvx9UzHiI+pg0fCbTECMSGITYaZihnIHqf+W67QzmK5WOhvjop
LcZsJcVj/XvdeLNXcyA7PgojXkdUfVm/90OvOl5AaofKT59XZ7P6rybAFPbnHqsD
UNZWESTckTHzr3x+Fh4MQ1Zv8Ij6oAm+9Mubkg2XCo7oIUrmVoYt/SYjh4wkPf7X
9jZ6peo9vtt4/fMZvf/utYLvR1x/ggE9vzulLUKKJIKNOpuJVw35GxgEPMe2k8Tu
n9DOhiwlHOS/1BSBNP2DLOStL6MZTUctlHh5aoHKnAZ0TzE6+vMDwfGLzWwi9idp
NBjH6U+37JYNRw87nyYehVfMp7MGx61SvARLvAjl8/mUBclVIjv/pXXzevyqL8i0
36WhXtxB21aeynQJvxwvkXG0i0r9D9vlWvDm9g7CNaKkxkGK557N+no0pudTRAIh
17pF7YpIW2qVWM7Gk1yPylcgDLyKKGrWyv6DUKyRRAt2mNcLtWX/MY8r5RRg83DC
L/Nf+haAIubAqcxzUQu5nyiw6facRpqfMAjReQyy3396BDp4tNT6vXxCplvUXX1e
fpKbGwe/woLH8hqadQDnQgvmpwDuC905i/6+kmHpPrUuMbm+hQxRP0R7Lr/cJkx9
WZ2hbaublLFQIytJMwb8s86EF6C7e+Y0PNGxwKdyI0xJ8FESW2Nl4tI2mmvjDFus
dzY3HfwkkzzeZBF68jcKJR54U8hhkXBOcsD7eqqMwfbY3DDd1Gk6UPhnlePmaLcA
y5aXvUDEXZ2+RFC8QgtRKNrHgB7Vcwh4QeIOFf4Z3ADtj46IvUPt5A4EZWpJUHQ8
o72dSb7UABtctkEq01WU0iQC2R5UbfphpiQdbLkl9EqlIwQa6+LRmjUNKsEnyrxD
5OKHxJjbYewqJcIfSmN02WtgRKv/jHrJ0rY0akKe8/oFVFGdBnGaBD+Hbkgw0mVh
ernR7Q5fqAY1eqWISEu3VlerloHCmyoMCM20dQqw3g4VkKX5TpKIMrYVZEsgoFtv
ATFYbY2WujPb3sWxw6EGEN7/pCSQ38VS0UWIsU07wSSB1fjFBqb3WSCO+yZFGzlf
jn36wSI3YKAnzHsYW4mOPEQv7vy8IwqgBUpIrDAHVuja9GHQgQkaOwxkkO2K9o7j
xPDw9fTUtFV1aDQSkf/lY7gfaxkqsXh7ATdV7AvqzBxqdUe6RCJtLDvJFAe6qpBk
oQJ2Z0QsAXXCpMD/R+ekNfIh5cFhVtyQ6/dwciWzMxAHVr3dyZqXK5/XbKU39QRA
lmDdwPUCQxbVTNtSBCWcAuaRaXYakfdkN+LdVAfzGOaDzxE75vwG8nwJqi8Oep8U
wYwN1kgpelvNkOUKFrebE8s31Pb+3TkldC5NQcLkX9Y+BtlmSAOzYAMHL50CBRLh
i02HSMC3Fxs9J1YgXiyv6oD+eirIQB19HfLaf3zviUSsHTUqTS1u8/5DBgY7RgM9
osn7hSyzxS0Yrxrngf4fJgZHgs5fgzpC0SQW06gaPdg02z870vADnp4iRkNXfXif
fjpTGL8bhNheI0LJm8+Q7oQorCgTViaBBykgUs+rzLnpUi5XTTAiykQl+7+eiIKX
`pragma protect end_protected
