// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:36 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hoWcYbQAQFqd7Zd3h2KDiatocbZJcbp2D9ufqY7gKhzb68r5BFnH9SzC/kHRF3xr
NbUp0sFekouOeX1muAmThaEoaa+RbGYQcK/ZFO6QsK8hh16bMsR3U/ouksFY2bZ+
yJLf4hdt7h+qxjtDtagozWHd500uTDuInSYpsfm+D6o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17280)
gXa5ubPTpR4DqVm48XdA/36ZtGSP70qi+DZSCoo6JXRwkzszBrjvd4WGZhhcOQSK
wElo07l8qUf7JXwBbxetKT9hp2yIpl7S0r8FtRpjtf5uvjhkeE9ZUCsVmCoitkzL
ERD9f1Qpefv4SyPFUuizaHP5OmSBK/Fw8SShX056zucscN6dz4I2iKvg2/jrZ72+
GR1Mt6+0/E+ZkV+7rbx8vjb63tSebwkjik5gfIR5oJFU5syY5HYC8BDI4qEdeqre
GaXlNp3Asw91a+8NFTUDJIm4lNNokUUdG1jpZ+vqCS2QmIsBm7EPbwLaot/2zFoe
1vkJIwtqc20XRLwqDTaqe5m3B8h6f+A2Edmo4QVukB4xHSYGof29tU8P+9nxGqia
wWr9x9XlMjsmrXCwZdKzVVDGPFqD4zoOo65D53c+gPaQwzCDS3OgL8ehUWMKb4lL
d3o8EgHGKZf2CIwdDbHAuo9/vKHbePPdPNkMx0pxH5vSE2UwYS8x2Ho6QCwESAS2
qK9zd3OMbqXkOPduuJ02svq0epcbBFVffi/JrvH86HPk/Qwc7DQWB4EPNf2ON5fb
ieA43qQDQYhb6qudQGhYAatnE0ALun1HznZ10xfIb5urOWVhxZkzl96DbJ2kIsdQ
bQMUbEOyZkRYqihRirL8m91HX8sYdK/fGOr9/mVn/RBIm5yi1QDN/T/oT4mNlV11
VBlsVP7sQN3kFJKXbnRWYrEMGoby5m3qztxK4iHh0+Im+712eGOK3Ju9ajqbGfr1
ERSr9GspFkHIfn2/gm+Ch09cuWF8JRGMfig7M1aEEqsjyOLjDaPbKjyPXY4ZPKQG
VknCCbIWpMseLr3ckOj4fUl1dHrCFgK6qXeHupblbNeGhRhHbPjF7YMBibEm8Vei
vEspaFjK5H3Sse0jGEAW7mfEsRvNJuosoQsPaOaQcKKJPFirjsl9tlW3kWJTy5xW
2oCpSGoZQRbCKXTnJrtFwIeuLaj62RYptM4sxsOyJYFXLQ64cGH9fEIlI+8I9CHd
4obMFIb26TRQFh/AFZwWUaCVPz8rAjnDmbCvkwDID95T3Icg44nYGDt0jKB6uzqF
NAVDGDYBFzG1aCu2/lgFehJL8cyg8OH25gM9nBcOIQK+UKQFHpK0OFAMD1EMRFqo
GgpXu28H/RxF4PURSP0VbCdnW7yLmajxsCS7st67W1WqVJANGrniBwG62uQpkAuW
YuyphnuUCCECGbha98RoSJhgfXlEanEXUPnkFg3JVqbwgoDjW8OnLB+E2lqxoWjq
FsEcUr4noxhd6tdPC5CoGEiHyZNztMecydgVwWlLt6gmbcc4RpE8pxuBYfKRRMye
Tqzul5CxOaJQpRz2CVRCRACFh88P8+QLbq8IaaLhVnUTx3W1mojoCan+hwhu5UEA
W9U2aYGsscElEfPQngLanH92lW//JpglbEE1ByFFMhTJOg9HHOT90uAEHZHtmUKO
u05QeZAlxVlZR2WZhim9LC10FjrlkR1bbOubw33xz63sjsFTNQz8mTjYdKKr49lT
8nZgh49eoAdJ61BF+akDA7jzvbeAVu7juLBz7TUkMTUxNNfXCAh6XR4b6RgfT1o7
ZgPZgyXeXni9K1IXXH8e4dJKQ6owR5tLP4sQaSF5fqmagDL4E7dP1vC+WMqGljlW
yBGR3pXNQ5HGT1fPlr+MvTPPpOJ9InXcJQOfwKn8rumuZVvknR3jKy7QpWNiK86Y
PTL3de2zA2plQ/3NavvuVQvM3ArGbGFhvSMAk1JYFmN33XmSHH0rhfJ+SQYmvCKJ
wEROFT07km779npadivS0q1cs/75LnEecYNdbSakueopOmMD5xTbP7A1PyABlG7G
huDubeq+8VL1jONuksXSV3O6tpNabr7qmf/RVvaDPb3csTa41nAMeIGslrmsKEhd
jJAhb+uGHzK1QP7o60wsxNgEcQuqnQWNJITH8AWLwo2E0o8H7tp5Dr75d4YRGGlV
JPqsFx97pOya6CRu9PwcZjewp39lAQZX6YHAqlnwasaO0KO/YRe2/mf7ylA87CjX
YySrL3LKKESGGSBjdxOm9ZCe6WzmrFbWpNxTzASOcmveK5Bv+i6QCMUzPYqBJ96n
MHqPK0o8qU4TyI7Q0cTdNe0A0M5BLqP1veBKfnbmaLGNN66LANf8CcPYevonTMaS
XhRm+AZ6jWYb0peCbckLn3WosHNVhiZayDt+6YShoznB/gatKbmkiKii+kqlA0bm
CaUUsqzhkgIPVxiTsLuYtY2ZqdWJ5w/lVpL7CaCans9goyRZ7qc6x+L6nRutFuF4
VpaRTXhgVsgbk8POZ5BWhuI8SeUwo36nwC8LWzrNJPtbr2RqW30YIP0YX3Y7hOLf
204zldGtqtFXFvqtX/ZJ+7EVkREXEVjQUlfRosD+oVtb+Fp4O3HBKBWpo88w7qzF
6WgIR6Toi0Up8zPATc92n2f+A79Nml9V7IYpzFWm2d6pUjV52pO++vKg3UgtkL+5
Q1vZKiOe1bf3/fHbXdspAITK/25ZAtGbOp334W9r7nuEnfQz1F8VWeAU+xLAHNni
cL7NgidbnZ1NsSuDZTuj04YL6F2Sbm2rE9mkvtSKwauJEn5aAEY3qUw7KdWjZ6nK
O22nhEw0dUNWap5Q01F+emLc35A0pQTPevWV5pgi4IMhwmiyoe4V1p7wP3dl1EJx
xE1aHoXx3jOlrpOrz2SjPowk6cWJ8cYiTYW8H9UGFLdygogYMpz67pRcNFYAPNXq
mZitemR2pEBb0lXmGLp/L5ambvcHqMEr3QYR7UGkVE07Dk1LR2spIHOKv0j4h/zw
Edpt8ERVvoLo/XGIOtY2mNb71TgVEW74dTleWDU28aXgPGSYKbDIiKy1gOqnDZYJ
d07kEr4lCGFR+fc8/7VCAijCAtCsRlNaaE/5JoLysFoFxDKc6iRfrQhy7PPwBaYZ
xKDkm+C8BbQsoenS835mQp0R1Yi7Xvh6+zgj4y9tMZnj+jXahC7QDYyCAl1IjViT
prIK00grCFAFexCnCqxp0RdgTJgzk9QipODG7VBU30mf3/wuQ+HYBrfPBtYmEjBz
zLTAH5bz4t/C9kS/0XuRgaTCAq7Y4TIdEROShCJzwkDO2kZY9htfGoGpnJId+zvg
2Zuh8794VKi1dg4miEQ50VUECstgV2YYm2ljIFQCKGO/b31BynBo3Kl6khasBogB
lr22NLGCpm6oce0lr83NlY1Z+fYCodeUP+eX8b8P/qJT+FNXBH+CWuFT7JILEiVb
gVfkFGtI7CaR+bhyPPc7hv89TZYcIk2aW9gVSDHcxc5kN751LzTebvieyDw99weR
sqQPeHA3zn+jK1/U1wK8NBuBITigMGIrsdRaAzww6esSp2LwrXycR6x4Df7lqGb0
p6fWy/qxVKQ2O5phqGeo3FgMFrpPXwXCfeUl9nqbqwPu8/Q+q4Ba77Cf0XbOGjk7
73yM5WXfP5GfnNVJoLC/tMw5w+h7ASvM/+d9edKHEHjnwvH45FFMuAm5AAAcnSsR
R26SSqQWHNQ+nNvhZD8oRy4l33FaAzNfzHI6u4d08rvYS37yCgf9dNydhMLwuJoY
Ev+00saftiDlm2t4oD/CyiA9nrQ6pc5E1s0jlfm09cjDbc7kBz+ULY7xBtKp9XYY
FxKRhoNqL9LC4RZLDu5KAKXcU1PMo2Po1owL4IdyLJXMkMSIKNiYDm+I680AB/hM
AYdcHEQaMLv/ACgw+FfI5/N2syPadMw6oM3DaCRSv8i6Ab7p6bqRWkaazp13stbc
a/TTpoIQZfQyH6Ginxsb7fk5ducjoBu9xkDmL55O7IHx7Aakgoi29PrvDlDYB99e
cgtyk37bACKPm8lwqQhlhHpodrR8+tJQho9ZuiUxOl5CNvc/1CBCOxGSlk8Mf6oo
KbrzQFuTqFa9YedV0VQjzwGuKclDLpFTUXdLTxUYukbc90FPgiOKoYG/5AM2dDL3
xfyKn2S5dP5EQpjzfJj0SZ8d87tRF8wDtVKCovQseKH4edW4945a4Ngy9JjGMiYj
SGFvSSG4i60ZsJrkmNVf2vVxxg7gcVaPyZOTVyI7b2D9LvtONXUewxyb35qTdS+A
zl610Ekk9MkerBMW9I8lnteqDzhKIBNnnrBPZGDvaDnArDGnPOYEy5kLyiHd6Wql
f603Mp93unAoP5gKQgOcdWQWsDLJt047DAcTZ/SerJe5Xmj1H95iBS+PhKLrBdJZ
tDTIYcEtFrwrhwg1Xymul5hCykCqihx4wIVVy5DPpQ5g0W+aFtsFMY6ihIOddQXC
RJSOdtODTZJ3KGpbix/jQrolxWYuZkR/NzJez7Oq993YEA8HIcMAwkcfUrpLumUW
sz0syWDlnmSnFy0e5Vj1BsJhntuiAfy8O6HGCQxhJWVl0xd+U+2mjUML9FilRdvz
f2MmJSdX+gF1nIkQ2lqz8/Rpq0Kw9HvrT9zc4O3IyXdot/+2dKpNrv5WtKZQr7iw
4XqTpkmQ1JCw3AkEVEvifs1tu1doPC2vYlsH664ckuQHnifjByzVwVF6axKEEe32
uZNQYb1N7ZyKw3xri3e8dSSUieG0aY9P3TDf83Y7oTQSbK3lXhCq9fhgChJAPZNI
6KCXektXyiqPQdRYqIMnU6AuEnRYT83ev7w+lUePQpwF7MsF1boiyXCMevWkrl/H
Cb7DTTDfb7QztfNC/PVA5t6w8SQ7/A4Z0Cccib15OsPWxlTQYxguOdIlfmhRfpcT
aWXmBtAvB2mfutMVJOKcLsah0tBJox0oIsPrdnu680A/tMQGv2Trz8C98olNMqEp
1Tf2Gx6vcVJvJuM3g/BYM6PdO3pQmuCDRNxo2EG5E2eT24terHfLtOWpx8MeEgF7
+KIdbNsDwB3fxE+7gLZ83UhkqIkF4gn5EDi82e6h2fv3qnDQJHBfwOzZ9SxuKF/P
vy1AnEsH8EY+oZaME4DVnWrFoaRfCCM5WVJ52Vb8dTlYvoyTwiQA6RGBOhTTAoYT
DmsVNlJzHg3Sw5PJ8D6FCDVor8h8sReyEh/Z80j6ke77sQNv043+ytaRVG53rDpp
a+mKIQeK7IEK/yIvoA5C1wf6i1OrAuajUpJRBFhdN3Ob9P4PxHq8PkMPwzCYsXbS
h/kjLpqQbJdpfysb/8wa7xvHKFpN/sbRpn/rk8AnIIFLjKjN1nBNxkSTYy1P15DR
RqD0JnMUYtf+/jQn8gALLnjNSiZDZGLIkGgME87dfshCgPWFDWqn6WZum7PW0zMi
iDCObIRpvJ9gTkp8Jt8Z+7L1NsL0q9Np0NOwO/4Xg62rLZEVcrjdO8MgGHgAbwKP
b7OwJG3xS/fclaseiIfxAmZe8GHQ5/VjZ+cVZh+JnfAK+/L9o4VjZIkU7jfsHJFV
PhYu9Y1yS987uUcdj1U5+nWDtnhXPqH3wLMtZ9EtboTDFqHNAxXLLW7lI7x1soYM
Hwr6v65ykO9dq/lRScdxh+RI8KWCR1rKpHHr+sfgs0GasEDnrXejCgrUINTU2G4y
/7XdkPTinvR5PrTbFQcUy7FaXd6RMGra0dnX5QrSMeHSCZAgLx4tWlHRdxxDYmEX
3+DQckMsrWU2Xs7G/qcwdRopz35vnD+xkJyis5JmTjdS2OBZq60DmDHOgRaEEzOg
qKfSMrQaEl9xwX9ZY+EdceV862kvaqRNmhDN6nwU+9I/IKpF8tuRksTX47vWP1C/
Jf2rem2oPn9gp0crqtbZyymVbR9Z/k3WtTTrcX+MYir0BRF9Gr6LFpk1QeKfOtP5
uRzYf144UpGS1hV4kx/A/Ilm44vZ3hBWbQHquDO0OA7YZbnSuR4HkVIyeemtL41R
EiUAndyJ5q7MP7iSniBQKBxLXOfEqUc88K/xdUeujsxME9mdU7sgkIJdDYea10ss
ososB4f3XidnoDciWL5s5dp3jY3oyakzDDx+vRoT9x0cY647yChcxf6tgzEB9T8Q
ExdL7F3SR9ol3t1fMy4n0yok9zh2XCMpsaDxywgLnkcV1IiozSpTQPQH6bRgWof3
OeQ7Y+EB57J1bT6BYMMbHm6mlDHNJxqSCPNJddzPOFn5Q/wl/xVFokw3DZcN15Ll
G/YK4tGvwmToGNIlrDbq7/JImDIZOXUBWj6+Q8kQlDP3h384YdzGxLrjnFYYyf3M
9TzLVxZoCfsqjX5ScfTxTopDGVKHEdrXFXCeuTaiaYNKm0kyEhQoRy2sjsJutiAM
1WfySxbmq7awT1F4dqZuVV3BcGZLdxYFDNuXXauH3kwCJM5WpgY20VeMPp/kphSB
ZwA0LbcD9IjpzQAcZrXmDoN/iZlqWoS9r5Ew8WJhTmQfAipr/LkxhDOVM8ECx3wI
LDjSyD87vDwtSf/OYaT8hmfave1MptoyGUmYsQO4ZEsAAZh/WrGGWuOjCZlcz+8O
4LuETA2dqQLiWWezZoxXlGvUsZXUBxzFNRRakKZMNhFNo29wN3EQLyD8RkwBA4nx
AaCeFuYBs0DD3wwewirquN0XOJN8nxlp7sfdG3XaK6mhEvfMvwJRM8XkRJmBkxL2
UPgO0YlOnovMlLXrXXbRKp2Jch/gaWBDEBo+e+b6mgACPJxId2AVZ/u7S+NyjYQb
fPqu5piEYBSOx5FGmPpJUXoUM7jid4aI9G7ZCok0uE7uClY+899/nv+YIbwJUGiT
ALIjD533/LJPa7BnsN0qF4nL0zWX/m6LV1P7u8WngEU77bFk45/DdgTvM5R8QV+1
hOxFwYBiOb/JMR1AWy8cjcCGGXUj9uCfxejN1aVdQRFHWODKD8q01YEVAvYLCgxO
Ao4pzXllb2gOdaxch7pbfkdaiZ/bulsAWM/oKkr1qzUVRhW538H8RC5TQ2SW/r9G
ZXm437a4563we7ZTDhoORiMQaFCMFzuRRxYxAJgvy0EcswSJVg+57/l1mYQ9EPYg
5gQ6f1NiucYVMhQJe+OrxP6SKmCLDv9ZUD1H69ui9rbrs3PGTWMZ53cgDAejNFw9
6vOdVRiRK0ZdVFW1v+3sonQSIJXB5GZud0tr0o7P99qA7GAUaa8odRJXovRplVg/
/SNfOZNi0o7RazMaXqreBRVuWu2nGtR0tOfLV6FWuC22CTHQjhi7+K3fCwUzDsJS
I1txlQd4Zu41c5rrCoUpO8EYBTsfhm5enT7dnmFAxeokmIqIpdSzN5upQww4juFC
mFY8SIgxgPlTaWv+/ZGJ+pZ5o30N1+TS3QXAnTUlk4nN6yOa4M4ZMFEqtdh0X9tX
wf/8+kjZ8/+Ca8MxNc3kjGhLE85fLBWiemOd5miM8K7zroMcCsvsi++naIh0cImk
2ZXdQjpD3csw36crFjwSs7vLgbfrWWbDyRjVgcUfhBsgGN4ObMXN4Us9g8I0xuWn
uBInIrKvqShbEqZ5avLaLeSy2Glb62rZyPOH5gD9DYJV6OhBz9Vio1u22DfllpQp
Unz9vkBlmOBIc8bAtmv/uEHjdljurZUH91GQhzhlOKz+VgyLo3Xdlgnt9yHduP7p
C44BsONgrdqf/vxcLzTE5syGxxFETvcaI00B64rRT+rtxg38y8Exmc+kONApM6is
xUbq9AR/yg6z/e5zJPcY0xHsTU/ikxaVTLjU3qQEKNaGhFlM1Jhzafk+rTyxZmEj
Z6hpLb7bZ7rXgOPth9hG6ODnw/GRb04eyugzot1vXnusPXG0vKKAEV58FMpGZ5fk
ziDgEqiSm5cYSURmS/DkUk3+xGH23iiyF9Rasmv9Rmun6tiA5BHGSO1++ajB6V/a
3hgxP9Or83P1OKCtd7e4G5tKCDG0rL4AAxPhmyuDb5FTKmIdhLN6A17Kx+hdKOIg
Qq20suSoZRQ+XyrLRvaA3nQ9HA5rzgZxh9hYIxSjLQyjxN7ToWaetVEHqyx32b5w
vZ0mPeX4QRyRKQ/JG++Hj46KE/K+rvJM1avVM+0eaAyKo7FK6xPj2xyZZMpIDb5D
JY+HBIwtLPGLCi3c4PGBkBkWTqQvQ3vBcegj3ETK0I5YP9CdpdWkNf41ZPQuHf5h
4XAt8gsLJwWkysGGL+WnEI9aemuXVwjShRURVUt4s4TqTvlmHqIkNA0vqj10gR2S
DDLraXNgC1Szksgp6rQw6cVOSCD5b+6lrPM4Y4yMK6HLSXKOD9XrYERS2nDck2y2
r55IP35RvzkwW0v9M4DjVU+Kko4jGjOfi43eguAzN5sldMs3vfKH4GklVp6dmVLQ
PEpk27wso6nzspsaCLtBbUFcVQgavafxrN0oG08YiujiLqyqNdZwReG9DP7D7ppl
BHaDAwlyFolFCqp0ZOsj6YWzCF23MVpzhjJdKgw2VWKZEyH64uriSOKLYkOOWtZp
SQxC9vu/NHiQ89ZqqSvznNZTU+6p5z/xR+QqmKjQYm0xMx35Z07gl3e9HwZbRTbL
J7vKf1Is21HAewIiDVz9Kls9Gdw5VMo+8W6mXGPFXKe+aar0aC2z1oFMesjtpPOs
g5/MfyN7KVOZ5y2gEX3ezeNv/FcVl6MxpWDt1BTEQbC4PA9arsd0ewe0j+yTzJ4p
Snuv7lUBDykmRPxcoqfcquhuRjAb2XLmg7hthBXfKOVB+7h8jfXHw4lBfJiGW5+T
aMjiqGIar35EnxDEKLFU9uSev72k+i+aFrEShcjcgxOcT2NtcXKSZHQu2Jo+6c0r
9zVlUfULEKmXeILrHMVvfTfDkLuid1ifV3q2ApdSBAHdZCYLZQWcEW/aJX5BYpat
pR8/3oBjslVRcxjVOv9MA+LE67q+gS4E9EUq+dloTAT6QpQc4I6rVRpFM+HcBM2D
fanpsyMgQWYhhRnPNQlp1UkeR9av6YKKXKlz1pnlp8TZR4Dkzmo6paWlbawQ6Ltm
36+SJyhWcbi+IfE6w2ALJM7LOu+3skb2aAowAGck5Xz3tNo8df+v6IXPAmrugynE
ZmcNSz6usHjflh0t4lf8v4HwEWODbdo446X0af6HvPLWZinvkvSs/pcjTqcS4P6y
Mu7Bs22RKUM4dVp5/0nUw5POo38EDFeVJLLbEV3na3kRYHqKPxbkwsN3mZkn8CIp
Gv9eP8GJzLvLfhx9s+4fewoP3c4laCxAamcrvrDWSmonfUVDOd6BBiDXjGr1vSmf
2GQ9zZR98hNz7cWfhRdf5UCX29oDcFdVWERO1DYPORY77oP4XkCncevXnNBlLC7B
mMKNCkoTi44WE+xDT6DW2t1XzlncN29QhxJfJW2gvjOgrwTtSGjczyn5PEXQ9I/9
VGutR6m2DgjbeLlVUjlNUpjnFsbyVCrFKYVeM/olPvbsa96A5YBKhdUvUKbK1l6p
t01g5y1WpDwQlratL6OeLy1QoHGGrWnNzQVUakvDkxJEtUb6WogdUOFZoOcyFHaI
bJ8e+O2488je79lGifrMHZEPPKzH1aXf/G7lOez/YDFE36q6IRMAMxmipvovuXMJ
pxaSeWgmiGM8cZnZAWo2JSElREq2YTdoimIVLyp+0P2dOsv66Flr3WbiyH5oEyVr
UMtoE7r9n5Jo+Z8eNZuu0KaM9ffWZ+N09+l181EorYdsfT/kWy/LPst4liGSA1L8
sKZswS5OFpOe4NWrVwNDUbhrBfE3IZO6uvHkRk6dKlKJbeQM+iawsBFrnWeouzMH
LktYyjeaSSVLvLDM0ap+o7y0gl/nk3u7G1admspGwPn4N2xkmuQI8Lw/jP3tjovB
3APFd/ncfD5cgEgnMJXn3C5kb8jmkv9WI6hVcsxnMtmzEGAvBLb8UQf/ayrhKtdW
W2tTj2wwtbAANMQjpwfG6M3zHUmA4eJlOPOPI0KlV5lfLRw9IPhVF9ssdfPPdVXc
FCeGw7fC9ByOFVB7PBXFwLp183mG7ohGIktYw5UaL9ZMe5w+f0H8dpABx2zdTNxx
q6YTwSAJ5+/fKZpWIQp2hw9cYMqwG4ob9SUvu8gEo8kf2/F/9HMyETt0ZnjnNpWO
iulsfr9TZ7LdlWVMnbPRbbXm6qRtyup4PDMIn3fBiAa03f6yNRcfXMTAqEmNu7gf
dpVnBLJ/5RRJSjetzOk18rBWGaX7X5VNgTgSVBK3eRg+6GZ99vC+k7dc97WEXjPf
6ZAbuNqF3cdw+OyJgjPDnC18lA2/U0FFib38xpEp3qELxap8/3Ai2WmuqmyPfTJC
7hmm1vYrOoYfMswsXYK8eZIBAZnI8tIb+RVXGt1bLBHroRGaV8Pw2+RNG1o3nWzR
FCMDXWqKNhCe9Y1AsoewtzJaI4aS7b4oSOwqiOlfjd3O+YDTZNpiYFCIcywdEfQz
cD9j9Zovw9cc/m/Vm42Fgf4hAJrY6AitN70dMDcB/AwZfx7jOIzvMa6jvyKB/WAV
bA4bIzopX4k9gtAAp5n3bwsyKanmnmXNsWNMtl6PAdoxLqODuMMKksEFtMSBO8Ss
T57NIFGYt+7Q8qJXz1bGl+Cht6g6HhCm2jJXyT1cG/b4wQBI4xRjrlrSfPbTBy9F
FbcgpFSuVH/4KNJHhuwQ5oe/TPz7WRuYDEuKeMlFasy8j1+P+tlaahUco3MyKUNh
+93aJJyWUhMCLBe5LLLNc+lIdQ3wMGtdzcm+znyNY9xUDPiHGQDZeLxPSf+MWbXo
RVBAdSOsb8bl6OOMoaTrsq+5Am1SC79hi1EAi1s/7cWV+TmTl5cBz8nuL8lMsZ89
jkwU8wzTkxLOtqnR/fbTF69YIucgvmMImh0vk8Td/rTbOm9i+S5B1qD+eD0DnSyY
QLBShSyKcK7JMx1p04pi4j3/hXKhArags6Q1TzSjEV6ryUMui68luryOAIHBIwAd
bUJYSrJ9kxWA/wJdG198AIOhQ6WufymCqpapkmbfpS+/QHm1PhkQRjsfo3+mfI9c
dnCh/eKAzOQ33Wl3wcpEtL5/1wkQhclrzIr6KFXqmgVlOooF2paEtJAoTpVdxrRC
RdqLqZrVNG0f3cjUpkh6fsKfm5c0M4xkxvglfUDk2GrUeVUrRcpZ7xGu3y9dC3IX
AqK/oO4SsaQcN2UZKqvl/t+VPVFJ0cPzaNlR8w5VNN6PLtVQjoNY43jCwtvf2PTT
JOiFb9MKQryp5FSFE0kSTJlUvu5cJeft6DyD0BLDpXtUyQNfkAzFFUnu2KtxS/VO
nN8B/YEtPBXy28jSCxUw/S6zv1sZxUQaM9xSM/St9tQddyGI8bV6p5+TcggnCDK7
FzHAQbYUrZSXP9/uZUicdzlel2cAWoN4T6je+gT+2PuRmFaMjzzB5oLRPpBLLeuU
H6JZVHp9shnnHXZ4W2zCu6KHpFdi6u1KsDi1Y2Nd5gSZB2o1UqgN/GIvIgu0nRmQ
8MfJszBgnVNsUNG9wj0UpHA0UndzCskueA9lfGZrc0hVohCtrotCycxPkEemfLLE
8I4c1OyiCIDV/vE0GOPYL5J7R/3odrqqgBc1bitoyMBqYdfJjE8TAFndIctNCYal
rn7ql3g9Kg1/I03fpcg13paq4gF5r9h+LZzhELUCfQbVuU2DuQxkC8xrj7ay17P4
taPrF41REBpMNqoopQbFZo+E1TN/ZHhonJ0rVmHBPMiQqnWNls5qA6KhS3h51y3Q
XUUoLZXP9I0X4jXOYmnKylECjURRpEdOucfwvLdpp2zaKJxO6m16+JgUkjj//4Ie
WGz0Up+MG42QMu3aFxl2kWHv0jJXE8k/RWpMErJ4rZbkU2r17Es+mCemHB56xBds
MyUhdwaMEDTV8o1G/OHf1DxbU05E04gS2hwFp83aICdWeEiCn//ESOAqeZCNvt3z
9iRKUWB5HM/z277WSXMWtjw6aub+Wzje+TnHyc9h52ERvZJx6q03UieADZznn1rh
9p8lnDn/04lN8ZH1PvAI3OXYVVc+91tG+CBZgl5y3rJQGg9qMBxNDRT2brEr+ndE
gKR3aenvPrknclcde1H/CexVBDFchwlK7P9SXtTGrfP38fZ/BOKKar8XsP5Di1nl
XW3fXl8RLvFB1sYWsLE1OwFhAe6i4r7oB/HfoKJ6H6jKAf15SJizgVR35CcnS369
D8796qkvl1Ek9b8firItL0UyU9u9PvSeO/wjFriDXiDEUs5j2ZemmWL7tGQeJrgj
yP9C5AztgPJ6fiiUiSgs2MiWmLQIncL5J67Wvb3AA2enKNHOL6DvUCvVT+G7rWHg
LhWiEuX0NqVL6qrYyLbEj4c7hgvx2SCBELJlBCeqXNcC8F2epAvm/qPB26Ykwpfa
CTMWq0gzJNtpfAB+DnUFkZA+mULdhfSSfm4xL1+iWNMTo3XLd4GYxk7YBfNIkQ8y
Mq2bT2+taVmYkcoRpHmA3wY0hjUEfsvCqQsgiQ4CKOGGuXhXJZHmhViHZJuDjjGm
6Ar4/2zGdRM6kuVhO/ny2gYi76YBKUlEiUtPZhJoRUZH1nbWsiPlMEy8CPhwuO+E
1/YVOZyZRdHGAmLOoEIA0KKx66rs2q8jxaEJmJN+JXTuaMSRhyzFqutWW/lH2fQ8
y9630f9hNrxLdORY955w2q+AWb6jqmPuaT0G6xMOh72ji5VMe5avRwV8ysnBnwCh
fW2a8v2gia3DjZErde3cHapd7halMiZiMiDQv/Lgu7iym3SjWDH6MJOuIz9+zGNO
3iCQbwOHH7o5hh91UCaO4l2rNGinXiOiaLvUpj5277ccjCYpncHckQH4FZgmm2gT
pv8aggfVoExsn89HO+5w3cLi7vUKnhBfi5SmdtU2sYe7LVO0i8egcvxeGLQaY6kd
X7CNNf5ay1Kj/2B9s0a6dunQ5JSPBVZrIGQ/PC6uQnGzbyrzG4wNXC39hrtZvAm4
MN9gwqZL47jCz1wXJcvX9q9mrhc9U192i7m7jX3ThWuXuPZVukbSCDssXoFmJYtr
BVB4E5DiJwxly2jCJCGeUjYrqsIeFhQXIRdwIfgA4nH8Tv6yjZwBg3S2Doip2peX
cO0QNSpvWV1Wr14WyA4uH4yINbvYsQTnLho1oFJk7qO8iCWJV7hsBn5jvALqRLXq
tC8AyePUZVkDWMC0cW+2YvP+Rxly3nyCnEJOHel8bfdJzpcG6uboMt4e9JwIYVpb
0IxhiyS8o2Wnk5ugNyWPzWv5rwCPRln6kWangKGL+ZIJA314rxSfYEaoumN13q8Y
e6LaMTGbK2lty9VtPcYwYfpZlnwohRowH40g4XJQZ01fQ9P17wwbjoQ3HrSeeQQC
RWB1Ih3Ta3NeAD7TDAl9sk/W5NtUNUdEWi/IXi1GTEVSwPAav12GnmzSs5y4MtGO
f7pL9DUtK7fhMOjJh+5uZwGeRB2SlZ8A6N1oWPaexE12InEKGhLg8KX+eblnG/8B
/xJRmpNJVoKV+7MKl14yUVkEaW0sWg72QP9ixh8ThCLM+yobeimdMKw0Lu+u8n9w
b5JM1rIy9V8Jlrfu1biGbNMV/i8KfwfIm1/ksrc3tv0Wv0TG96etLlKqDnMF2jII
BNKscNzbamuIDsPxJBmND6QfQXjkrf8aT5VNm21HTk6tS47KeOGWLT5h0/aXsGeZ
uSi1mAX077A+9qjNPSxyqmuDst45fdA1UU8m7AqKYEQ3KUy7iaxtqlUJWZfioUyl
GEqUOVZwqGhrt20Q8DGBV+LSuBqm4JrXoWOAC2dnYoikZGwkeQUtTnq8Kfe4wG6q
fgAzs733Ih3IKS3tC5mc5v82BUrdrkNTkTQVejS9FH8COYT+yPUZP4hlJZElTrLy
4w1tjZ4UZ39ZfNbNSSCtNO1Tt+LExAEhZoDzMqDKWIhXybm2Fd/rYIF5C1zd5F84
gWSAA03NMweLw4bXwo4H0YjLLKJcCriVQL8NfSXTAKvOUw6fNcNI+32KyeeJFtUd
FTKfZYDJS0uLESL4Ih0QDkvEmIDE9DOOg0f6+6EsWsa6RPRfcbVs3dwkKbLGiFjy
7uaF4XadQMppJ6bOs6RBlFj5CQPbSzsL6dQzWFjtTk0wLGfzz1Mvv07xxyGTbE0K
OO3aZc9EkfU2DvvOfQhhC89UgV/nCuTla4Puwn2Mr5ag9VO/CmN90833jdRpNEXJ
4U3ufkywaMGqiPctEKsuBYrZC6yp11kmcZG8c7hwXeA3D1lDWpeWlZXgYqSo345k
jsh2m5QtsgqTGJjgaltIhW3apgy0seoGl9d65osHyNrdi4k73yiWYMooV9u3hazl
DGUK4dfVu4ofrGzDMWN8dQjjObjG4qicNdCswSOGAfhH5Wa4m7zZemgLWIus7Tsv
eD04hzwFYFlfssC42XaiSwdo4DHXTmloaDpdFjeYD0dc+EvRgjaRbb5a7Glk3zJA
Eq/o4VABaCVbb0eTj5HgSKejsXxGv9i4GZ/QX/4TufUtpi70DSoe/qy+OL4CNcZf
NyzYZ67oatKMJeHUXUkIqrdIC5uQ9zbVwWcttn8u8ecHWuD/guhEA5eqHhnuw4UB
/vKbpuIrkcyQvsrqagqkAzg3PumyvA8+/54o7aI63ObkGpR4UpuGWe4KpMSJgiXh
AOkZNftBcNAJUv7jp43K8Bh72z0ybt9IoBr5Im6BY421qqGpJ20nvJx6gfYyyncd
LSdBjUTwdvUdscyeKy+d6stfRxAkvvy+n7rOHanR4cfOXpP1fzvVMVgqDKZunkVF
g3FKK3K5e0d/6ynm+GejzwdrFTNSmZgW7M7HXXkYzRjQRe2h/BOq6m/nBfb9mqE8
dS5UQEoZfwLKd0oW7w8m6BZwelckt7qp9Zs6zoYDSwhGg3xrnQU5h+8KKGu9vTqk
mBeIM4eQJv/WiqLLwW/9rb4dOgimvwXA1DOqnECFFB+//2IAiyNt/EFEHjeNayfv
rfrnB86OjodRHYlvtdSwku2WkC8CssG6XDypb3aQPFhLJn2TlQ+bijduEa21gK20
389EBjZZmxCSIYQpgxR4xLr/ejGv6tw/HIwph+nVQtUWqvuTHycGW03joTuok/r3
qBtrj6e10Y0fZlhgEo7p+RQRuxGePioRvaVm3uJFDcnLhExzf1i7TAOpteU32Ir/
sozeqh6JuTxEd3QWQJ56Xo9uKAJN3HMue6vXGFXLNEapbPd0TyfXKCfgf74Vl7/t
rBeMAuznkI0we8euDpOVJVyVt4l6VP8CGGWIEjHH8wOUXDJfoQoEzoZZ44waQ7/2
8jn0l6fBDMpArSdQKpyIEDTgN3hzGTer+4ZdEqUT4/XLiTMaQOcZIj0a3iQ0xjaI
MznwZWHCdp7Kjo0MIL21hfFUP5UExSqOptx/xIy93H5I9wm3TYss/ReXVzNiFmhE
K/AJg/Wpgj6XbOI1eKeISAVXVT2SkqXGwdkXGnHKpKZZUwXP51q92mjZev/EKhfC
yCKZjs5hdyX/0XgY10zSXGoskBsYurY/dVlZqXpKAaenD0owpx/AwfvEtz/DFNda
/TPwROVkRjtn8jbtMFrOHc5TukfKMW4yHumbugjoO6ZiKiI5QtCp5FMMUVnZ/bxk
RwgmeCGBDkzA76stG/ieoYH0MKowYzzah5sG/H50PyqkPfddC/q9wSwe4EmyOK81
za7Zeqiapzumslurupfm9ZyH0tAR0uKdiM+stBnIQFsSDCLQ/nULxsFAogTaCPdP
KowAkTrrdMoWfe8zkSJDQOy1tywoLo0C0On4E48vQ2e8PEs0d1JFolhmVG+E5OBI
RrgTdC2IZ7fmK0vERJHltyhrB8kRds5qaSTj3qxvtVXC+OKnG76fmhxlruL+za2h
mYQMRg9j/njNxxrCmr3WkidhIGTfHXZ2VZeh2sdOXrmV7+aUoJrPmUTRIJ7iO6ou
EypazTkHe7fnJx5pSRMZBX8EvjuFVTbCCmpc4I3Pprn88+J3fnhi3JHCsuxZv9hW
UQxSAq+952WoOU1zedbevENsMzWskYwrkGO71gg4iaoqRs4/z+Q20iY/Ub0mZqvc
b/GHb4vT7ZhmwYqVMxGWpB2Vom/ofPFjkitFgIrS4v2JJp+qpeCZSQPukfo6ul1a
mSmNfnfpnUZmEYDAoBOh8KiyJJzA0H1gm7qazcLyT7jNGwJx64YueN3p7UzmnMrH
kuptyhUJBgxN595QzfGusAd8JksBejyH1K26dUOJvMgmrnACE0XDDqoXwIo28aqw
v2k0QtrjD1gpVtNwUwuxD2CHW9iOhS/k5jp1txic/Oho7tqnyOuSpgbJFu0L1bWt
Q+eW7A0HwwfvxbZGnLk78JPVhJSHWkyglEyj0ZV1XQIItL7dCERoFeG0WnrAUleO
uVj0Cg9dBbgiVB13zhzvGTitXdXZ+cZ50XDodDKu3QYgEY12GAYDW3Ge3ctFUC4d
o3JvvRbuRPtVKtStGTMgXa2HLns6cafzYWorNybTLx0tYzpfjZIvZJmGJ6lsJJ+7
vQSAI8ZPabnsskjMPId6EzfqBV9lmOA5uUgt85LgSP6DttsRpbhaTiSESfRDYab6
jUK4JI/LnK3ZNb0q8vwH8D8Ie1LhSkhMOMPFE42hov7FZy11qO384SzPqanHGkXo
I4s3PkcmMmhhDOa4lCMaS9oPsgPzOspzh5IFWCcCWRu6kEYcNF7/uf03kzBqX5x6
UWhEzyuUF0US4LdkQEBgJKRdnUehRtR2+t0G28If+yA6p7RxYGS0Po1wWHqgyGfO
NL3VcoV7MwLcDZL1O6vxf4K9mh7yDYCTA/65iCEy2eiHevRaCenmSAq/7fGrQlVD
0lZivl0f6Zkb0VxbENaUzRjX5wGcMxgasX6+FVHbs4P15FOX5iQ+iO5KQ5wulMJ1
RUmwpC/Nl/xz4dleNuyRYRK5jm2wst8AcRqvhPsAn3JLaBUK5pT+t2Gu6W1h16OI
XddAbyRqustTSot5zRtJZ7OqOL86D5J1pMNeTuh8ZyT6Xd06pHHDBrZakZ4C9EGo
yb5oczNTTQ3tp8giNXZ5zNiG/nmA0wM5pB0NymzlsdDvQ2xJe3bHuNggeewoZnKi
OuBqC/pev9+L0tZghtgUxV9PQjoIgVtzdcRMWOKfx0s+H3uawZCvjJU2/3P4e9sL
xr4Dfn/lZrU4CEm2fbnuqeX3Ty7GRaeuzk5apdRZN+c//f6BNSJ3RIHvdLOj1vQh
Uh6peGVI0ajM6m5OwkaQ4w4Mjq/9zCATAUpdXaT0RfroSlq/3g1GG7OpzDXi9crk
Jfh8LhE/EEuwKzG63S4dH6Ppg9z8uyu/KHm/iKAG2AF2P1QQGY/o+Yzs/sGFh+sx
zaFZNeL9Z35UmaMqW+QXasPgPF6310vhyp/VlARVfAc2DwpCM3+gahgGyhKJQl3+
1JzzxdqomD2YN7lrvbk2E5aY7oJoedSBkpP69xqhebKO+KyIMtsk1RCjEXVDGz9Q
sIAjPrxpBKNxkP52VPyT/5vTtFQ/xU8xZnFRhAZMiJm6IkkFFJ2c2sH9CQBrmcQ7
8lU4RUJutzQd/RxUjATxo88iAGBiHfYqi6nm4ZxY33COp0BOLn4uuOb7XL8cxn7B
ARpGkOurpvyGUncj2tQ2tjCRj4QrPNRYCfkH5PP8Q62WVD8llBfX9EwuBJ78Hz15
BmRIAkADPDoOE7JlDQHd00WVyWEKToO4/NoZxsFbwu/yvx+QhI4SoBU10kq6e1jz
jK3VZvWNr6cwmib6gMaoxJGhqc26wXARPCT5+cv5gMDBsJOpoQAfnyBKQ/C2jIXu
Xq9mK/RmKVbyuvaDLxRHvEm7PmOdP3EJvkfVfRooi37y+rJQ/6EKdSvMbR10/zSR
L2lUnkkv7eIjOqIBQMa9E7Ynn9JsXMb1sUnl/JiQl7zekzZh7ShSFGavEpQrHSuO
mIDSLTwHrAeYAGqNaPcbXhl9vQRUOVnDhdz2KHMIzPhvX/NYmpeKINxuumzPcY4Z
is/7/+LkOfvApnMKpwjI/veEzenvPw1pddOlF/e+MJty4QvL7EtYebOwc6Cet2+l
QdiFAA7Gws0C2/1YLRONB2SRtUVir+lLyOGgz8Zj+EN4iSqXTcq0VbXYTAvgRGV/
il3nlDlYhCO55UXZbDej3r0FnRUTBzSwKeyLAUkqtDKuAixy3/KV9CdnrfZoXdyS
iGExDfn95HySUkgaqchTAGX+BxTT9beMN8mi/Ia4EVz1YYm2Oh1rV+yheVdkUg3j
QHBm3R85xOemHjsjbSKBloaIkMt+ET7GXqe0OLgip8XwMpped5YzMxIVwEgXmgIG
xpGtriplGsS3ZiX8iTDmCQErimuFSIlDWGyXj1Fm0GrUQxSF9dkK0B97w4qZ/k41
IdPy22vRWpvJcf55aZzzfP/QVb8HNihUGkXev/MiapMzMT+ySekNEepx4UHODvPW
BQxs8GsKzRcMnTfc9wV7JKawMnFhdNFIgEMC3T751taj5YeF2LSZ334UIDeTbFBr
yKLO+EtAkZLyK/Ia30L1CjxOBCTGVuoL6OT2QXBx/VdIXhcWrc7vDPEHeeJJFTRO
3pJkir+/bd9TECVQBAutuxe+iA2Z4i2UjPm9nflb8mf9mEEBxliXPXBA2bTxkOrC
QwcsW56LvEeMKy46z4W2SW1BT8UW6FyW7EHk5kRb8/V+aWQs7USl5FLVY4aT71L3
5Gk8ni7LcA4r8UiEOxe/UcbSehSyoGl7AP9VHv3C+6v8VLOl+hBV0juoTr1UTz8M
K5uOXmiJXBLMsIu6JpKEcJbRIX5nSme1eYqnsTbxghUSFnmF6RA58h58Tg8xGv7P
dIEAJmqQ1MloyO7TIpdmUhX+aPLgEp5wzGWJvI75yD/yUCWCTq0Ru25bBtpTiV4/
5IDzvxMaqeUAmCpNaU8WAzsL3SXk5fwEXYY3XHbBU3icqfpOM7t0DKpIK/WLsWpV
4rG6uN+ZAId7xBOy/PZmDVX6t4k3xDql3+ZaEAhoZmE9SxmEq1qoRl6K1ynrqmCN
wt1cE7+1VADDuMiP5X2rFQfR6kILrkbx6NM9h0k8TpbsieQoD8NmOi4x6OMJSOFG
1p9/HWPW6CucdHymAk0ZvPHCTd3nsBSi1jJPrxAUvRtQSlgX+8r267EAD8InZ3ww
sCS6UxFWbFsAQS4sYkTuqcgAnPR3p3oL+rmgOxTu+Ga3ho9cV72ofQ1t8kFrSt93
PY3NyPIcp7nTxGdbbxRPUqzmH/X+gNqcH6P4S8b4ze3KBSJDfY9UyJjvDIIp/EhD
QGiAzdCzd5OWPxy7QVXMV3AwnaYz+L2I2N1rnm5geOpOJnCiXOxJZCSPnnzSqEI2
oB43yJZMM+0NxGBBGLQ1+r4uWToPe2j6PYdJqLU3DqEvqVUWxxqMPj/5A2XSlm/d
eu1jYZtifQnWyKOWmc3/tzHYFU/zjD+qBEABiDvX9miYSobYgU3kjG29AU04xCPA
YAfVZCSAX0h3KuzS4Spqg8A8BOgEtgv45SpECIqXCnK9hy70WNPz45eoT06wA4Ks
PZslGhYVI9bYmd/K5vZ4MUg2hwPeddM0KMOOs24ax20w45PvLCouJfhGBdL7+Ahh
EBNyvQRGhe9rayW4cpMF+3dLDfSbpBDievxK+6bh4qY4mp7XpuIcxe1qKk4jHtPj
sIOP7YqjOmp9DdMHA+liw3DZoJIrOfaOVX5XdZtibsHGm40UlbKtxjgPAxfALg5a
e3FryjFfUJoBk1DRm/hFBmONIXtGjimL1drIK7n3cCWnGPzigijlVeQHxyhJET5X
vfHRar9LN4uTawhPErlK/ah4KBOxmwcoNaae/qlTN+hnOfIjXylrOXNoigpswxWG
ZubBD6CqlUVK+jgP19Z6TAllbkm3klp6xObsci3vt4JgEmeW+KP4OeB7DZ1usLYF
Hh2/jjLDFHddOha8j9nNCvEMW7KuVe+a2ApuckPhFLmwkfuRm4SzOrNIotoJLiIS
uRlOdo3tqgmw63ox+hpJcKxuydBQ2hoOSSbAaDHiSQdR5UM93Il5JldN5rT0XW29
WqMAxrCo8+wygEFKfLI5SUOZSeDhGqEej+tvqKaAKd21ykNwI/WivNznHxAfjH8Q
YYdJHgodyPCyOEOU3SgjFQvjf6YEHSikIAZFHl2edoJBfItuSPv8gN1l61+T9WgE
Y69gS3pRmC/awzmBaxaj3IyAo7e9cI9r2Z1gingauUeQbCZNXUyjSdbsqVqntt4w
QmDqkgXLjbnn9HPsjTKGjv7f4Xt1unDMxlOcg9zcXKQiJxaxd2QuX9L4GhG1DJgj
ySUzcxyFgPAuNGhlB+afuDRuhMQsy9w4ksRwz6dSK88LkBPF46o+DNp+ZoSh9/9i
oQ7TC5EmJui2hvhCpdu1qvA9uan/3PXruOBfsbZkfdH68w2q6BaLAnFHeD6RFp2n
4LEJDyIDk/cZmgJTNwh9mvxQQ/eE3sECp/Muj1qCzUqDjhTiQPe+XTdGEmce8N+1
VdYHSeggAFJeEbTmRJ1z8R/pe5WyjgkIQvdTHzVeMXopw7nEIKkcEEUD5xb1Az6C
IDBmnOGyoPXmHVpfqMEko9CbLU8wWqBiJq1rEMuNJ5rKWqjcYtpI3CK5o1vrvJx/
+FivkFsJrE2tCo53nQFGZL/CDm/gHKj52uEI4IulfZnWcuaNXiuls8RvFVZ7qwcl
Au53h0NAVywmtk/IIeJF0FFmdQIYzLWyysMvnQrW948PSZOeZGyqLJCunv4tlaWO
zARnVojMklDH3dpKRaEsa2AUgSBFy15vp9ADcMCCNMn+/Izo7oGIdZ/eAqyZqVDB
+g/4Lkuw9t3+sVpHilkjDrMIfbKCy+HngVvJzV+XK7p9DAkBEnyYXZmOfDiN7pW1
3sBJaiz2FwEKlZpnTO+Z3PtnpJpHUlcipnRxBYjr0E36UV62dzzDj9K0bxnayGXp
SFXqjg/jkIeaNEG++nU2YN8ZceCc2Zz4fKRzr3+RAascA9JlwcN4fNkW2FJum4Ib
F3pcrhgFLo1+bUtbjeNIm+45wfd5ei3V2V7dJXMvS61li5j3aZssho9IFmiclvCv
I742nf0OOBCnkG4227v3Mrmo2lmwGWRTCmk+gYnan7m8M2hDBmu/xMGVDtYa6Alo
ePNfq4ZaChx2YDbcmt9lf4jLuKgUeexyOHwVq5UAiBChlt0HE3K4QkkL/DlkTmps
Xg0Y2Ej6/e++BjqSiLRIyOPVdEvROFescLMM9yC+aVJ/TSadkqXXGF5zKVtejqNF
R+WAvvorq3Od+2cVUI8UxF5KtXxjWb3ea3dwcZBlsBjFlVD1/q6SQnVx2R47h1zk
5QkP8vNIQBXy3n8HhxFzgr0Ynkqc68MNUUbRqUQnnaOMcMFVQGgXdctZyU86hOxt
qBJs0tpKSMCTbvedI3+DFirPBztfvyqX83HnJsXrYQ+FtcpLtqCPTBdT7SHqbDPU
6ch42dzwiMq2nOthQ4YSX5+uOYE7m4XKbcKYIGzT5CLq/rg/MDN0tSMLSczHfDEu
No5TMG31sUb30RS4tFuQddptdZ8rVWE8LmPo7j7XlHmzoLcl44VEGODVFgT096IO
8lkYFj0/Cwt5R1MKXT3DTVL4YuLUo4WiKW9WpU1teLNE+SR7qXXH0OTcaZeJxOMm
1Mti7yRFsVnaGR3XhXR7LLlwRaz6vPfHC29qtiaCji1j9ER89zrjj60Z4FMJ7thN
KtnyXSHJ+i8HBVzvDBtJYg4L4gFcyCbDqkxhkhKO5IagjYtE+JDVgshwN8fnBTUp
hG5z62B/YJ3KnYIQj2Gu+d7h21KqybE9vAYbUj213dNgAavc6uV0K5sl/niNtFUo
5PvgZr2yE1LXiHqi2bFJ8K6qy5o9sgM5tqDjSk+yKijDPOnoKMXTAuSAspvUoSP/
sIS/mGKeVSzTfkTa/0zGlN5SoG7dVt+CiIBcoG1Q9x8qWcbFMIujYP0+Kdh67/Hu
Uer/IxUD2vYW6pnAF9dUGXAHeAuY5znC/9zZcVltNBj4PgVLl0kEhA5Yq5NXKA13
3UNA0ZAEFdTUCXxKmzeJQpwDIPWGymFkXN66eoj9LOjRatInUnJbmLKzfCU7ohMD
DVWRsjmrijbCvlq5JLaq5qQJxXkC7M1F0sdRjlNhobbx8XxLumsH7VZF/2ALu/ic
8qkmaw8kLmmfb4MheMJK2y72I/77Pswy5XT0h7cn2cDCa5qYleZjYuFqNLGQiIXV
8Zzp0QDmQnfHLz+0KIfqAWpCzn5heoRYkj/SWsEBDonepON+bmh1BcwbtF5ijWG5
0WtLckgyGs/o/aRmBYiQJbHPx8jYGxK0TLWaL3o1Q88br91u9jSSfyWgoBr++z7g
xSx3Z6GWvdwxGHxW7B54ZTBbLi31V/zUi/0wcln6oNvhAfz51XldrGS2f4XqFSB3
iwpqwacUz1a2bl5LfcpOMycVQD460Dmt6bO2t9vyLxonWQsP75ry4/+lAt3wh2eh
Y0yx0VjOqtW01mPQ8syVJejH963IeK6Jih5xopGFsEG1bq1Uc/bSCILonHUTjwv6
HORI9f3GW7+08fBS/Rt0c41OtNChYMcaBL8lw0JdDdcEJMyK7sir3hwYDyXTApCp
jiEi2xaUxjeRuItpmuidpb3Lvt0x6NllUaeE/WHcBufdtk326g0jg63NkT3Tscb+
M/ScEq6u3ILMugSmAlUOU18/vr9VxSKPqjSyGJisbq1CeWxNZyU41Vk5bnbdVDBM
t3EJGPK7+N/mA3TTdIL6N8Sv+ep/uj7+bcjnxZ5CZPH8DSedU0DLsDgQHWOlWoif
Sq65R+zlVQRS3Js7kDUshsDjlUk7Wz3mWLL3jRZ2OyrX2kuwGqLvWunHcM3TkOUI
FHjo2/PO7uo/EbTNvd2NLadFbsXnz6HwSb/2StfN1Rqy9N54chfJDTXZENrIAh+U
51vRl+HYh6X3U4aa4jboe7J5OZv3EyxKThO/vAMsLZ0iY4C0Q7lFxnqjvyjLGuWO
5xQEpcEZjNiRjDVVnzfrEg6c7DZLpYLld+FfmJS1OkveiuDry4WwxsN/1JsDPlr6
cycnGlZZBgGWHVzIDLnF6WNcDH603N8ckKxK/iW4SRJW8F+fTjdx8b2LPaRHEiUt
U/xI1K1Z0T2gP1v5ueJX/EXBdA+igZgf8L1zeYP1C5vvWO6X5ldiySNlm1Yo/2cP
jv2WOpES3y6bu0KY2re5or0jJo5KTnvRNLuUrg1OwoNiFv4/EiXh0eY+QN6zrhY4
72KQLcLtmjaaNjGX1Hq5FC8Du8cepT5PzeDKDs80iZCroGRTJV3wP0lQ7CbqIDef
`pragma protect end_protected
