// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 03:56:36 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Hfoj954dhhY8A8ZnPV/px6XRsPJ53z7ymCy6ROz4avOAkx561obuje3rbKycIckL
bAx3iGI5FW0XH0ivsSj3vlpbToTBn7HG7kLu7I2IpgucvWDivoNcjieiSer7s4W/
Zy0nPwnTo3VRgM1uwaR6IcQ9Au47h7H66m2GgXFpKuQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30832)
CIeNQffJf9zESRNYcBi3IFELmcYOK80tQTTDxI4ahXEGNnCHujfPMjNZKPLf/mOu
+geIP+KXyEQ2MJQdKSDwwwOoAgYSo7luv28WXmTWHzNPY9dQ0nKLgsh5XPflig26
xSoGew2yWWFDI9iwIFCY4svOWehu2upNXqZr32kKU2B0Xq30PGOWf1MNfRDdZS95
hs+Q0UTvOxbyHV0lVmM3wOnIGVsIJ1P1d1UEt7esK1Q8yCoxNgoj9K1t5KTCVjU2
yFcKoxUJOn2wxfQNlsCG2XAEGGym+3AwcJg7zsyig46WsoRyrWN/3cj+4+GlB7ch
K1zGSpqVgBm4dhGP0VehWfXUAliHdK9lR9QFyfv03eDazejwCstSCsQWgXXrN2Gb
l0lFfQT/1Lvcv8yDtwE8qteZ86vz9iBOOXkAVu+QdT5EC7VCwsjQ6E85WOipqADU
1iHXFVA1G4Uo4PVKJtKtNIbdXYc5IUVd/ft0GM1b22k3BK1uUW1TaKmMtJdFK+Ur
gK2k0FVk8K8vFUKcd0FKjxk9UxfxP3W9/aH8NWyRF8fXevvdwA0FewM84YLJRt9J
IXwa80EiOSOncwJ9ijBwxaVh88BC5QOX23ng+5iZqUuWB19+0k3JK0Pw2ooqyyc9
IWweiuUveRr8QogqLnMR+vRJCtrjJB0qsqyK1S2vsvVFS0YhbnLkRdi4p/QCMHDm
3Ea+KFW7D7H+jZtiaZHMI4fM63GFNQdyAV+B53Mtftpar8HpxpMfWsCeVZ+9TJAp
ULWhNwBNqwkNT7QfmlLUpCJ6+BI8SDxEUAveRouqhlgtvwSC2LTQg/un4f5SSMEX
mi0HLTX6grzvz0WUc0RyizZ/sMEQSEoHUy1uuI3q5dKen4AFguwtVy9cUnBuE53T
3OoqqSDd3SoT/7Omk+Bqq4FIzdJ96tO3UYr4bsg3XvgnDFfpFIxE76vAbHD4A49d
dpJs0V9Iv9R72/nnQnw1B5dssVygpQshBWwDe9e9hcWLKpo8deRU2zAzd6qoJNiL
8elnWb9ecJxyd/MmJymBBFRamwXH07ilCPRtU8tthV0tCpRdZfJ67h50oNzW0YTI
7VSED5qW864z/oVqkpjA4LWROEI09zB53TGAV7ujD2uV6sZ5hPhcd+BSZN3KId8r
UwM4kdOf36RVxSpZ4WKrd3RidxZwPtpp1Yv3dgCImxRSJ888FLmU2IoKOOC8hfDt
U/1siRNbCug9FSKXY0tCXAr9XR6KcJdp/USHrFyamgOgveoqICLUfyL4+q3uHpzM
2FzyCxZGY8sUyohIoiO9dcNuWRiO8D8U8dpK+gAva8FUAS0sXicBhfoWSgxJDusm
bwx9hBVeY4vuVjV51i4akBThQzoL9BCnzoZs4nUzFRHhpmZEcdQAysK+kRvpq5C/
/uHDkfBI+NSeMLfU/M8lSdmkzbh7Vej3sEtcA+iyubH0vbb1jaiWB0l8gyFq7t+2
pceURA/VBt4Cygq5t1VQFYvhfxtx4WU0zAVMYv7nK18MgrVUijPqXnSIhddgWjZj
LOXlVs52XAzHrUILS7a2YCbnVH+FXgahk+SgcA6vSRcrF6doof/WHhhDwoT3gatG
DdJaoFTLJ+LKCGuDjnz0Qs1tBTgZKQVw+mXCsIUPIMbQsLQiMt/l7vMsWzqXuiz9
iYexd++h8hzY5292Hd525atNgP7GX/yYFSivlyxB6z3fwN2kOSFU/JgW3s0FkjFo
M4SaJQru1562N+fR2kJHNfIp9QtEXXf8pq5OYqonGhFSqKb+apJKhPK5a6nnFITa
XjLE5uhIT2nlfBmGyoOIZrtgzDI6XwypgVt+fVIGv3BBuUzA9iQU/zJbls8F/HZa
wmLFmcgvT/Dk7tIv4RC5CPr3jOj/vMFi0Xd5TAKEY7aOh/bRiGiGztpdO0NZaDZJ
BdfKsBOk9bqO81QVxyIwixgXR7K+StTyXBg0xKbp0mmqqYnuONRTSBiJwqKUl7p3
d0fX9VtPLxzQYPoSmNTf54rIeVLDP1OxXnAkORfQoXvplMHP7yGr7r4GRIPLTJ7E
fpydlb3/Iq0OGpNUGHo61TODVD+Jinr7Nux4bomWBfpkQEIj9krfXC3cd4Ddm/2N
qsLH7DJXQpNt3LtJ/YRvFkc1VjEU4bUSNDUY9pGHLv74E2jWe3Qdxjx6BLiP0MhV
piZg9pS1K4Ja+2DTH8mcQhfVZ0jsag9ncpc7tsEnc1SchRWRBYuWG27DZj+igPHd
IWz7Bq6Lk8L+LyYvgZuN880Zxnim49WbYbXtz5689qz72acSKdNj2rlK0zZ7LByI
dl/NpqETXDCCmdwOOUwVNQ4OGJ5y/Z0+QbCMk9gNnZHGH68BQjmKdozXBhCUrmlU
YtGIsJ0CNnlv66zAxkN+Y9udI3B4sqiHfK0BtjlvBdhsB9ajV9ai0RXNyamFuaGE
3lMACXyGerbJNLBHbKAf83Y1BlPgJ02c7Bvt7vq/kfA5hA9juPLiUfS2QT/yE6Ki
DY+LPkS7FuWYk2kpJWmVQLoooQja+0YqVoIbKWu6rvQVpFOEiq/IJ6F7T37m5RXu
N95eBi0ErChUea11/U6o+cB8XxwOa4zCLa0QrKbYVF1sc2tby9+uypOwqbEjv3FX
zhzQwOXzJL0vIDbcxmV5Y9bGdpYvuF9w7e3CL6r+GCO6Po+nI8YrpGuiwRFV+kuH
e4M5IeeiRy+T7chQwuAerKJK8NvKniNfyMBTmUZHefMpj5oR1GLnO/G5RCu+Y+Wv
ulRNfpa+VFqNStbAo6grOjwJktHx8s/ialIPxupjl0NvGpd4R4Qgs9ROa9pc/RXm
7AIic911+EKienL2KyV/Kquzsxi0YAsxhf/IODGDMAp9t82vIuQWqslX4N/Trzzs
tJtuZ/oGVh5QtQv8k/uNBcgzy1h/k9c4rJf27HMGu0mX57PcuWP0LaOl0hYUQdL1
jl5p5IpFsfcZoOcKW4lsCxkrXXjsr05CUD749bMkZ/f3TdH+oPm8UKbX8KGfpBO3
cKtKwloUqE6oi9ToGRi2ePS1cJexyMguikOD25TBj9z6YvY6DNQepwTfFyNaECO+
6bw/Ry5XqAapq7Zzzkhg28xx1MKWoNBXDtayN8W65kfNSznQariE6GJfrhZAF/8t
H5yxu1LxMWJKqjEm+zS6xqbSm7y/vrKaFklKN0ynSNoVdsb5JmwLGyFyVq3kO7Np
6fUd6ZWJaHFpY8zVI+tU/SqMxB5lyd45ipKafI/ALzW6VbBWvBvyJk2cGZ6v5YTM
kzQpAdcii3nQSPjK0cNr/jagYxcZh6BDLeEnhK0C0kz3TA+8TNJWK1m8HVJFU8Fc
qd5Zck8PhQgx9E050hTV2LWLcC8W9nAgOhc+BpSitD7m8xgAhql1LdD8q2SjqoBr
BQERWTcIQgL95PvqFcWnV4Q0nn9mnQW5s7oZbAmNo1PcdnNU2dboben68Xm9GiDV
afOFqkTOoPprW9XCzS/bmvAhMW1nE+TsfJ4ZO9+0m5/KEN12983JtsQPUNLjiOFK
H+AHwF/9qERG0Z/PRvhFHNdQs+MUDafF7ojV7EpXphn/Do0UE+G+7N7PiepkPoin
9Tq0HQ/YtmK8lF9Sjg3FdmyTs04EFoF2iENwB6Q1IwzD6kWE5uskKxNxwUY6jjpa
oMqgzFFSfTGXX/C2OccztVAc1DRgRLyZX8wTK9YIcMaxq70bS+n4ok1lLekNfD/C
f5F3A2cOREV2lEPHqkv9+ByM8yCf0+rM9a77KiaQbXrTbT8m2sS+yNWB8W79fyC0
swTiCaDk+TBB/EJzDUaJndLJ7YpgUgQ9DCtUhN5OZOXCq92rAd5MkUZBuSODz5DK
GvO1yLNQtVtRUDcVCd2RCMr2uICfb61+PNpY5JEBu54UGokXqA0quKsxVGzGXyFT
JwOxHHVmlPvJOmHl+0fHafSLo3KJmb6Rft+DaaT/Qo2QGTMA6uCgkfpzPRcONcUt
X3KIcOxBepk359FVGzRLkrXbM55Z4+92A2UdE6hR3mlZX7EIUlGKkIqOaLPQLbQP
ko1xGtilzdaoue2nf8kaR0B52xpN7Hx4M527dOwOne+PbUhj+6yoJAqqGPB3CkVX
4sXpWsbdejSZ4IGiWUPmuT151yLG58QdNMXCr3IVGqicwJcf8/opyPZYuEaOwNYH
kQfXRAUqJKE3qPSiKot9mhkjE53AOFEd5/tr61EUuH/T/f3wTheOvvfjmor8uC1r
XMtJiRzFi/upvTSCYNRXp57RQDQ2VYpOZjlbmar1iL0Oxc+wai4vwjSfjmYUzOJ0
B0T60/1XTxHj0YWE0P1Cf4PKJ7PmqOtDN/ryDy99WT6vt0RfeMYvVvm0Y9u4b4AG
Pt9RbjWzxbuvqDxP8ZtVfwZ2TTq0PXlc5fJ5Qs8TrVWouOinRHNx5SvtmW9kYAHW
sw4lQQEAvPK/IzjI/DPxwmtGAr1cgQV0c7B5rYWYp3nYnwLkgul+9SNOgsN9GG9/
GH9GikBqKDLCaFFuSh2jOHYbOCzORZp3+T8UbaiU63zh0R2Lxz6C94qZ7cTNQvGU
4kx1ojOqmRuXiXLonGrPjdOnjk8FO78zXDefdhulkZ18Sihq0jte4f098eTfwKuV
YuGl9ksCrRFi4B5W06nGnG0mhDm2EWLt8fp/6cU+fZ9GQLGBCzNc+q12b3KJGoSe
5sC864pxyMWFYz85Po/K3M5/s1SDDp13Nvv14UBvZ2YXnBpghtDumrsbhZojSTnv
Zn91uvvYof/zi9Y4uHza7rO65eDQKYzaiEkBdyLDU716Po8esWvwvubYwNXlFeQi
r5OyjeSCccamBxqcbFSvNYlF81uHH55JubxyNrbXAIrxAl7oFhNV9XxqbXUA8DF3
ZGI9cEnwGdlKWIJxm0ozQiso3s+J4uv+dN9aj/7FVGcTRYpMuRx93Eq2HoofaSMY
rfQMumuB98s/gPbwxSp9YLl1+DyTmiigtCsnnHuUtHupzAxHx23xo2jtHwBYS4pW
cnk+6uWuvssO987lrMsFgluRi/nYSxtaIW/t+oiUt8H46r5xWONdK1N3hmIf51LV
bhpWIIFXAWheJ2nfTiI3sQ2eVYgK3WW9r4eppmUi4tqlfVRsv7KNAbIs0GQR6k+T
X8jblP2q2UDFEy7nZ9PHsnYFNyRGxDOxmYNVszGYIdJ6aGibF1yPN33BIBPvkKS2
1V4WzggIFWyM0DllAhmgSkRyKdxiadChFkUbg+S1kCLuDCi0F3VrQNb7JwScKu5K
FqNAWPWMvCLdKYk4u/AX+wmIYf91agmMGAOp6uR/Y7vBflRBgCIZDMTfH5c+iRvn
S1hDB25PTurzxgZuT/i7fth+BXAiYbsJJcnLTovblTRrnXJ9ivBphG9gjHxikIOp
AmMPHMuUnII/r9KB1sgiDvJVyZ2N+yRPdr2++gb3dApdb4lrahbLKo2dN40zENZf
K260bKNKVDzUMvAnI/hXXDCBk7XvYxDDodZFCEi2F1VPrmdJW5vRTdBqs4XUy7xq
w3KyQT1KrIgj6uZevB/yrh9Yq6sza6mFqxCAVNv6t5bsoUES+YfkRYTVdSsmtrkb
BcdB3dmlLj3/eBLyGszFJbVP1I6jg1wSSwEEVGO5MY8Wj+l3lhOdF54LbiaD/EXW
LRlJRmoatLthyn0IPLXF3pKj+BWPMTHDaTbqhsOsXloy8mnE3uvi29TjdAF2JdkO
pOrithFr4i/9Zq6F7qufrvFax4bJl/5+5CGbqkliOi5rW0AyxXCstBEqgHeVLNk9
r9Q5hZjS13oLPWUwZJEPlxSbzKxv7k2r2GTcoXWXKy693JynDC08W4LTHDsfdVTQ
ZsKqPi0+P9h8XZOuzkaxEUZlMueKk0ULBMrOhkM0BDIdXl0Ft6pfETxO802dvMlJ
utpLdzqwnzEMm2HXc/c6ni/ROosF4lwFq48DswmyfVJf36MaEcJKkwxn8kxqxeOk
Rai1uuGolgi3bI59Tj5iul8xIHehG5XO3EZoBJRfYtpB81dAwe/4mtVERkF6rNul
7wBQp22Pp/4EJ+UgoGZF1SYLnROybStN/s1JbxLcwfxZl3u6PlmpcxdmWG7XADa8
Ei1RJUYZ4aH3AtgVqJjN+kyvFP7t2qH+1i3fiYB/qxq8A2g/BwDPaM290Y9q7nKh
75sd4e5QceBYywWaF4N9rjrnnxmNnAld6bcQPOISNbyv549V80KtxUdsZCqzhNZo
lMv/2A4W017CB6/1pP+OC/Zz73P27XqaRuFyb+Evr0lCZG1DPnCb29K2dAfHoqMp
VDqIdFVsM1zlMC7vYEZA+a5cMA71thYUxW0kD26JY8TjAo0YD/r+ThQtlXibab9X
ynH35Fo/+zpSbcqBFnLS7BGTH9aymSliysvFRB5w/P8J7i0HzSPsN7Ab8mguTV9V
mxMVZVCjEHWXNSHV5BihrsyY4OcY5R3dg8Y1Qso4gqGGBPEFA9PXJKk7qg6f0Zhy
CcRmSH1mtuFDbtgTEvGd2wubSyz8HIU7C1vrU/Ifr/Q+gV3RWtLgqOJJ4Ld/7plQ
v4f6p2gEXwBJxrOWkvgeEhaiqKw/Zi7FGIhKhY/712q2AHDDaRWehJyD6Bz8jOM+
GcJUbVP45ep3iX2UVOLPd4LSbg2U3+bqwvFEXfs0ZYsNKaj/SJHL2utma+RiMhWE
WQ6I+cjyydTaXsK0qDp9SkedJcz5uLynKMk2SjeQtgCmvY8CnvXIHv49X+gI0c01
+eZOfXGvZSBvCJdbPRIQ4BQvoGPjZH8LRu4LIv63NxpDtT/0J9L7ThiZCuBtMWd3
W4QPtcxxFwmeztS3zVAF9qbWjQL9wz5LykRc5K8Cdv6kjoQrCs9o9R4ixikaC9EC
QLt/h9oW8OGvLN1Gvv/hDghfBA5XHEMHDqkECj4L3GRynEZnrk9J7C1zI/08JBhZ
oU03cC7By+60w34jjWL4b2uXKDAcZGahuSRv1ovNj+OjMkabd7AFlEm6VD/ipnjd
+g6jUhqas4DHWBOz8YXL1LCYQVclHZHWrgs894UTG6H+vQodLzSeyneIzwiiUkQh
Sw3WGxvfoogA1OSc2S4Nyy/yFRMmLDCX9GiC9G+VRvcUUn+iHVLZI2vlkBycVEPC
luzM9o8BYaCPR4pm2Kgxd3uPisO4VSAWzKNYHbtNl4Sl1729U0SuurwDIg/BEPjk
RpoNDFlMFDBF2cx55+xeb2OCLtSepHzMPOW8H5XeYbudxq/qV8lZqWO5rWWgVi2+
Vofpd++guoEendWaUH8U0ppKuApNN32F6omAVydr04GjK1mm4wJHcH2KAGMT48Cc
GvvrcZ3YCUwFHNSfdfvxqm486e1WAxa2z/+OKfjM1HCFNqoFmVyxQiDxlNE1Mqzo
u37f9Oj5suK6g3FRspo1d+Wq33S8ZokwTUm9SZVJekLGi4VFXAwSY0ABqzQL+e7f
hpPDculmrN7m4qEoGNplLrr3Z3It4RvPjCbbiMb4PvNqPlEla5F31fav6o14gdo9
HkJRy5DBXzJfPvt7+k860QtE3r5M2qCFt3fwII7xtIZSFr0LAMOte4wlH6F1os0f
tfPYNIxMSsYPvzoizg2eFc5iSuP60RwVJQBSE7giVEIQ6NRteRQhTp1ur6Fj9+iv
i6Jh76KrYtSThQnAFgJtlpmc19gEBj/23QoH+HIoxMbFHES8vn7tfS5ELXyAB1v9
ZrE9+Y0r1uv0/qSugS/w9JnUnrY4TCbcg7R5vesTxXlXzQGFeDtLSHkfLLt6N8rD
JN2dqdNKO2YS1Gvzt9rT4i7jKbsOO3iknVbNRHgMPgbFtdIMFCo/X7Bnr4hbKaLZ
4WZtl0aLRuGZfyQmXDeq7xi1RE7XPGK5fYhToCnvj1lmLriG5tc5Oln2TERcaoLG
GIiQON5n+ns6c2o6ABFUl+aGusgGTDH2MqUzlUAI9XMU6hp1xgcKae9/7u84uIgH
BqFdZYCb2B8N1+HPH+FXnoF06pJ2NA6aMSEaJscEikzPV5XKL2np1XWvn4Blq74k
QKQ5cT9R58NvBinAiddtqIWB7bCI4X5YNUqwMMTjOQfDCSmwKC7GnqnEjhHR9pTX
63bxg+884FjGmVhMbcRfm7PfBTENLALXBSNtjGkhqwViwaEh316orNNFTB5qJC7p
ZnEuBjveu+TO6zMKZqM3/oji3xIRqv7k81T8ShVZJZsdDPQaOBOp8uQY/pj2YNpR
B1h4ZUedSSnojHxiLtIAuOCru+pg896LXxzXfb4cj/XYNSWitFLXC//WvhPcj3pZ
HIFC1a7FcqEZzJ8/nZ4P6VrMV2KpoZS7Aylq76OYCwDE3Pt/nxiJA8L6EBtFsXa2
uyTQVK/N5mKKcKg5uoPdUMv2fdgTWXHz9Gtq793J2hgn1QDnoVaROb+reQ9rpKEx
QN0ULeDLWkjwk6t6j3wIdjMOdyRrVHN2qMSXt57h3JZQhBmvRmYsl40rDS9PNpmi
dXdVr9l45T4aO3kiFNUGiiO91+I3uahFLwX4eUOoEb9PqhwwWlXnzkgaqsospd9a
AmYgGvlqYq9R+4zKW6xvO6HM24rLa3WfPaAVt1DVy07LozOi4heyeNrCSh8LmzM+
adtfSgVJachWG86oblQ80jGwjL/HTaNJKDc0T0svVBqrU/2NtLKrE4xDSETjITL3
7KnoLxngeB0fEkYimi4MdFeaWBCvrNjxCYHusGwnYiWwWyW/OFRoy5V4AX86rdRe
39RYY9VK6wjZN3+RQx0y6CVY1pQCycQT7tKEBVOvpDPben/vv65Hxjsl0OPwNvRy
NxI8J1Wt3NrdOJJzrwHRl0edmTcrMepzxAKTw7e6RbeeJbu6OCbjHds0awNOlhas
hpeAQT54IhKPAv2U29SGq5/SpLuAcWwgghVhcs7a8mc+l3PenvlsgqeSLdH2Aih9
XksjnnJ5pBlrDKtqVpt4HpTh649WfnFAQpUWNk1G5Rac4e5Qohef3avgZ0X/v2hT
kfKZZk4ZUymptlhJbyrCk8RJXF/9nMTQCw3QWStcErNTKQyVukcWM0edML3XYaS1
1esZXRLSPu8vyTYqffUvXKhF2sQhX4zi3ZEpedYjxKTFlSn/t8UTDXmOSPfu/zGl
58DKoGs+9nHmM7SeNeGk6s0xKsDOivzJm0N85nWVDnyaRx2QJGMmuUnpg2NtSQRG
G0IBhBiHOAI3IU8DDuaEPjC3vGIbg2ynSSGoMgr/65DmbDTo1BygdpI3y8ZQPnoV
WUH9dMzPEeXaFB9bcOSq4yOujwMIXFlUhOiEDrjxcDtbNl400J/uSFwogdYIwIi8
ixPKf4k7iqDNFbRKCSC3tZHeRmOfPN4Tv8uYTg3EJZQiONrAxAMRxnF1HHBb7EBz
aVd4PNM8c2ps4NWtynXHs3oFKY6d1YBdV8d7ymtmGceFp5rQUrRfsruYUG+nFCOw
+ZdCyg7pLRuTWIVTW2gESyYmGxfjlevxypHikxOjCbomdUk9DrCiJZnWmysDXemN
56m9tGoBitmFAT3niV/4Kfn4fTCOOwVuyurz0eS9PNqwNhYGTD+TreIptpI80xTb
JD5xniashxynsfdYSzvuWYv4AplqbbvR60MieVGS4xrewfltWXPZxViJPRJZRcxW
03vePVrHERei0wdGK+cNqEzekl73VqzkEA8Wudn+huoVH7JpJ+40O+FSXzZ/WUi9
wLI+TUgpRyHWU4GgXuXp1fAPYAV5Y9XRWYCaET3I8VnzRNZk9zCR2iNYvkrmn/R4
VyO7HF3lamkgyP05s3Eco2mshxq/NA3GjptFinbv3D7ppun/lIPvpzLvf2Jmv3TN
nii/+qF1VLNhVot89kDwEDXl8vcgWTxJAts/uOhN8kQAiGjYkTP65nDlbHPgfG98
W6LK1cAmFiWd/tKGJj6ikrhnNdf3oxX/C9ScsiLytgjkkyOcbIttmxK+R11oX/mJ
yYBvR8I2HS6Nh3dPI78yIfrSjyKq2OnJYdxjhwlkax84wRnD/0TKhvhx8nNHexhj
JT4oF3DIzCXlr1hUQeSCjBjmti8vneRsa/sXFbZMOBV0FaIuf+pYBuDqLI5ScdD+
ae9V5I3TsMrFWERxbKf4tz5NnLtL3cU1Etg7Tp0n3E5jzoGp29XY5jeRXC73/WOz
pkkrQz4GC173furYmXunzkboUlmanVbMi3RdfwIUzRrnJaRuQoTZFEdZ3k6NEAkA
gHsdhAl1PZCpK9Tq4OihrK1uEAd8jn567WoZpckD+O333Tpjk7jDlGMKMES8Wew0
ReNcn2lrXnr1xH8HFrfewgJTjZe9Xfecq0EZ5iLtLr693YhuJrkyhwDhAOhUk5rn
NmQNFdQOigJenB8tA69iM7V1LrDIY03VFs9ETJUxYWngh2RPKNiVw/p7Bgg3W7uz
azJbRYcwl9XD5V2Y+PWZDz2k0CwQtlX2p3DmsgkXtOZm9XxH1AjhtgG17u2K3vCd
SK1xLsWYJyqQi6j4K76mI8PqYVWr/l3XR7CNrko2pbjXIzVa2S0W498ZyP2FagZq
8cUdA4Tm2e8tr1qltJaPHDUEYDmuwiSxzdxG7iIV3NAaSRu8MBNxD0hv6JddiFWa
AHfTZLTgg6dxrJUIDjThw6jRdL803k4oOGwInlu+rCt2qMCaEzpLjaiIu0Habe5z
H3Y+ViVmFiQOklAjSCv+VtD0y1jR2ZCE4ObGAXECwWSfU560sHCUn9atV55HsIhB
EcuEhMM4b6fsYOKFmwlc7egFkW9l6vaRhn7FQgUVyaNdphc73z0YxgY7rukahh2b
Jx//h8flD2sc+61NrFyw1U5nDEJptQ7XTji8uZdT+mdxQphFQmJq8BgO69q6IiY6
l1MKH7psiT4erVyoew3Fi/q2UPG14qBO9aFyRJEUYf9b9/0NMV93aPwvYYJ7y+lQ
WBv2DXjLWYc6sIAC1I2pMs0iOKxmqJAcV4930KF19izrEWWU29ag1DJ6c9H8jTWU
WNDjRLcN5dBCyyM0XmHn82DFQ4DssUKW8CjOQKmDEGxZTLfZ5eij27i5oRHzg2PC
5HdhEUuOsNKqrhjEb1UoPZdwOqoYxD2cuROnBe/XQLBvHbnb6Vz8/HB6DTpbId7w
/IbbFFGPaZ5847QCuc2HF1i8eUQ+vPQcm40y6ePOLgC3FZyQ36+D7DsNRcBHxhVV
njAABcKzoESMpPKhsELVY5v+2IWMzyf2w1ejq3UPTWMNuYuVX6B1xx+mB5R+WxdB
IH64915umOs2bvrBjNtARu8jym3XYkzKGX8xd80W+xIhLN9rRCC0GbfWQSxg1i6y
vXXQiySt0O68/pKxDNrEo5EQ1e0FUZw1dsREnIj7pmpnJa+exsp78ihQlY9i7lPe
OUwzRPbTRrGhLabJO5IM3tCce07abl862xF7B4fvJBZeCBKIojSVbT1Hvs+Dkhnq
PfQxqIUY92okbxhZ+F1s30rwkszia4EAwZl05T+/oAB5JJRxkiMAj584gwM1KY9b
wbPYmHMKfPY50KoQPT/wrkAm5/tDeaH/qHsRjXWN28TPbEq1mdIG9aGaAlRzoh1m
sYsrbrm3fNPRaswpmiKmjJalflrcdX8dot5fdFDOrUCsDfCBY83L4xrDHdHr2Dz7
l3X4pIQIOeI7cmfnrvtAbgWE74MV3B4y5PUQiOayM9N2fXLos5vC3sRUB0paBvcP
E2yTMeL2JBnvl0bhTd2y1rbgrB5mW7PAhTHFaQqcX2oABly0exq6Waj2MWqHfLjf
fiUg8MHvrJrFXr3AOuIpGtGoFq+RSyfCNCV5ywSvh9IeOGOvMWruIhxLOfhNxuya
RA193fe+MqGYECyxRt5WxPLx4EMiLEIi5bS+3jppwAtQ6875MipvPJ7bxb0toi09
solwetAS0NQFzJ0vrXuAcn5jl1mMdhy1+A04Xofeiq+gFnZCzzWKZ0WNgWxdmpmM
gCAFBlZpg7h/nv0WohRot9DvvWb6nsRjM6LnhGiw4tNrQu4nhCgB6myuKzrnenfX
TEOECYY1bc3kIPloS6RiK14Fs0i8H194LT0DGQJ/ojIc285yp4Ree3kKuvy+pQbN
N8UXkTaIwGJkGUdNPkmIHtTjR2yIreSOhLNL6fEh/JfSrZuhH56zWI6KA8vleTQp
xYdbkiCzQXA7yKir168tkcp1M+uotP9tiMbaPgQ54FD5X0qmQBezwpMGXFVNTsdk
77wW/cd0Ne/UMYWEsdSGIEN96AxP9L49VqiE51r4t+4WCTIhtTqKvl1/Ir5XoUfk
ns57Okma5OugEb8lMZHrQh5bnar1gyHR9h6g7WOsii6ZyomNSfT1x9gIlO8n96Rl
AVe0xRFsiF3HnTYTNCw4p6zhr8zOlaXeMDaSh0ohplBcw/XngrqrRU84PFblhjsw
2caRdoBEzqG8R9ighsIfnqn9vtymnL9pXk4HU7rXh6l2R8dCRzNXTi3fJ3I8EOtx
Se0L0NgA/tKla73KrfI6nqu4SqyaVlZDgJ+lUuM532NIUk2qDzSMdv7EdLevGfnt
Bqch3g136n3FriHcIUlKko+JmpFZMtDGnUW2IhgZcGpnB9vo/yx+oIYwMMTv0Q2Y
xDt1UZgP46v9JwzegRxvuAbhXYdKYT5tdZAPmTWf2jL+04pfolzZrGqAYZ7iCisn
f7VUV9764Dap4KmkUQGvpIh148GmGhQciMOl0k4vVsa0ZehaPAGL8JL37lxdHu9j
CLwCFi9zIdI2Xx8DHwm3v7IITO8B9Hg+LG4uM44StoK3g8uVfClUk2F5W0jrpsRk
TBc+8tJlKNKheQq0d4fNqD1fson0/3ohHtAfavu6ZoU+WAv+skcajWqFCFp+JG4G
NbcdUWg4VSL43i50ONQoQe1xlpQbNSZrqFR9o1CE7+7QfCr6IymNsl18lQcVBUAy
l1Lz5CSvXWxUN/hLpi4qCKIC4EDk/iK6OKJwsXsmrz16OlaZkkILEHED11EZXkzd
Wzk1eQBXrkicLLEapE859GMoolApkYq2HE5mvn2cgmp8wvyF0BHDcwur9kq5/VK6
rx1CfK+5mX66dATCail/vxLyxJVd/dKIYAfP0ICRyep9NGsrLWquhpLnF0NaHOJ0
KhyRMc/GrADObtCper4S1VfOTMku2fWfqSl4/ygAst/h2nm3Q4IAY9Z6kOl4V9es
YYIVxJapcToTGfKjjhWOSOSijpkaC0Bo+jGtS6TB0kWTABX9BkU2AqOsbRnGDHQs
nsq13PHyiy8panEcnvCrbV3HVuWS46MxvUE8f7F5ibxqNylP9Xers3vplMxRiowb
dRFDhzoE2Q0ixfB0gv/G86UaYXF4BBgKUYc3cn5HRnRpfBgN2JL/WbU2oDGprzXu
Yoek+ocXtsMD3kRkaOZbYVoKUPydRb6H6QXK6HFqlhW6NVDR5WLJTVFLpj9AwHXz
+/m043hU+ePrbYbM6teEDryO7BRcxiFMGIJeX+ABaT7UM/ZkcuOa7OrbORFv4OHt
0W0i5TSZ5RvudToaXw48TUlHpWtULeHqzOww7E/WWKIRtqg94TjTq6a1Jui3X3Po
iJcgMHrdkjgtyvSdIWRTI9xzNkVKPvpSYHI7DPyst4G44YkPDEo6yUvdYhDuXJxS
fk9gKfuV/D5bVYp7GuYBSXaAPO6eBYvCEZ2EogW4CTPIa0vf1nkx9yHB6E4+N11U
0UEfsstxf91J0Up2ZpCeXe5hyKv1tPvsO6ptMvFkhNTXuHT755z2fiJ75YqwVKfM
Y88Pof74vWRBFqiTlQwhKxb9LCFRaxubsPwbDOtVQaKUTKHe5ZooAM3G9xiKD+c1
0Nb8RI1Jb52ERht6UUq6bplrvUk53cbY9lGVztbJdnWDiEef19mAJHgRT/vQgvqe
Zn3Wd/ay1BSKc33E6OsQKVmLesrRCS6Avgwh9ryp9Z/tamKBeZtiOVcCb0an+1yQ
3Le2EcxhoAz3T+snrZ3Oo38vKygM4bQRQ/8VGMqmGoHcqfXmEUGpfDSuXEk4ilY/
LLymP00fxp/SP+aS7eQXIJ+y9MlaiqlOusKv94LhGx8kpqDnaYDGausM8cRKSf4X
hvStKmLDnz7xhQCzHOhyQdYqhJdH9rbdKaBB86Ywuyq1ibRWkvYJn2TjnoofuOJu
wpuSK17luAQFV847JYOBK5cGur14BLM3zW4VPoQRUM0jSQetKKCKtLrObU+UiKap
9nE5BLinCNVKXH1FpLd/NjvFxYDhOrXgbBY+CHMA6JGb7Ok7GrFphd8lFSB8HqH2
ZQuPwHxuU54DHAeDz4ATj8yknVCtpFuLRkDcN5pv3F9XvZpxUlhD52nSuzS9xoa/
8VYRHsuVfZpnQiJY/ODBsDv3FsUeFIcA3f3QU2gdQMnWaCA5RKaAtIUpK0TdurMt
aaQUD/XANooJDNCrY/veCQkXZ5vEJZp5EVIqkNAbGxae2gY6acxFI2S/pa2sMWmn
IFI19f0kvyRgI77lGL+cedS7Gune40MzLEsLXh47DySkxjwb7dcjG3dH9Yn8k9JY
tlNqapqsabmzeFt0WK+e06uNphMB3SI5iOMIqfQXgJivyv6O1JF2rkhsq/rPPgSA
DT2RMz9+p0wxnaO3v96K/xiuMDQXIsEaSqiU3s4I2ixyw4u8qvTIdTx1tLCfSqUY
LhODOExS9fIcxeYICfCcGEuXtkndeyoqFYSY1rGaKHG/TdcOgC1K1/Oj2VDMZVJK
yEh1nfwGtFGu2IpfZDa+8N4X66W7JUhcJufRBi/3XzO6XlfR4cA/hz+gspAi8VIP
ABmNqhh5MQLwEeF0zWxVGgatLCiyYrFSskUXdy5YwQuxrDmhfUfTJrnCp+dWQw/5
9w8SghcS5OgULzT+DC1fG7GAW7OmwQsZqFqIXZiB1a5am5Ey6QqWCUA0NpaDpgwn
G1wZ6C/MS1se0ItBfmlnF5OE9/I+5xGJJlQyGhTTPizQ4/K1B/c7ukMEG9iNxun5
LAGdgOQ8uKTgmuQqvL33uA2zD76M1OV/Q9fJofOP1CId3FZ1JfLxnNw79lLzzrJG
YhpwjNc2JOAKh81nu+gmxbNGZ3t6fskX2P6G1f0tFkeMBH75T1oqt2c/0HIeTi4q
ScEmj2+vo/IuazqfKd0faidjWXEVrTNZoFXAK7et782o1Mk/eo2txNq7mSiGWyKa
vBp7Ib+kcv67ZiKBX1aqE1afTwQvNFVGtHUlMSpjoV4fKTPiWWqzodWGoEmrtlPr
xy46cETMhuZCt4jOgNR8L7PAxiIWMC+4XxXnE8J+pRoblbB0lIiq+IdHxIBfF8sw
zlX4eYt4YcOpwnwidCPelzcW082hUjiCh+tymAqVDHSP0NaQbA8Yo2ljaqCd+zIZ
0T6qo+0kJuG7a+JgEBxOTK24ikE1/UEz68uD5PIB/gyrHh2Xw6YtZ8TDHLW7uCY8
S5D9FBmHXq2V2XFu8pR2G7B2JlHBdSmNp/XUAo9LIYnoWDb8LadrHvkuWOuAdrwc
Uh5oazrJyUlxry0ObUCbSfkWrwu/vw3yLU+AIDLoQG7sot+GeZd+w4Up6Dh0WJxI
/rxAVNHY99q9ECkySHOg943w3/AvuaCOxifhLSv/eWqnbCC5NLJIhWmtp6zRqpWh
r36snsj9ozq7b01EVLLowidmoxmL4cCyBJtC0KUIdbkvq8JoKWZm2iE/4S5JWUho
RbWqRJVVhyZsH9j/woX2YH+UvAxsZRSyxGMH/ju92hYJbEtoFL39zCTShTU/EO8h
9jis9S0qW+Lc70RT/+OogRUcBXYm0UZ8zyFxfAaKt/5ReoP3alT5/dpNr6OBlNIP
S19CZCBybuygmtoR7tcUlccwFqfA7fmH/ISQV6cb8tIPRjOvlL+dvVT8InealArr
0J2bwB1MgPsSJbf1AQNs1Yri815/IkfkusRZfNy2RYW2c6Lxlz6bucfu3v31aWy8
5jcJVKpjr5ooL7oMbHxZrysL0OhkmXcTprxh/66+Fw6GVqUHH6fNPoknrbWfXann
oMFZbmVYlRidGKofw1+6+QQgjw3MtAntBbxs4TEf/OQP7REHHUkn2qoHrI8NRWlT
3wzHzPIhYnyomOgwwpjkB74nKj/IiJu7qqs1XeqMG7HCXSE5xwjudAYa7nPT7lbi
mUJGcFfoP6je5YyOMj71PgDsS8P7RVfEXYhOZ/ur9ADPuTxjGf3J3mmXc57UxhLx
g4XdSO8+xLx65NR9mh90Qo571i5pPKsjL4dUD0WUKf3nFJZjbvg+7+E+Dmugl+kR
qr3O57xbW3WrHMP7gnpSAdH3lGpXoypavW8NB2YVpLfFXNp2lCF967fp5Do3tSJu
MVJCAQGeo+bKvGv5tFUT3oQkWvFQisG7y0xgjqyShM4qkvxTkbuPGHlSAcmoC4gr
UOg91sc6fc5WK9usHsn5y+eNxe/0mcHnlXmnYNnIH52ObAFQQl1BVCMo7tvuOA9t
aUTUu+WHuc6h6wb1AA5SkzxzCQ1UD/iCatoq+7FGkBTpnH4idIHhMBAGbI+f+rBn
BqBZYRpvdd5e1GpSKF3ca0CNrTuN/VdAz+QvcCExrlcwFA7gSQ4xJDAzuuTnJQgn
/kjxNqQpN9sxCftR7+hQk+2UIopDnBkaJuiO4JaAbNb9+0qbwaYH9yiOM8P2aKEU
UaNf3JvVy1UH+lZjhQfAU+s9mfHrOXctc9kAlh1GitAeirXh28Nuye+3XkVlkY+v
5W8veDI51kYY/gPljOv+jRy53h1a9pSY0y4pfpPm1PZufx/Us5+Bc6vECYmK98on
0YeDrZ43mchjwNaS97C/ZGHTtyiTYs1jhjIkBkn9AjT664c+ov1RnBNTcCOyb6v5
GnnXfScCoyi9GCepeB914P+KBj9agKYKodDDcafd4uplF5Ed9WJaDOoFYPxRA9vR
93DQ9DEQ6ZmgITIcam5D6WQU9o0QWjaF7+feT7PLRpEjcVv2fNr+6ktPp73/zfbv
7B7BXFufRxM6kj/lcT1eO2HpISO9xEHDkpfqvIgJvwGmoORLnLnJgTrc8x0ojr5A
r+WtqvotEPMJhw1UICpW5ClHWEvXYbc/KCReXMfZBhu1ZrPW1rs7I5GUKx0hQYdX
jcXVHBr+Aw+wUxQLos8sWBBsZp1QBD993L5hN0LPIhDnzJr99xYHR0qAj7OF4v9/
PRtTTVHrQzj8Uz7vzdN5IacXnfN+9jYm8TIw2TDmDf/Ggef34A+zSgKwp5vsexiq
sDboxfJiSEghqxmZ4yQfa+eFgTk5xm0jOiU4G/UW+lp030YKFSwC/mzHydlrYkbY
hm4OqH5Dg5Ie4s1yMmMamTI/EZZ7TK76d0Tif+c5CBVgbZLdJ627oJXo1WK7zr9E
QC2IW22u5oVMrii0vCrgySeycXDkK/RWchuZF82jyjzdh3MQSaxYDOfNYB5qYQ8I
ZxFidxYLqFNOyeKL4eQ3uhFrbV0TzjNPy4BNpZ9iMA1K+gG3F7D57DyPSWcVYEPl
zqy4HEVRiKKoWgfu2nUVVr/vknlUPHwHP/TOXPsUY39D+8kXuj03LylaXnN0l8PR
xwk8Gyax30+m6CX+lp0vIQyvn3LO+rluOUe5YI56RAjGrBP6Teo5Ajtt0fOyu29i
ghyKa8c6hLTTyJM8Hoj7kZa1zLxo0LuLfRKMkaG1Ab3LMi8CNln0KaTro5Ug/0yF
N9Ec+Clv6ParJraYYyt3XH0nZSKCJX3YHZMEmgeaGtCSN+P0XhBLUmrEizbxnkV+
zwikfVgOuVemUsen9OobUTyE+UJs7wQ4QsA4xSK6BXfp38G84Fl/3CA8cL93U3KO
crvAIRLXHtovFWJeRiuAiq5vEtsw1j7C91WoU9e4hcAWbwUav4SUlvVLW1zCXSnG
TDJSAF29kG94lmn6sUe/QotMYvxvaRldXJdRvdbh5ebk0nPjiW/hSCykP93gNhSd
IvFbAcqbP7xENWmWzPf1uqdBfuKdDm0sfNHeA415bT7cJ5H9H3V/YpVJoGl2mDh4
KUf782wT9XDiylunfACodDkY74PPuMz0kbNpPWm4Ks2DqH+Hr4i81mDQhMRsyppw
D4CHsSAgNp2JxjhyF2rmg5pjr3BqGZoh2VlmGIbxZuBBPeen8QHAvj69CRLQRVTj
yYYOLLeAiGq6zjYJi0Cnmv6uSyfVFcvYaUn9LCrNz18/kaIp4yAZRHCDXLB9vsCr
apVOTcgD/Pi7ZJra4UbhP8irX8BR8bLCm7iBXCim4AEeEzh4334pFsm1NPoZDaC8
AzD/JH/1cFmWkLOMpPhl/cE7nSxh/9scKp4ROjHh8BhTdqPCEYkFr2raMyQoNZkV
u3YSgaJ/uvCugolNXWupvhUXs1kQp/dhdHGjJECWCOIvnJCFDzjVtLWYD2pWV9re
aOR34v0HcsIxz0pKmuB1Ahj31rLHmmKhZGn0B/2WB8BWOq5oKC8eKHwh2fzFLAQE
csOSg5t+mSbkuRrPEACOngloMYHcXrhj3zpW4qczPcRHFzX0QBBi4D0fqeJDZPe6
ZyNRqRFVaoVDzWcRLYrWyAxj0R2hEx+XgV619GU9vov0PhtCSRQTkvZWLXQLPNAj
C7qQyK8YM4NoMb8Aqj22aRt3/xPh5kXRV/Oj5Wv9zxFUf5gfDcRXE57m67W7MRqW
/+5+3eyF1/G+D+4o4uRKruDK/Dy96vKXvOA16BYVwqY/3tdD2L6aRUHjE7Gq6ZZN
TdL52AsfQcXVtQA7dTytDv31G37bECS74bwZcczTnQs1maIUSj4KO3XNqE8GndvU
QKI5djR5TM7hhFRVlkb77EfIEGt5KU0tQL1KSP86SS2PwmAph31334uibIuXki5u
nZtYpfxTLmO2KMXUGCOk0Xr6cJyoDSVULtRdTdpxzzdvrmivg/ZZGFaePJfV/qiq
lcfuYIealRvj4JuQMiO5bPsGuccCjHKiY48nJ1/Qz6LTv2n0W+idjkqtAAlAkj7C
f8Oishgu9zBsxe7GCmKFU430CHdfF9wnnW/y9ayH67FVzrWNzb+JTSKM6yHc2vhQ
WadAMz+STji3v28i2MrjaeENI7rEsMI2ZH8s/jtfYJb8WV9zArYekzl9DwIC3+yV
0jmUe3Ik+dQdutyKL8D+oPyP9XSZzyitVyI9ZRav+JjNV1Lh4/EgLTQaDhtpxNvC
/a3RMetMLBy1kvLFeWY7T94UJXUMQf21p9DIwZjwx+kFMKwPtYsceWFyf/FWVVPF
RPtxVbAcU+gH4iizI+28SWJnULGw/qyQRRZ5/qf6Irc4zfSLchziYrUH/WDLilgK
9HesPtt18iDW3daiH6pE0udoJw7Vv/1N4kbTSr85qGEMeDb3jl/Hgkf+3Az2zwog
bRSS5imi00Axgtghw190o1L8C7+uUaR7S1pIXPXUoFG95Snbq4DuUI96rMn3EvaI
7VufjlK9ctcJlYJ/B7I/t0fFvzsSFWxLBfNpuSDiD5Pn1AdoLk2I7PxDUEwjadJy
OW1003fSpZM2oQatYBGMnZwap8SxyxjlyDRqo8Dqyg3/eMdEkchOwHlDiZk0TcnJ
wVhcN60sXDv8+X1HXnRhw29rFCzcYSSHJCckkkNGp47qOjN1a5GR2uZ8pbVBaQpx
pArTFdbS5lMzRFSnbRKgWJf4oBzp4sIeNLnJ2kdG7l8ziMYhVWObdxE6pZubZCNP
3s0p4KYtxv0/AhpXWN+esL+MJlfRjEgWnG3JEJhZrffIseY0YBLzK+EtUCD6gc9P
OB01GGH6jZq0ZPfN/g77F3kn4+2iRNscrPg5V5su0TrHk/GYAmoJ8dpKvklkYLDF
mSMpxQp5D3wWBL3pTe0hCJJ/gWWuzbK4FVjSqznBIXmEYByn8foNLBvAdafi+Q0R
uJtyBZppX5iqXVsuJhfiZaQ+OkZa/BBeCGuRigGNUKm9VL+pU4mZtcmqZqu0vN8P
RxdHo1VIemBsaeZ7hDxzPHieeHj83viXzvBV2IZaujVI1fCR7X9ACRv2nsHiCvLp
ek+oQGy7u/wv/WQvp/4mbIvUPOip74ryGAq8ZfepHaAGQ1iEtAe5YOy8g8MdH9uj
DwR2XktLGxvMuZyRXcRptTZk90uwoxYmLrPj96Bi/tgOmv/l8MFRBK9enR6W/AFs
6BQzcxyo0/CyKCkaCTskeRmGFeKdIegBlm8GN710l68GRhf9Lm319P76MLUDZMpU
Ik+4wWyV+gvOKzMA5EOwFOhM9xAa6QUvv3iMVZnD0DapjD92KQSlQoRRrKox1xrF
5xzCBIOqwIkDPHZDnZrqdKHz1G50f0I9mce0d66rIQ4+Imj9ZP0Z0zLvqdFKkiFY
7LYmNiPxFrQPaUNU5W3AX9b/LgENb2Blgqt9NseWH1sfhSjXyLflVLbKY04tugeQ
2rxZjvHf5O2DAGnqebHwbfrqD7skhC5yel1dxCHeBgPcOrVrXYPNNjmKwgWH8TJh
fUFeL7+f7qpfG71Cx/q9cdqQsX7SRBAMRHQGAEKHab3WoC3hwI2nD1Fk/l+yaPMD
+bYppcdErZHzCg54mRxJ+Ak4jYwsPfFb7uTWWHX73FXHDKdgWFIq6i73wRhmRTvk
2jfMb45P+SOklqad6YbpvCTMS4zYVX9HqIzC+hslwgSqKRkyo2nTwvB9B8Ul2hBS
jsdHT4l7bw/eQo7a4FyTpg/q/XWXE9vFKB8lPXvTzfVJxYQvJwhlA5k+ldajR6nP
/KjJjbeqVpCWubeqhsX8I0Ut7xlp64FZGBMwZdHuE1F4XGfVbfqmJPuy402hpqhs
jCnl/u/0qeMMiyT6v6zWjfUxYTguLOOqOWHU30IJ0GtphQZ2d8X3QneB4wuxyrvm
5dJRNAz4lOhAL2oHQ7uJ2amubu3by2kwlhUMaJbi1816k0cTLmbxsXdt4lfR5zZI
c2F7S6syEDpDqal7rN4exSJRi5RYikpGiCepyiC4SfucFMEAJpoAyxqTduJbbkWR
jCtbTEjBrOcPKhH5BUXqAP93aexIeHEyglclfE8bzMbHvpgQIGaPdX0Utai/qSz5
DLaQFefJZjPGo/lB8lku5LXUkofW1Ms17c8Dm0tpyrpedUanFCdHGAeP+ueJHtB+
BWSLFTL1XAPUlStmpdYEcyORoByARavekBAd/yOWRqT4x4ZkcBfyJYtF54pDJc1X
XhBRJPRwLRf8V2g5DZjw2rPvPiHNcvqVLLu/MUnPi01I4+ptiU/FwvmwXkaPhvRn
gsMcGrythpSVjJKpgr7b9/G7XBmlWfVhxTcgCAxBH+HvEcTsuNSRQPFuMYEuCxi4
BVbzA91IUNQW/1+oXaFT38rUNmbo29wd29nW2X/OYL+kIHzCHyvrvipyMSX2PzMY
DhPO5Ce1hobiUnLE9D/lQLb2zIotR9KLQTCjYqVF53aQUzM9tY++SX6B+DuPE6pu
GskpR48S8/lvs/3rbqPvj8J8Q0H90iTrZ0Mpt6qyzlB84EqEKOjNjDoR2N40EOsv
3NoujY1OZl6zlfxPjukSrCsyH6OVIaLAD2vCxy7r0eYTD7eYQu3oAGPK+FvwAb/4
i777HafPu5PTscLrR5Km85dCCmHdzkF5HI13etuZTJtsFZN3zngj3hqHm1v37lJK
Gj/ZqG58deklpxIAgTl9bDR9/qJm1wk8IbaKG2FkhbSGU3kGSZLIwxhn6Xw+nU1P
F4UVyTAuCeIqbW3s0xIvBDyvU0HmmRGEUIwlbMtVjuCahUetHLKmE4+SA0wi2Dsf
JmoADJ8xAnpaOR89GzHI8Eo+amQPJGty1tq4xew9rK+rWhppmcjTFgivgtuFOwZl
dZrBgm5qcy8Nq3Me5LlgjxCJ1Lg3pdm2HjA20/G2aMVPGe3p9twG+AIvu4qHKCCB
fe3Px+YE4Lb7A5ySWwZTyAB/P8XEjo/yRwbDx1YkMUj99sPSCquIPWnpAp0/zcuB
1OK6fBS2eUgh7AOfDj95go9xE0hTElJg+TVYmcWI5pagzhQCZFsLftiIWSRDR9xI
4WZQhdf5d7YbPdeTrCgGGT/JhfsvXswdXlc+MHIgHqO+wqpQhfLcv2bY1T7Q+yKM
1qm0A4gStvSBDCNUzmud8nNzFaCUTYHibO/+DBywZY0Bo7MSRhdi9OO/sbWa9FrA
B+GgQMUzYLyCRZUV64sV3vmf4nODd/ugVmkm6PkcXshPyAc7NEh9ZWI9aBBPfVEo
MD+vLkJmbjCegXGEQUeYoPdUP7pT+czYugAWjnnqvA/bUSq06EX70A3N7ZaTpPCq
gDWsJJCG/ZFFd4jM5L/X5nptgf4I6o9kLPlLhyPw8hNyyIgje/fQDK3izaBO7xlZ
K1fAG3SAvpAes0hNYySC9Ckg+ujm0DoVxtgwIymiI+SFxBhyRtPNsh6WqbnNhkdu
LaxDlECqMpPOhqD9El8GZK9suzAf44+AcvYZYB6DJKbQeDzfDUGIK1Lc+y5t+w59
QStwuwBNq7EE4oNOtd6KGlOGrXa7IEI6tGe+CQg1mAY8ZGJDi0jajUNqfDvqmmTy
g3+JsBC+oIJFBJlY340BTMRsC4lLZclORczEa20J4+tHQxCjC6fBbgr2Z415F4DY
IC993QsqlS5nKnXpazHd5mCJx2WI7iHfBmamxmCJ30TQLyvs0GUmoDfpWF4Wg4s7
IZdnofh6xGkqH1O5HtjStTaQa8Yr61IbxP10g4l2Vj0Y/syHDBIrgjB63yakzF3h
GHWjFs6ig39qtdhmQns4qcdsMjakrXf2QCpSmLUJJKXRMR6gEuuhKsqrUd36intq
jv4Wk+V5npn7lyHHfGt0jes2wsk3XyTxzF27HT5IM7pFZXpUe7NnREwCQZMUXa9V
XV826NHwsz2nXzGFPgBdFRstPOpmcithpEuB6yDd37nP+3jbH4stwYIG2DBLBT5s
lVcGOgTquP/6IXYJe9Z2ZNrGVTb9w1BJC7VTrZf1BHQyN7+43F6T4ELsqFFN67lp
Cctt+UAM3JurFaM4COyrwZQU0z6bn3hBwWAjxWTJ46FImZ/urSuFmqO+bjY0wH0h
W1TwUZjdr38lG4ehf0+rONmH+v6VoDVSorahPDjTatg1HIHSxmqfn1FCouHnxbkX
BdqPyU8164oRpVAqWraRS0NiMDvnn1yWsAXp3zwMu6IGtYWD678hud2PHW5/+CY6
dvDHn6iCtGQlZNfZ7PnLuxPPK2yrzIOwSzlksgL+0l8xo+XLAtRx2+XuMd00X0Bn
16rvfFbpbU/6MY4ej5+r1pSvr1DB8xrA2m9rQdR9tphj/NWN95rXydHyK1toeqhH
GX8PK3+VFEDB3OtJEck6W2lsTKwINXQOJm8o5Y2pzJNI2Hh0o7gKsVIT5wpj7lDg
dJMRb5QBbTQkhf1Lm/4YDeod8iXknSHUeN5fp6iBSVxp5N5yTo+fOAYAdhd8fKVl
lMXRSokPZwu/jjIkm+OCSqK1JJPjvVD04L82bphHbJ7ucIjzZ5X3yNExKtNSP6rc
svdkYIzoyv1oa4UzBMbu0qwgnBGv+o9BNIEk4lENU6o4YyRVtq/XwPm2VsOqoAH6
lTOpxEl3P2WL2q4bz4G5AjOaKZk7Q/1KBG37qyUOSh0SgqB/XCxIRLy5xyuDrPuM
xTozz37sNSnQZldo+J6nWEn7kYTgAK/E+eujkAPNSeUi2/tTcTCMLtAZDbcezVsA
sQJ0XCFxlOjkx2qCqw2Xi/5iWWMr/G2g1vEljuEXBOZvXW/UoF4oGdNk4NMy9OeF
aS6B7/qD4iTsM4H1KiVBrQBYjbLrnbq4RG8jBfxyMRx+xIDbwzxjgZO4SDpnf0QC
BWyNqMEkXqxgdwwxGOGHSo5uOxpqNuItqRydvdGICx0/xfO57XoSV9NAwPHWk7E7
Q32cK9svr0KVUhVC5plA0AcC6a+IgfR9XkCSNbH8BTx4Odz2m0oaoT9IzRo2Uwky
hhqniOqxqnIr+ngQ0gLSvVtQD7LeWSxWN7shTuQjwH462s6zKswJx/Ld7M72edF6
WkkdSNUSgyfdspxE72g9swmYEfgPtomi/1Hu4klrPcdTgFrd+IpKg2qDbrJ+YuyF
mrPkBKvRj4st2md9qCE7FJ6yI13gqfZ/pyJzonMfyawWeAsIMIR27PRZPqxMAMll
UjBQc/ewvu00Ht8HieP4lK/1Kfu/WhCyqsk1v62K+4m5MxEfDyKyZ6tlQXjmb25E
3+gD8H+oeYxZIxzOexvm36t3WFbi9r17WCrlyNR6qC1lwzB2pvdC1zD+z5SWnNHo
URRU4sPQYYbmMKFcI2+marjn4tg1woQOAsne6x4GxvpydFEXFlZtQTrc8t9FslDc
mn/GRy0G8ThdBCcjr/yov698QWoEEu7FZoXRjG9II4YzS9LOnZLlA5/WHsDZcWKV
nSf+egBv18XakQkDeJLdHh2wF2H36G8G1HdSB1zTySlHin7VBa7SOvDhnzDAmUNH
OfcUZ7DyP5D2Wmpa9Eg+KyLNH1OHrvGF2tP9TcJx3fJYygPWsrtyGwAHh8VyhRwE
oe7GeGtja+f0lyU7/STllWnvYIS2d8s5IJl5R8oq6iM8zvwydJxV4Dwr5HkRkOVH
bhTjmWkT22sjPLYB/DFmiUtlbVxMGqQ4O8KfOGyuXzHjJLQneg4J5nTrzAOE9D0I
M/di2iqgjIF7PTpGxUs+5sQzhKUpgwn+c6LatbAAOqy2xJwus7iCeiyHs1GnKX/E
+KZTAhHbg5s5xM2kqbw1T1oUZrjj6StCcpkbl/Po3VHnSYhQm/sNBbm7X8mg2EVx
LTaTl90a26aC++MdSu7ZNpb8vpUFom5OMpi7PyYI3j3Jq0x349X2bWXX5U9n5Jux
uSze2v16eQvodJiaqSUFpNfDZBcVTBsGTSYnUHozbgpp3ekEiPdrZNNXArIQvTIn
w6fpHNJOswoCSPOMQk1MsH3MluaLHZ4PhzfbqIsI1Cu3KMms4dsF3F/9O4KLB6zb
JiDLC76wwM4mtNEqKL2X+m3gQmmRqI6XihzXCloPqE774gqA7DOB+5J0xTLMgHam
QgtkNaL7jsxFdfb/UVOxN0G0g7OSZW93qiLpxsxnwqLXlggPJ7m5/AAQigurS9Cy
EkopTvmfKwdJxTBf5j7bY80Go0Npa14+qjaYWqwinKUpGokrW7N9XqXScaGpyokI
pKvU0aM4HSKvZxKNMLPiZ0ysO7YKIXr4By4Rh7RMQohMXFwAbsh4AeKbjS9/Q6Bi
sDML/8oQvUGQebAKlJBzP21mynVf15QjsuEFip/Oa7EJ2vs6V0rScZOR42RMfjgq
tp+FiIvgiPRs2YG23YThXeyZ3SKmArM0ShYAZVR/w8dF75EHG/YjNbHfJunzs6/Z
qufmzVRoRRy+ISTjd6xQA1d84GjFRW+Dxug/QS/ETwhpFcbZzxvbY1cbvQWgcSdZ
9qUYACUqkOb1qRkesKV9BgrrhRNom+ZEFmDMnP0k+tLlU+0Faw0YamP5qencFOKR
vd/3MSabuE1DgE/uCKUGdBqjnWDS0nfbj/gfgNDWT38SNzSjnU9/ooumy4xpYGWu
3BHL2u3/p59DcwRUiw8VemtEUuuwYUlrZIIXbsUA66Qf22nxuF7XBXISXGxHA0Ws
dccbae5QNszmMRQ3dYBdRAzYX63ilcP04T1tCQvc88+zmdILcQt+DtT/LE6tg9ms
aIAZGbPtgdqAgSOUrpnqKEEkwBcc+vP/gwP0Z7HOgIc71Ns9ySoB0TBj95H/56VL
hxhH58J/hMAYwpnEtoazAqwU1BfjE+S3UeK/37iGTIPwoV7na9DmSJNtg6Ws5/hb
EC7Oyzio0b3Qp+E7HUnHVNkTERUFs1XcRLWpFpbcXiOmdGAQ+nxD1NTqTRENIkE/
BpPRlmfplIgqttd4s/INEjKXzj/3bSYZQLpNMoMqWC9CLLBMlpVLRjLNbbibsNbC
fgXoDOjRscP77Eb8RTao054LQilmP67Bj/SE1JFEJoFEG7EEKVE3p+vhmguocFKy
qO2LKY5cvslWOqJ5Txcp/Y89TalTvSUavvgs2HbNT26fmjBMEhRJTmkfL+UYeG18
2MQutQ3gw/U3zX7e5EHiDyf5PFeTotSVKu8Ragf+pDEjM5hXUXncNCaRd03hzTIn
DDy2/anDAC+9tXDJB5sp15BW2XOz+69B/s5CQkjje96TBAr/044V/WpSSbxILGz0
a5HVCKqmcnAKvd5zU2G3Yc5/cOalKit89ONFupaJ36cTNAqFu60SJgliO+dMWy+3
lSeaxzbDs3HBQ2Vjs1EAbHnD9FYNSK9GJHeSWWBp4bfbXTOis9i8Asv7V6Mwc4Pl
/Ly85/V/z5QaRwaTcd3V2ozBouwwg2pk++Lm6lvqz5QViQsvHG3v3iETOyyIuNDY
46CxgKJxzNFu6hxmIXaY3ffevM6diY7frbz7eRHbW19TwfByNQm2NKU6IoqLrlzs
u5NZkL4HRnu1GWElSzM5GSX5V5gzperHZ2z6z1uso+i60EXgpy8F287kUg0m67rW
l0WEa+Oc31lYY83+f0dqUOgTeciQcKKGAHjnqO2sD33j+V3vfCm/JUtFVNkBKwgp
sXxHtwh0vTV+S9gFO+ieTXiGCrDZQpHEn2NGy8dagSBsC3ZBy72/WRzWobjBqc+K
FbLiW0L52/whnSXiThR4Mv3JsgOgNBLUFPNUk71NMXQIMAlBprlqrd9UCcSH+7au
qhemUxZYw/nHSSmAXgCQ4HArllPouL9svQxEJB+jUM3j7RsB+UWb3jLPDLN5zfjN
w+Gq/htl+6pSde8F/FkhwiALn1xOQkfXMeRQXojCzF9TFWFgvvYpliyWJ9+fq+9P
pwP9CH5enczq4sREVlBj8M8ug0kn44o4XeP1nZFWrxn+TLpGDbjxkttcZzFBnsMN
LnrRX6btDoNjLgxY8zygBo9VYZ75XMoHIi35ksjhIlj497Jv08/4eXEOK/JSNLrz
VzHjv/IAb0qZ+sptgFvxOBuKjT+MIvETWmgoQ6mCGmbTNPa5Kk9cWcBv1CRj6cVp
hfEhiI9BoR4Vmfclmakxr42XTj7qC/IjubBzuPH797lGrTyYIiiEXlGsg2b8SxHi
kb/T6hOtL07dNHDIYaGV2S6vtqzcZQBkT3SGRawaUiCNubcSiPtFTXGEu0UOJDGm
SuHo0mvrhs5/iBocrq4cRPm5Ol+fV9QL54W9JQQH0dvxKEuibjCULovXVtTMPEJW
EiodDqbPXpmd4/T2OW6oncRdWuPMOOMx7H8dmTUWqLB9HGvso1raT92vkt60cM0K
CEoXDEdgGtATL6Bl3WZvMD+47zR3coPq5SSqiPaaUBTtcUSjsSj8eRikhB/aSyf1
0RPVjna+xLd5Wb2SYZwDMOXjgR40HNq1MhnU/L9AcrJSwYID2QtAqOyB1GdBouTA
AOA8yuTAj6dTSjMgOVK1NoHDMglBebUVfcduon6tnkd54ua2zi/9b4+zEx7lDl7v
Q7361MVaJTLqcxW9ByMAbsvkEhzbe10SsD7Nu/olHu6MgrccE3huc1gKEYugPTkf
ymHVr+61wmaNYHR4mIaDc6Fm1AS0sMDMN9iQ9N/b6QJDn3B0VnEZ5EXGsLYXrCG/
jRmq/bHSnaREcGToQ3h1TFdW35zilDTaYl77cN25TQnXsjN6WFIUV2T9tGhn+/39
u6G1J210RR/5nQ7w+349jT3/f001PbnMZTjRSG9VmUbRmwJFLkftmKa8pC8AqHuL
wFugi1VuYNQKBKz+YRFpVLWDl6oD+FiEV9mH5R6RihNO1cc08brbL4q90DETkR+1
FxrsvcXs5hogkokgH8pG2EpiVmP7Q+2G1vRZ3MfNsFqrtLolLUsJb2s7q9jgo8TD
YRJJVrC9OBYcZhGJLxwSoeERjKUPOUi7SzcILIOBY6q6AAw+9Zd4sNzx9pJyBDY+
qRmxuebM4PZ42smAzxTvYgFNo+jCMiox2SpZ9rt0azcYd5qI3Xuf7r8vBI8pFjVT
FKIFe/WLDwX+b0CSCowmi5mOKbUwtGlnQjDvjEdVJrZFjGKkFhvVqqFZZP//PtNH
EF1i8PAFaTbMo8ky9vd7Do8TmqfmXS+Qbb/uRMkDlr4as/7Kn3A2mlPRF8iPysBp
mF0s49iIOWr+stbBjJXpnCx9WjHkNDyBGUV9s9EG9Kiw909AaQmBTHn+BulOBbpo
mHGPwIEytnTOZBJw6jEn6KpFFMT7CLdOci81+XIIiNZ2lXMRcAr1KovINGdz1LB2
FY3hvLd4l9fnm6F2PT6OsxPyKLIrdmGH1usv8/eQaMXjCsLcO9G8tyBVPbmjKigo
j9Ki0hpsKKIRc8CHaM8jSvP/E3N2ziAO57D35aU28ankFzAT6fe3Bz9KKnGGyiSc
/R0FyLDxCjQXvMFn5LmAifXsTG3eWFLhdZr29UBlXJIRXg9sX0IjqgJCNxFVX2lJ
Wpc4hYxjmZD8Acl8xdcwPHYG9uwp3OAoiwExScY8kRa6w401CgH94fBmzmt9s9J2
KTvOs3k91RcFYgcZdJeHEaLyNRajAWI6o05rBrJ+hnE3LvZQpG82bPELd8jnit7C
gcN60nJ72U6strwsVvvBtFNltejfyGHXpcNYxVE1lBAvGaKguarYL2kfuSYryZtc
VYNMLCa0hzEb0G3vXTuzdHV1F5qRpOW+hgCYPrBOG+8ILD7veGui5JBjFPAkyW+a
dQE4DMW/HHylYDJzImI/V5rqnV3hIWECZdi6xoS9FIXUaJHEJIRVfhsRQZV2imZW
8bkxBGy5pDQMmvJXKJeNj0cyInQP3PvOyXU9iGIrVBseIa1nxnxN1+YjabN8ufDV
ll8o44OfXpJPjQj/ma1OFW+AORJtJw0+NqTZeIJnGdamIFcwcR0ISi/08UF+gu/p
+zLSUHoNfxlUa7vKVpzabKKVIyMA+rV17egfnNkPSVRvCEuL0jY8QgynQq18mCYp
g9+iaOvBs8PaRxNT+SRJ+lgkm8GieXgVKve62FE5/6sVc7Yw0PwQnw6yMDbGqAMY
nKUevZdp+fG/fwgem6Nf2rLrXuLz/Z/rW9s+WEcQG1c/l/6ozf+83Gh/mVI4D+7P
0KZeHQIxByLWFEp3Eu2eBZQAVJbQhBEyvSdWpfg4dkGe66Te+Qupo+DBd/ofODfh
U/Z1K29U0ABpaBvmbVRUIazOhHHwY6rVNwrsgSWVuONsDw9Z2BOR9wS+4VJ8wVke
XIqRT8p9Q4q+8dDaD89jgc8lR9ItZUN9HzKdYpc/yZ4d8WQKveB8A4znapjUTIX+
LeA0Znbd1ElLc1tGpdQhsW2MJRo5pHGcDIMSe8tNYIuixMfh713bGW6Q7pJEaygh
+jDKOg3KCNhG7milHrDE+Bpz7Sngq+9oLwIK+2VTob212cP6bIK5h7qtZTZxqz8T
DI7Mfl8RvIbJGI+zDV+I9Bj5w1LWsjFIgai0ME0NDIc+4pyaXEWuQmsnZUERGon3
3M1IhlVyNmnGuGd/MW8FIjSrqd1Uc3L6QUwSYvOlXm7MoBa3PM8HGmGTqkZIaV9H
G/cEG9twWyqgGFJ7zL54iqenhydqQHyq1oddhPNY+8+Sn7qetEliIYBYja471XoD
zQoWYfP4WfFzuTlFEy3XYuHvoYbTI9rGSO9NOyuWecVdWNiX/lKkIP5wdeTbQFvE
vDJYuxCR52n+PozXTaY580ruMXnDEACrXVynQiKTZ5Aic0tfk2dDeMY2BJo1L/Ft
xzhgQx6HPh1z5YYaSH/1grG3VDTpdLZOx2KvL0wmeT1AT2Guy8SnTL5IbBwcdH+Q
c2/IzPpwlm2fEA8ySyzdnryFjl4cz8of12GR/buQguv4Qz33zpCdupCzbPj/SSF7
ZvZ1XnF4M7/0QJDOGqMHVV1NcFFF3NzwPvnSR2q4azr0s1y/Ofr+s3N90WzcrMn2
bUOIBAzSzYUKvH0AFkiuhXNXINYWyUDF7WNX+Y+NqWeqzt4UdRthgFev/TMIaGoZ
DEmy6D3bB2auJnrpxLfzzdmH381MuYog518iTzlJ/RCxFs785XmcYdQCZ0w8LfTr
n2U3JSj1wRGmTKs1cRTYM3lpC7FWxhAGtuvv1m436RhFw6lEVbTWTv5/DYvVc8WW
PVC1w9Zvx7HJzGRYsac1GUDuYYIrcZU8ivuk3jucBjlXc3WbtYSyY8iJJmu0Hxpt
yYw+cO7ZAyOqmNqjH3QZ1y4Chwj+OBpyYYbmu+iKEk9vXLD421tQpf1sBNhPkf2m
x5oGxOd2ugVjGOh93oxUM7LyJtrdBaRNfJ1CnQbEx51yHmPLj+hAPhznK6ep1gBF
kQhQoxKSmPWeCV2UtWYu2WRccbGaUuCr4ByKeLqqecvan5gUsdYgMVp3ANoIw4if
6Qnp6FlFjSrq/FCRgGZ93GzPLsWkSaL1ekdRw365sJ8V+bvRrVLyu0oQR1bSdRXy
6XrhNkhuIoJQhRHWwsisrtSbgZuf2b3HDKMbItyMjGEaYkxaPQiqd11qKIXvjyF7
vpRf+4sM14VLwazUCL71hRhEI9tcbGqUC+WCJOBt2+ge9YW7tR2JIaqdHhB5Hnw8
RyRfLV/Z7T2UwjjeTVU+B+n4xJffWQq5rsikZUtWqUSPjjuAQHkJhYHXvJaoVXiG
lnyvqLls4B/qqVB6fn0Sjrm26yj/jK4AIdGH5zBF/1q+Xo4HnwuzZbqfxqWA7nxr
fUunaSmK4f668m5fJ5P4v/thTofdd2PxI/2l2RV9vChXRppzNP7MHKLrxHgqKf6o
5ewiDGsWQSNl/a7tOwjTfZf5ouTqOISzUIiQ5DvJEgGjg2ZHobnA+CeulPC5uZpL
jpGfPW/Jt7uegI992/aHGq5BmLjdFvOdvWbrrIEzUyBFiUpfzw/LTqso4TwiV2c4
BSxHiwuHjK/w5DSeGocEeSSSdTyYUxyyP38XCuWbSNnl28zRpLzffpcg0dfM0CBR
xJ0s5R3qdrdaTcdGKas7Zk1i8VU57xhopAS8oBNVX+oIHh0aw1HLlUkXBchwMejf
UtwV4S/tPYwCmsrzHCXruZLa5PJZDw/meUBc/ReSOP7Qg9EAoSnIeNNSuySwOzga
WUMFO6MI6tFFD8sSZXClWag3KFE0UmpMvxQjYgQNiQKHRipx9b/1b22ttBpvPRik
6fEIzNIzdxFRRU6w81zUYPCYcKtithbqQOUdc93Sy7c+UZKtyUVkKTkrWIBzqivo
I5CnYtIekTJFZ/KE5k0FMKxM1ExT9EZcIpB/aMRwYp9hz2c8losJAEI4CAVNjFFI
0rx0wrruyqg2bpUbThpbGXlYSBdMQiIbTleQCjnnzDGddNBb4GwYtBZfs1MSQ1zh
ZcIsQixBYkIPqIEG5eI6/nP13CXIJWWnJQp5JwFwTPKGjiNt1ibg5hayAAA3u6sT
9vqEBkGevztm3fhO2O4bKynFrbKiewlWyJ2MkZjvdCOcv/lztHWyvo9J8yBjIu/K
fBNjRp93HjfavaFTJu/kj1hh5IeqBGotNqJBHL7yzVdLz6flzlQFtYrTzPrH4+on
0B39qwSulonFk6+29YFEJH/nNv95dcRgpPG4Vy/kJDVquwEBf7mvF68zBbp2xAzo
Ig0W22lvp2aGCiyGPUwp1MpgPrz7cQ7isckmYJrgTSFi9Rw1CJknpaTuwE7a/mwK
xLH/IfEcEM5dOEZYKbVEWqDl697ZmtvreN8FLauNZg/wQex1QEnqEO2Rs++lfAWA
+SpxuTZjGixp9o9RYuJ8WJfSmglJui1xGNdinL/FjbF2p3iYwp2ks3U7W2X3rKMa
sXbHCfUYJ/A3RNfqV2ASoetqyFh1O956kA9SQeOuoRZW5NALO20bVG1KdVu6rzwL
wyQP4weq0/Q8i66/Dr62Bq8UiF7Bwb0BeT1t0J37vY7B9rnM3p6QfcnHT7+IoAtI
gwyd4ewGa5i3ADk/sBwHzAJjKO5MB/28n2l8X/W0zCkaXx6QKFZqJOBdtU+QBlde
8CZJKM9qm7ZT3ZucIwq07z3Lc5GnHN7EGYFgJv0FwDptOVUa8zB0Z2J4g9amptwS
AicD4+Jv5aFXugfbmVQPDZTjaGNpU42EpCF6+WAp9QblXltFUOhOoEEp9KmdbL2a
dZxqQHwYnBTzSQPinEhR3lk4N9ZdlaAGWpV1dsnBiWJ9g9gaQNx5x0w4TK1dzjET
WqwECPy5qXlciTs6H1P7pyvba4tHuV7KJ94U8AfYajUSl4AsN0kZ6OhqMQBbFgd7
18xlpqILmXuBilQFlP+ExShnxg+nucMTpZGSHB3CllzOe0N374v801Wv/4Ktt46F
eb6AK1WmUpu01yvbIUrK8RSO6DYqAjiE1c9zqWCdQTVvyT9IwcWndzsrDrobRikF
U++h15+gTfeHljCe3c9WAtvaMh335PiOIHXveI0Q5hWP8vx6gx6pjCR47LTunPXW
5EUiQgACdm9A2UpO0TMiM3rYymk/nNI+8RkFtzTJ/hmWSU0XGJ3Om+y4wZSNJbr5
hSVivloqKgX7AMqiYqUd0qOe7VbgayiY+4KhJUkPwIYaBFDL1tTIpu8BlRm5ubsZ
Skl2RxLVH7U8eQDDRMHMnEeTW8D42DWZIHLnJVr7Ll7bHz037flmBEh31UqW3wZy
u6X68lEEK5XAdVKjrwjGcLa1QTahbV/KMTimRsOe9W7zfuBWktzadZ3oZAZaP2QG
MMHHzznrfFXAdWEtFG65CuSLkBKmhEFurfY9q3bjx7i3/E6gJE8JvScK8sMCSAIT
tQILmI+3nA7I2Gr9b0zF66JMHMkdMSg+K5hor8EOL/yjk+p8f08B3g/zLgnUS25I
sRHP+XAaFUJ1ch6f01cOS2TSkFpAlpal17OHSxGNwzk7kuJPmU6BdMayDwOr/UUD
WApNI3UwH+ugSNmWBkv15TZ7zvRG7xF7t+ukZzOYTYFQ1jertpVttCDQE1JhPIl8
VwPfDsfvLucxYl9Nlxt3KCzSdGpJwKo80NHRMMVApqjPmdCjYUdCOxpNm0hp2OhE
ekqtWASPhiL8w5+3K6LrK6YLrb72knQuvI8AgtY+EDquBxQV0TMzHwewZUxw1Ytv
qM9FMb8CYkMghp/sjZn/1qGQmQDHKht39GfMIjDIb6XSuK8taXlYuA1PSuFVk1/D
vNp1daR9+gUIzioYSp4yOpdjv6ZieVnmAn2xDsa1zm89YJew8+V+u11IJXZT4Age
s+u8nPAxoPlKLvLLFfFJsYPRbkp6qf5QgLgeAX1D9lhVLst2IlEAgCG+rJBoHXUW
DJ9bhSkVfPyGB/2d9dH0gKoRxzqj/on1N2GCfGWgcXVUt9zbb+9V+E5QCYtMiN54
Dx+8+XfPWzEneWmwhD5CycfppWl0lt1GSfSwCo8QdGmHfYBDrqo6AdltVd9MDkm1
znikoCgOd64R3bpf9aGfCX7mzt7IZ7ADehrOEKDi9Kvaw0bW561Ddx39Oqj6Uvbt
M3J2WwGHJ5DY3Wug4aD14LewEoAzv/XjtCelhTrSAJBEnqJZ+2GijTX83FEqc6MS
KM4ghPEzl9SzFal2aGJFSe1+mZ+zAu+PFYChlMO7Vn+/v8fUIjc7LsCc7gfCVLEd
3JkloyY7Kno0ydTDFVoA5wVZq4X3PJ5hwpKoD/P/pcolhm+f96zAIQz5lh4zzkYc
ppRzErJ1qwzNZEStzt+5kMw6BgsinNKCbypJTcf2VrISB6ZoPewrFMtStCiriN8n
PGUk0pjBujavlV3gj6wqwm/ueJELFxCBSr9wmOgC41FUIt73mlh7heQ2X17/02nJ
9rCZRtuxYKD/kNmBd5RcB7lzp7esDvN+fj/Z/1PDc94gZBhd20l87NyN9FTrGJH0
VaaLz+35T64luvlPDaAtIxXDwKuPsr5jMzJj6FuKxubhqIyj/0YSUWkyiRXUUlC7
do5jFHCZatGMBKwQlyIQO+JkVMf4ckZsVo7n3zYmRA26INjQLKacDlLrAnElLezJ
B6HmsNpFz5gbDZxH4Z4EnP0q/WAuNrQhc9U0mdt1VRkpyBzjDXcVWXGGA0G1l9JY
LjaAyN0bJyxQcZblz6827713Ng5Vo1tjUKgzJw1jjZIPBr13sNq31UbyB/rWw8gy
mAJtrZlEXwZYs/NH4cnkLR+PDpO3L6UMGelcsFgK0H6diO536aHZIbkhdhK3Lw9v
nbMR1NuvyOivK8teEo2CXvK3VnAQD+YAgotYCHl94hCsMxDbGuFzmyoq4NdffXIs
NJsm8P8y9fbI9OkOGx911YXoY2QIW/tMy+IGD+nPE7Pr9BgfkJ4xjBIOP5tCi3K4
GMu2K1W99YuDPfD53gZNZeDl448GhUfpVBgZtzD4XqMb/IwHAqF0XJd/CXHwSRLc
+hdJyq2OK39+Qw2EFyjrc6GyaK7fRRH+r+cvaa8x74Xb881TX5MtGjNIu6iAQzIi
J6hxGGJgaKsU5+666pTQFJ4OXE0lfxti0Ma7XsSgvEAqJpbvfIdvA6FzUC6qTPVw
rb3KQcCBSE3sGU/zlyfl4jATAgOcdcp5a28iWvvsZ8+pqrpvt1tIIsfIdls+TjJB
CZsUHcRjqeYKXp0cmRYBHiQhJNVA80FLIH19VyFQyHx1CjK6d6BWCpNwCSz/1xb8
dNFTrcbzkqg8fWMxVvv6I2xHYzBvD0UYT2/2LK1Z4QV92FpL/QbjR73QrUlMJUkq
379kFqDgyV+AqU7IIY/S3/qGTsokaq7Z8VEAYkfaYaU1DRAtmrRPuyAB2eH6Deca
XNkh+e5c22i6PmJuwJGngv7vqFefcbP+Xz7lKKYNGOONTJaq+4ias7wMZkmGXaKR
pJZgfh2B7fAxhn45Vxann8Wqf5izHFM2mU27MrEjMc9kDM3xpC7lpKf/Sfp6Q3Kc
pymTMNs60lxwhAp7zh7jrN0aE088i/CtLAwqrCgsSzGnx8TD2VhVCLcPwMEPz8MT
3S0cY7rSCWqNEhpZQrVjMcK3kok7dd20TmPFK8CEJbJ/3PIhWztVJpJbBUHtFYK5
4rY8L8HvCzivrYquuzYcOH6dWmlUyqveB3YMzxEZIziYfhoTQLvUdKKAh6wNIXBm
I/EW5DyXktrGsLxms6nC+te1BVVtIccqTNtOrcSNRGM3rTYTMSPojhk4HRSzG9sa
ZHFfaWfQcS3Lh2Oz+tqaI2cpNmwZyY/U2U1nr97jZRwBm6aVoFsZlp45tXMmADqf
3wTXCqtfzfEUecibfWg4Ck5WA7SkXm3nvBcx5iAIuaZAVUybLBicxw2bNBb3CQIz
UU9YVqf+jLMUBIjO9GugKpqYjEDXhq5qEmmymYHfBX30peqoE4dJb8f+MQlGvNi5
PpK7IRbqv6NqewbYOCUU3cSCjkUuB0Ft/UuWshH7JMgBkysUtJr7pvXVxu6ipb+8
NU+wNSslHBp/jU58WGiT6YE0ksn04pVkjt62CjWL3H9SVzFZgDeVCyWRgvdVcTE8
PCdBGBNpsd0gkGGPgbPvO5tCdB1JGxht8/2s4GFX+gS10dCRQoCALloIGbb78mzL
SsIPJBOg4+ADfkUiN+GuCu+jIWevM12i0CNjp57Irmg3D+uZm87BbVy4L1G+FsNw
bILPl5RXb0DxkEuIzLWOi4X/9ZbeGGzJbYWUtM1n416qlYT9xoDivoG1XPbwxQt3
XyTH4Gr3QKpimiqpGKj/3AbEk2w8OLsgjo46z6GbCIN8MkQagPcagvMnpt2DBU1O
xUu0Mzlg2IBcWE/+QgJT+Puu1HJJjXRG3Ztc192xi1yuc1WD0MvMGaLSzV0uxvcv
YoXxc6grNevaWeTrD7hYbdDhVAezPkf9zy6AoY7vBMX7eEWSKaJFIKjUxvaHNpdC
ziXMSRpDzvx7ZyixgcuZ9dgRkDrDt2mCeT1w6A5MKXdg/9OqsP495BrXZCLinh2I
97cjXnteHmKF3l6BZhGu6ZpAMuS15Z8iMVhC3iw8ft3pU7KXEzMwcxH7RaBZTOsc
Vo7BdE3xQ3MuktrALhRaUwFuO9Tyyh5gq6ZPyfixm6l26cEaf+ELsVg7yFft2ljQ
Gr33F/VoODb/4ipBJS2+gJnbWhz0wjJ7/lq4tmz4OsrWdteI2WSsTy1FFMOSrrU5
AjH07mtSv+jZmoiJ8PJbCM2do0WioE6IxJSPjERqTwxEu3Z95UAcdehY2SvglAT+
qkgw5ofNHYePafQ4UbxfoD/2Uxhcdyb5B8dOZ1tHIb+CkmXppPulsm+JjxqlO+o0
n+w6Sm5NxHaDfBbDCqVrQU04hjFrJ0pvIqeUwDV+CzjTRy9y9fHcgZXgeVvZEZzN
KMpe7XtWtMWnsd0vXCotmlJqks0GefC3bDGq9Lj6J2aLcg+cK2QkKpxsR1udv7fK
F4cS2qhO0oyqT1OuoZ9RsIcBUJvYdnK99tS6Z7j1UjotK3MofC+h5CGn1H+RI0cs
FWyaE/Yl3Q0mgElAe3I8Z+pxdvGB4rAgnTPlQg2V7kJY/TLsnoncaaIGj3ZFXUmv
hY6SiYvadK5icrHs63W1x+A6N5DkKLtLrV5x3vT3vLfm3MbNt4TCrErw2mEQ16W1
9dxGpUkKMD0qfk3x3bpQRRvWmaJfqTPuzq47KXyq1B4MXVJkjyNHK5wXkDkevVwo
uZz9d/RxXmXEmaHUE8vVFL6WSUW1XTgbFMjnzUaSv9g/gIGnw0RV00sMfYqJ2h7k
dpy6fKHMsszHEAbtl0KYsJSUR2aoe1UuGijPB/TnEJtcI4xkLlO41eNG+U+UjgTY
y6kyv+EOZLP9tNm5V+3enwZuqBRqowidOMCmGbEOZ+uGGk7EnvyEuSijhRSHXgQ2
7QbTzh7i1GWxdmDjEyuiDM2zkZtmAjke6PPuCZCazzDoMa5fLNe+loMdjy35Vjn/
o7uqPrPqjL5egdjh7MvvrtOh3nvBmVykb/JaNCDQhBwbiBFd7Xh8eZOHTZDhfa/u
CUB6NEJZkD3Ex9qgtUlVyHK/hX94RjwKXThZ8PwupDIRgc8nw/SWMY6n7a2W1puU
KrRYPYIEVu4oWhWZ4FhJEw/osMgmxOnMjExdrR69tnNcQScZ0uGDxvRSf0jxZw9D
aAhlfLJIygZLH0RCkLDyL+leo+wqYoJfgBsb1e7Dctf2bRuo0nWDrhuuA8lUAtVO
3Mv7+hWV69grkHsCHh6y0IyZH19uLbCTC1edRhYVqnRO65GRd2ar6VLF+nZwCnW/
eX/eroA2dhynwXVF97WV2VtlhTDf+H3GMtc75P1k0vpnlt0RMM5Ts/DQk844an5C
jzFwCGm5CWDxxY+3wVdygF9MhlSRcoV81eHlVhtc9xY5NWfDHV5eZb+xuKke+xnd
Dyq6TkfDuxUwbp3O5OacjkItUqNHZgRAnWucurkaAHI3VEUpsHBQgjDu9cxWCeqJ
2fLWwgXw0igla5pLFhh9V7VGQPdvP98BKMxCQlllpl1t80rLzBXtPzhJ1A3tjSjT
63gqv+6I89WQVMHUm2sFv2uT1v6qxmQtpXOctjnevo+xYtulyQTMn8Y9EgKPJqic
gZAwSZEzgIO0e+FuGDavxf57i1YbLuKrcJEmCBwWAUXP9uG5NLVyv6T04750bP80
ZxLWG0xpmVjvOimtJrwysdOmuc3wfDtHCEQYRjinhAMwCIip3f688KSUg2/pE5cD
2boVjaaqPUe9ygEshn/1qkIRtb7sQU7QVw+W4HOlYx080NZClWv5gzrcis0S/2sm
gsmEiFpagxku9FwliFjdM98aPYm/8JJin9FlEiwkNzgKe10tcJzW60AFNuPwf7Cs
xaNGBZPj/F/ez6wRmbNwHMi5sWaNQ1ylnUQGhlYQauKW3zXdC0kx1e/vX4pbXcSG
zPods6cxkYt8P7HxMKhgeCUddqAZmaIzRDF5TmA+Q8rMJYEENf3J37cBU9NZNXKJ
0URowShlFT+mp25KYUPsTMd1iE3WExZuZaUwEKmTYzhKcdCpKpH7MNDma/KO9BHo
e3YElkCDLPLh2ybkPMVgb68+fwAKVChOys6ahdlZFZspBTN+p9ORRECwKeQu/9yg
UXWFBBlwP3wCUohW38fpxSOWqx3lLjK2Hz40+zHQkeb3oXueeQ5P0Q6bjN6EycDc
5oK9vd1+fABFfwArBMUQdRKvjXlsRLYqvTMOZit+Lqw55BOw6FBuT3pyzo3syFfp
T7yZoFW0ta1edXQFVjW0Vnh4zbsBrWFMvI4cOEhTAhzAhRMKkXRLmUOI9ybl9EHU
yTwfe+skGc/MGJymQO6RtXpAjjLClnhF6aHWe5X56Whf86khQTaPx5EJtEol2w3X
3z8Di1q9I7JlvKWuj9g8KFkDpL+8tw5dczuWeS8Ffk0x7Dm6OdqTVWIYUakMRiuY
KArlZXB8hbRjP23RJnCGgh6uG56IPAvWEHEJkor1AM3YZzdjmGNLdjUQ7SH7EXSb
i7RIDTVB6DRVE6H3AGnfFBgF8vv1DHhqUJ/Kf8v3g3DD1cYt6tg55R4Ev3SYIgCl
60o931kV8Ffc9X+YFZ2Oflkc0HZ0zq+Ubmrsq3AylH/lcvELCfbcFCTYM8s19k19
Q1sTdZMEVk4JXNVZ6R+f7z2no+3uyvlviSLlLgeA9kZQ9CxVyjV1tQ6x3/xgLmz3
QqjmFGumWMle6+mHAasp0bRu9nRk+JRG8BpaHqoFtSuXJDd5YMqBzHBRgQGIN75J
fx8jWUlC0IXUJj7G/O1pXKlCDC1Y4+XiqgYRKBigJNhYud/SsxjpFU7Z4NrClac0
/6I1J1XNl90WmlHmtvfxAqnTAR0/Fpk3A4E86t7j0CQD76ej8BXWxS6yOlY6QrNi
fvF6QXcRr5Ap2wfhZLtmnYOleUn3F0fyLjEImILBm5ian31ghFzirWdyJ+a0uhyy
jWqPJauz/NQqqvJiw/f+p/IpkIcO1XFXkGgMQU95mr8R6YgVuZnjOTLIHt8hSyp4
dRKkuvcOYZKuBB2HtgK5X4aTUcFxGg8MUU1/oBu7ZT+1DZBdlPrT71p0AB3Vf7rL
lrpRcPvbyqt3r7pWIPGsY37Gp596TgOMxwxHjf6Wathx2rPGnJI2KwvP7Zxq9d6J
QaIat5vB5WCW6f8dYGa1cK70dHxiuF0kV9lmkTaQ9QPwlk+ZQ2Hm7vr4DkggF7V3
DziDK5dbiifPKkwiRJ/5sCPCEIibTwveFP7WgtdXQgFEs0Tz9KSeVtKaHttgp1gw
hgaPjnHUxUCYUaRBn4bLxJtH3qYHctzEumTdYGDTP1cbJ1iEQXfXlWpltcLtG8T/
m24qalLrmOnC+w9daaonYe7Q26I25LZ4/mfyDRGfTm26mWvl7AFkWDfAZFDTvFD0
foYUlLHnbVyGRm5R4EloodkOchcbyN3u7519HrH7y80VdnuZT2/cYWF2f9Y+Y06j
vz4+V/OXQVBv7RlSff52vjth8Ok49sm4c9MP2ho0shUiQZJOBlncF+Owm4fdxa0l
pKLeoKGhyFuWwIYdWXwbrEWA1k8R3OqFw7e7UV+n5cBChRctq8GB1Kp+Vddg/GwA
FTb3a1YJx48qm4/SYZr//mhx1B9bSS8bUUfZHU5bQZdvzGanH4vyvVafooBWFP4y
IFZXb27hAjCaZAqT9AXwRq+FJYP7eTfEVgMZZFlW2KUwrj5BjwFj/jwD3FfP1L2m
lWXpd1deu87ficjYd0MFIljPc54vo3HGMaO8X+xWZb4IN3lR84xB4Dwa80fec4PB
GqAQvAr9VxxTd29EqUsvpfr94lGzut7MWCP5KvrTBbl06ZVDgIn8Ez/O4tv24G/+
0iEW3tQovPfTTeohbhquww+Lg47qCuQEH0ChOInsnK5nx8L4GuakIJpuqe3OCPa+
pFSPDoWJaobGg7bXmyOFQ2ku8daxQkYZxBVumXLCfSOGXUMQRiHHKI2FZy0HORtI
FfEuHq9XzMqRSxx3EEIl05PaQwHAncQ2Zg1MpebYiMZqy+Kh6atXcN1Th/srobJn
l64ECPiA0cBpwpbErgRQjUu0cPCv6J4kV/K652BNz3krgZoCzDrOPGaQoTjDSt+u
2KFjCsuysYP3Q+7ATqlHBf3oHQMxVhFs6Wz99pSQiTrlQdrLLFUQKNv95m/Nxu89
ga8UUXEQsT9o2ouAcKFLKVc8vv2HLWFuYKPvQY0yZvd8m3U7VfepmF/ljxtqsliL
9kzHyxq5ueCc3eK29vQjaFlzRpHG2Bm42B8JrYBrLfUoFnUBVb0IPqNE5WeCGZGJ
1JvwKZ6UOmStH6DYvh76SqJTr4BPMPspEmw/D3H7NpoXm6hjozSn/T0NtRokgJYy
6rPCWTrUEcewTjHdBR17Wk/wL4kEkjgTCjda3OPmZrya5Lx78Eroz6lavO+aQqnK
XLh5Zt1YTcPugthb0pOSld+fwIxsPffRipANkbNEKW1hLamQRS6Om/l0ZoyWPyhs
zcPPCRBGsuo88NhpFazZ8zkP/SstCNV70+Ssdu4Qz/X3o0FHNSeGNN3rdfgRGXwF
WJyeCc9zm9f2FtmHOH3hzU3Al5DIVyP6I8kqQiGjXGwyxqnO097GuoClEtww04+V
2d+cZVpyIkaKn6F2RHtSX1s9E7TG7XQsiVHR/FD2mFUppxOxCmFvM04w48fLLV6f
La3gmTVcHw9VL/V6buLENPDJSwcAGogbYbcFxH9DJHREVc6H5tPO53T0V6WlvBo5
KJa1DnnypVzRfLRx6y2jiPDUA2YD/wQru/AmzPgUw4jpCfzCMVzyG9ZOIEDX9v2Z
eEhbJjhGeX/JraOGxw+EEFchTaCTs9b4BR+fWiHdCEpHGopELbekZrsXeoOQ7ysn
CoHK0XKzsFb8k7Ov2JZPOSyVgStAfZPr51lRnDrRN+9TFj54jFQqcMG/zJU6lzlj
+wNlH3lZp7aRZptaZiJysIJjcyFrwPTx8PxKhWFbvrH8UjB5gC7GxBlWjL3oQ4aI
z897aXPJi6q8NKZyDJLYtsNe7vVwneXbZfsYnb2NUc9uvt3dab0g+UC/jcT8Qf0T
CIf7aHuE8CiFAKV9E+7EVMneQuE4RRN9e6CgPKTYsxTvasnUvvNio40w8M5+Y/Jx
2JAERdhQZI/oeJL4CkVtUstRwwAniiPZKKWs/iXrHv8h0jRB0xlGMOo88nF7QADe
S2L0WE53uqPX2Wv/wjAkmQUf0IaHF6nFG3nTRqQ2YEIn1cz1TBJfOmFrHwfa+gTI
fK/kubiWihxNtJbeo+snUDwQywdnsEwI1So2eX6vT2zrqOCMPxpfXetDugvLoExh
8Y0Mrxz+R7+/ebGihB0tq+zraeQXniTN5xhl5bEEPEjWb+CAVRVMxLfcuUYChO9o
s8MY4m1OshToLZ58lXO4xQ==
`pragma protect end_protected
