// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 03:56:35 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AM3Jd11ycw09n6cQLgLVijKgzIotz8izjavxXX/PKsSLdbnmof9QhFsGLrURcg+f
Y8wEicB/1c5MiWoQH3k4pD+KX1SYGDWflv9GWikbR8UohUN+ofDPqkWAf4oLGbt9
oe4qJlDFQavWLgqh9dMJxuhKY84hL+WCaTLJcBXu4aI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5584)
LIxiEPzqdAlJP9vW6HSgCcWsbD39IZ+wTktuYyO+ebrhEhcZUDTp86KgEQQK/wD5
vBRVwZItJaFdTtuQjO2R1ar0FZ7agtZbZeIq4WfsphRbFWJJMeNSwk3g82v9OLPK
fAQpaDCQO+9538+zlfEYS1vouTaV1br8qeqp9bkwHv4BMqg8keM5wywbEluz98XG
F1/EDM3Z8P0qslCUJjNMzzoqRrJAFg20czuD29dutYUdJsiCvuiCUNmiyPLS1Uiz
6rLaRosViB+rwlOlvmK8gza5tr35uJdmQLm62rVwa7TAKIWxdgsyc0YNCem+j9JA
qD6SDnCUg58qWTqRSACI/x5v6/nPAabNWrdBiF6CFjO0pMiSpynWjDV8a3FzGxEZ
HX7qVVyLJyXWrX7P5zlTCmITkwZm4EUDJXeU2SgIoCWf7ZJi2FqHSpilV4HjzWaq
aE5L2rSqelhdvFNzCjZ41P/LFRR3a6FaS2Y/RzqD2ZqpVIGVeYdIufpTNP4N6qj3
Kd5IH3dQsQqylpN00zImjPY8J9bOmbsLQIB3mnmNb3XiOLny9v8j6q4V1NSdCpTK
vJLYnAs650CSMRfiOCXQzu/Q3E+t1Jz7HVOCSpP+pde8X+ZdAlB6cSMvxcgZBk4N
QyLni0FfraIpSey9N4ofwhBM589cHp3JdhVhoR3DjZjtGZHzFnAw2hOHLFkOP3+D
bDBRIqcc/yCFBs8l6Lbz+0N+zzWKsnxitY5SBWvr4H/O/9Y6t5mjA7RRqaNZMfFe
fRv4+lrHX86TpPS+Ec0wul7khL3JLmleDX4A1zOl51NesaSJzhrWphiQkPVfWgW4
FUC+Wo3DhG8SeFIqpdoJSeysIiOWEh+iB7LhoNZRrIJDdqXPjAkVXKmTTUxelXx0
ir+MVi+Rm0ucOrSVjFBmbfIkVlGSL8MXaZlFojRE4elfEdtFVLhpiUQA3my3OSUd
jOFy+Z/WXVqxLs8sz32OQr1U/CTrvWw/w382hfY8zW/MoRNfGhdFJ8uSJ83cf0OP
TPbBAam/f3PVGegUgS3/a2BLdmJ6fHPIgtzi2073gi61XKwowC9VIb9LgRLp8FQr
l9Sto+2bvpavfsVJ60d99/3Eq9UESoeghfSZOAACwTPB3aOmZc5i5U1aMM99Xnj6
cyAd7QSTvHkm/kCdtdPoh797B63wNK8g57I93t9rMvFCmZXEHgBqQY4So32upd2B
5Q4+wwXcB38tkKIrXeiAzr+ACeNBBTdAm3zwx8BLYX9xyVh6pubrNZde5PCURIhh
YucrgYm2B70jFsqUFn0bpmt8MlO7QLtPJOSpbpRmpWERTPGC/oulE9oD9+fdcH9O
t8275nzHAa7PMvQi9xwMwCeMS+fR7U7lw9Xj3iIwjskVjwp4qbd8yDWii/KK4S6d
qbI+rn9gRhtBWrJ5dBOTm4A046luuP6m3HqZePx7awpWges2wKs1iptnBhIw3WUd
0gaPVChmMWofI74cmhxCGMrkvxHxJAnGuNGIMznJhsSdQQv/iCBdL4aM14VCk6KD
2T36juSs6HgGqOy61KVTkiN4omRUUpo1oGiSube1+9b0gnztYajtOkJIYfYyZwB/
Drr9TH3L5BWT3KG35wl++XEGpsdWnfH7LlN10Evq2r127e6fvXv5VRYtyRd6hLyg
4bKCbYXIlw12IDOhdh/7GhsOXkMMQ70kLhHSR3OleDrt/cQGytbtE3WvttFfqZEl
XvoYsFRScEmZDr9A302wIMuKKqgEDEO0XyeyzOhsiHYpmHTFanJlTWvJiSGhhsGh
0kfcqiDP6JLdAtTzG6wAwDbHwhgWEMNnhvjETzFwGljn2qAQ+/x3nHvBm/XJafRw
dj9CyRof56yrUJzPqNpmw50yVyYkPivyDDXVJsLntQyqYqj4fIWS6vSUj6KUonPF
VPvgV590uITQV+9SKGMDdBL6NP+TzMS6DihUllMUQ9tgQ4gimiXwVW3Wt07fyxnW
YGNQ6QOM7ywLHhqdn/wgI5evfUcophpk0oOlQSvA2fV15DGv5+3n3KJH1VIRY/ZF
EWjY9BwRF+p7QpchupJp6li8KF0h6/KjTd2jcTkPgGvjbJmqF/LZsUHjvYvP/CSH
T6hryCXXxUx+YWTIt9mLAh91DxJERdTcO+t1gBxko9n2/5hr9cHzdgbRh2IQ6L99
6nAdcv6PGlyGgDo53Trwop8PsCZJXaSyE7F2tiWxb9dAK8hTnvjinDktUxN3tri3
7djYRNu038wO/CT78EXDl7sPNWi/ar/Ij+4qMBFEcNyq4ak8tM/+V3d3RvclHY3/
ocdiyNAYnnr8Hxrnz209HteHPe7yIN0mT8UCW18JxnysO8FVOsRdD5SBRNd3LXMe
4YTQ6WdtVSIvGEY36wgw0ZjHOIEyGOJdmf1szMPcXBFzPGuzjwqnJ184l5R/7KeC
+Wbm8UdOAYYb2GEJwX5shx94uKxdg1fVbM6JxlKNArNEYzaN2cjD6U8m/8NpOvFR
I/vNK/wdyR2bwv+CpfOosL6olP9vSAVqkJDtUEn7hD7ie9g1zFO97osCcs5C8gMS
Vt1yV9OUFuptyxpxf5BhySUC6VxZlRunGvK6R/RrXwSlpngJbSVrPjfRV9r3PEXq
Xhed5e0a1fUuNvsKHg645BZa4zQNuPh/XfSM0AkRSEC47jngjZWuc3tEms2sxHDm
i24g4dFqdksojjb/I3sV7F4iAqMIrG5tdT8I/YBL/INBePmhoQD99gxBGLy7oRLG
OqwWu8JgEUCSYOUqJMHj22flhE6FL6t9r4irPiaDYXqRQmhhHlUAOtjonPq5C9M9
5hUYep1UkbnfeMCz2JtcR3Nn8sdnPE4N0RmXWMOGDEdEhWrAVvnWvfuh2tyQ74Rz
7teOAkO9n7gDEDYR0+/rqRToQ4G8xJn4c7sbxy9XJX3tKIkidJURITybFWZ8I3+3
S8GvRFwXOa20pd1VZ4aNla64zeG7h2dLtlxdF5xA1Xz+pXBmjLm+NIO28B8JEgnF
O4FC83lr2yupbA/AIHvEN76gugTgUxp02h0m6anzqOzmWj5Pdgp+Hhq9P/zuG2PI
SfNDirwidv8LY7q+rb03Ik9w/EvAytD5MqRUikGbNN+ewmg9pYxqpvIpfm908KJH
TLn2h3UqCGQ55c9ipy2rnhPYk2Elp4BOLJMMogHnNlMyBKwh1iy6aMMMhZXs0hqd
1d0fIoM5AfZWpls3MUy0adu3ZvP7ZMsRXIf2SZ7baibiWU1Fj5XbqLMkvztmYUso
DuBWOQ0ykDV+dRx4yDRv5ajlH2IArI+2drmFNpILMnnugkH0RwQFCVdX5GDBsRAI
GTpDk8sftVES5rKzjTzFlo1nkAaWMk69z+j3XPUqjMw96MENuqQ4nAtAOuKiLaQc
ElUlwetWd7A8A2R9b88AET6R+fnKPR0DEN8KeLLZ7Bd1oQxvNMXove5TEUmAfExh
o/gm+ltJlwcKSBsbPFOTduVWhD2hWC6OJVMHXXIr6BwmuRLXW2MxbejYjHU23dOF
N8C+hy5L+XNAeD/CuYIQXKs7Yb+437pvYs+DYaFpV9BDfqPFVjI2PStl2Yxx2L+1
bWY8/l7V33Aor9gQ1pFijEXTlRxmfOhrykwCITW1pduMVNdyannHJ+Ngw7pLZsCi
k88F+N/CVwci3OSmrPuWqT0Qz4q7nmVDJkS7q7DJntBAHL7xdBE3s4QnbRnQA5f1
DGPluvywzxxWdgEC0UnUW7c04eGWAAtxAXWH9IWZ+YtD7ntl4W7FSdUUD7fAVGDb
WSFbSkuUj8DZ/df1LzWrwYbXLGPSsbh44rUAizGh9vq/qCWZZpHZLta6UMp/lNlQ
YkW920LTTCfkYzxrBEn2bVJstyFS12QM4OVoRQEidm5CAJgcOEq0yObTaJusE2vj
HrkhRwWC1Bp8J9SdAEv5GgbyO2UG3qNXfEoimUudDhISyI2qCoF5gtwiOIk7pNxa
9bzZy8Uo/aV1d3MzB67x452oo6CS3gCAoPiOfKrjFKoHG5NdA0oMcNCqw8yOfaMB
DU9wn52uTz8PvpACGkyljFhI5E/PxKCLRKqvG4DjDCiIE2jeNVIrKPPrxcpVTbI4
IOLTp1H1wrjf9AjlePZpuUAJhzM5tIY3RmijlkuRSIDo+cUTrHYa0EcvkzHJsbwj
LCjtqxfNfeVREUij0OWOAuwAk4nV/lX+t+8X4bxPEvBg0mxEfn4bWjR4/AH3ZFeB
UgXgpxj9pm1n5WVDUVM+HVKCJ2LLgwFMzOPctQ8bnMswqFxCK1SHM6dXoikQgGHG
jJrYl6m+xDjbV9BIB4spG4Xp2i6OV8+9OkLz6TYS0qSpFE/LXYllKlrVbg1sXaV1
V307w67gzMQl2YCSmjNf+GD72rtF2bgZzvlNVs/o03Jo4f8z6/Lak+F+xZZfFtHj
OOtddMSSmngZ+SaB1zS6WnyYciTFDO981wP3rVUkUhK9O3qyGNNJG7XbWf4G+Uup
yhPkwJKK75zxfWJ0B0sXVUbWD9Z8PhfJoZ8Qx3inRAtRqx8eRx3rSOjcu7K3hGQC
TeQUFInSjKdkbwtLuxVRVECOpDWecDzC7UDnmrgtGu0j1WR/Sq7/HyMVlyX/HpzT
Y5HOotmS4SIni38qffOr6UFQIMDfQyUcAvMXBlB5rANuUI7BSQqj1PSPvepux8q2
m6remgzstOoo4h4yBl8FToXbBxLZMHHHayG7DDZ2agFJwlURW6u5YX/kYkgw3IvA
3kBnJqRRgLXj+6Fm27AoCk2DLzxYSlBR13c6DAGa4Bu6kqjLjtG8xiVEIFR0Z2oE
coKiYZ3ECmDa8+jzYC+Emepe44LzLfltVb6M75p/EpXpfoCmxB2kXXupJjh/7Osf
z9WjpmPKt2aVVVgXC7p7fMb6TUnJxp9kxqP1Hr1Ww3dPSJyU9FzXrL5eAOniJTCn
1OA/VlptvKXutnnvMsy3fw4DvRwT/Gmo0X8k+54UfYXK0emIEu7HmXN9jvkGz/4g
rzIVM6BCNGCphsfcNj1j8J8wXG+ifzoJB7yIxP0wvWQTuk7E+7T1SFkBXBb/mQBA
i4bz8RtV10lZuT/Sl/3PsqJg4gDaEixKPkJ7hSQ7YMZD9XCni0ndaly6UXyrRQdK
kNlP1om1zOiq4sw0/ptBndipCiDtOdRoFxV16KvnkSdCOtawKiJGEop+DF5q5RRM
95zDsoHz98ztVlDxEhvZMNksBH2uTnG6DMxCkeEkLudOJwznCQ96707A6DKnr0f6
GYkxtAzL2qW2gW5ZkZKq6mpoMYMpLmMGWeKcxocwUVgJfuqNmTUS/EzbeVLkoH1q
Xez5U35DT7VdGKpyDkjXpCN9JII2f0OQlQLhBuud3P3G4ng0YEfwveIkZRJ6eMLl
NmR7S0z5MW0UrXanTpPMU2j1Kq2vOY/L9mGDcs9VkPPXfTuXvboog0PocanWBehO
dub7d9aBoJkKQ4tETAqbDqvUePQAjQe5qvUL8tCA2Gj/uSUP0yzE0hJfWUfWMhEB
6oifRMXm06aH3otKg4Wv2O/HV6eJviUdd8QJpE3GS2QPfXVvaLUUOLcB3f5ZyC/P
9i2IoqmhTWB+N8SFO4bprepggHZMfomqkinkbbkN8BARnLZ7KHYrCx3gP4kH9vIz
bteB1DO/mXGmFwdIeq15aQQmFYsr0PAwyp9+yNRvtcrhpTSG/badYKWMUzrx0Ldl
fuXrYLBk9Ah7+fqaWSlG77EZ9zyBzeQ6alQXVogqqxUK/4dU8KcXyTs0K13vxa1P
252YpKjDCxtzZwrTrNisIKKtn8f45x0x+geQHwEaPRCW5gB6JWKmjCEs/P4pu/4q
dYX7Uy6Fx/OI5+TeEqTLvZtgqDCFPJ9JHN2nOj0l48ocjW/tVhecasv4jQf0FWIH
y4bCEN6jAeu0gm5frpkvZEfgRiE8GtOLCJ8JGddNcTXPRs9d/H1pATOVoepJWy65
XyMmAjR/uerqZBbjm1R1PTVByDpmR8bEJ3dU/r4enGkTt/7e7Cd0ChIgj+JIkOy7
WgaxXmj4rNA/9BWVt5A+T5Pn2ZZKood5vlq2Dh/0LuhB0VOq3CkQ223UpeA7g3Zx
mdEIsiAEb024SXnMfJFJ4rU+1SUbWFoFnYrNnQcsQW3dw9wheSgjcfIYZw1buchX
rIt/bBefgLDiTmEtLXRe4wozVUM9bkyUDtDPsYgdrewvAs0CkX0qJpXskSf0E8pB
QthUgCL3W2kCZHLBsVjRbbGG+I+KGwaVMwTI2dhJ8m7N+bLFgGX5TDrFsRVa/ool
5GLon/naj2Tb+7QkSHRTj8MBOZPin4KvjUmyw2uITqtflU+qpYIkrRPFegmkjW9s
h0Nqk8mqfKz83OXEIZqE96ZxuJFBi0g/0z1VgPO0rRcPkFFFR720VdVXuut7xAQG
acSdrffeqq8eQa14R4w1S0nF0IgWcJnH8NfGrcv31YUvdVU/8nWPHo/F+j0I/ETg
+BSVOpysPxqt0Afa5QOdkPe4T04XBFzPU3NUra3Oc8svBUcO6AcwQiOTl5lHDlxY
TRZJnigLTGdT0J9WztCYDBjg1eLARvi95LP3dSSu6DeZ4iLEU3Gf00udbCDahKN2
OLBsMRqotSsboT4dJDPxr5PWJHScTX+nEWDC/dbJHam9kf2YyyPRm+fm1yFn3yS5
rL56dYogFmH/tSl2SvmWMWRbjg/HQOaLhtW51muZHkh15kdMgqvRZ8wp1ytc8NHJ
n9Pd7uEFY0ltuqd6akFPbPHsw1X/XSfJU4oDJ44gXb2TwsnUaegnIa/jte4QdwpZ
AlIb3yMGZGbR/PdveSo1rMuCQHT699aw/hYcFs1JQgVxX0NDDDiUIECngPS9gtl9
U3hkB84qVcCTJ+98fUZRDBFEgrGt1dY54HeplQpmnb7w1C7/OajXD0DZqIRF0exJ
goK3Wq4Sgz1ZHUsVWrP0gXKQC7ksRBLU9NxRTryVm0hCw9ITIxb7wzM3jFsTqVaT
zXynoZtnCb89JVtcHllv13jDBwGvgMExaSjOGD7vGojlSUNxoIgFiGK0+yIwU+bW
BlqhdXzgmjo/MYb5fjiX7hkUmCr51wgH078eHjDtSs95V6hxGEYuxu9922iJxrDt
ovF06XvdtdI9r0LV/DA3WtO42P8Eiangr0XzTnqVr71nDijmctGfyCv5d+b+pTSf
YBjF4WD5/9obFdBN1smYc+w9fottN9qKjDQKC4z6oauOYEEiXkpBrd3MQvZHBljr
nas3F9X/ZYYf5ahjmHrdw6sjY8foLyqAUFtp4yLuC5htWt4KXO0Oy+xO/Po8bTGg
iL3K7v89gXCOdViMOgLdyOvDmRBJ/YFHEtSTS26TEg0PTfGNT3JSdE57zaebU5/+
lVeXwA0b/GbtL9o4hgq9QHFgOMHNwJJaQDt7aty9WsCvJQu5bcTgOTsKhqvEubKp
LZH31gNmeZRn5M2nHJSNqw==
`pragma protect end_protected
