// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 03:56:55 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
X0bhRQ4sVW6WDf46Cl2MxYKQgCRpmk7lPWTzK+6IkqgJfgysL6UIpKhoaev8WU+v
7NxvdcgJsZBKaBAaDT/ZZqW9+UrO7wasDauXURLK83mwEkhPB+Bx4TjUDD59TEEM
2aRnUIqBCsLFpNpLxLLdPLMk3jKHdsfx1wfmNiAYp9w=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5408)
Gj9v1WPczs0Bh/eUbfMKuCaMNAHYGU/7pvt1lMtT8uWkfcVnsfvdjr5HJiP5brzZ
tZnEsZj5h3ZL9P6Fktie5TacCeiH6GN/109wz3ZGcQe/OHxozoW/l7r4Al4kXY5k
VLurWJpQXaVZn4bWlHssfUlvskBb7J71ky7HACTQyysFbWh8w5m4ByZt3R3Jqsah
Y4hMOUBUKgW2mmX8zYp7P9lGmcGfHh8oR7kro7JQmchiY9GtIfdRV8x6MsBbGL51
JmdBhNM9lTjJLLgLlK/Bb9eQgoz24mZ5jUZFo2QqsNhyrYviXh3Ln3mBF2hJZD6M
kme4AsYwamtUnCRLDIqviifWPEcALMZ9Ez5/bCTgO4RPnzQvrkGSVNoiqGsm2mr0
MoKOArYITdq8eC+mculljysbu2wZGCjmU60TMwu9d99PATxc4SSRBKsvMZ7HMMM7
2O90b6D7wgsmv+3EkbMDSvHvaOfGstnW/8mF1NCPo/sQ9CP6GG4NMqNJqDoyv7qm
KMnx4TWuoeI2JNTWAyCCf1zntrLBtUXT8fWHbbU+LmVgY5oOwfafPHU1YcQzUxUv
62innfMveFnxf3ke7DvwT+Xz272aO9N/I/urLf+DQolkrl6fiCt+QJBAnjF7CeSg
ngXeFVjPtB5yh9iXwSpNqw/slozpZpPJ5S7z/60CTq57T9gEn7OYYscKLmBBddHS
P7mHXoD8GzUPp1LxLtLnIF0I8c+bBkfMxa7zMI+0oSLlO5SYpvTjUi9wtIJhXWFx
4lnrn7wowzWO42VgeTha9Oz4huI9dy5xeU+fDlIv03xze4KMPjuFw2cOuxi6zFPg
gLlTDDWrtyG7tNJchu0c+QyMhsIUNkG6oghU2djntac9JOJeZrA7kBpE/zeTWRhO
Gte4vpLb5GOC0BPTBQG2GY2NONcm2u3k2euTF1u5VONCyAfhRZrKdzCQiXnubvRh
T+d2gWc1gs049twoOat1ScuveiOPWnhaFu9MCP567qN5er4oeQtQbZSTEc/llg6D
rTVZAe/Pfl4B5HQLRuOgmBiwVmSZ2+rskhcw6GVqLPB5GcX+WL/Ebry9r2EI63LK
36fKE1xrUhiGdKJbKaWdex4JBgocigQlRPzRf06Vs/oWyAyrAaMUNqJjF5/0vPmZ
fnm+yl95/plc55tex4J5ufVbT0Z/ys+zL1oQUJjAuT3K0uZ2gIP1AXLgokKDcgm7
s59hgmXYle3n/sHG7Py5UijTiiysCAsXwyETy2AOmCEV9Wv2HIR8tEEcPw1mlVhV
N657gSaXa0rZ9Kqaj/Ch5IKeJ2LjBCQ8tjRJXJ95HC43lRYYv8oiLK3Qq0hyco/g
KK8fBobixfvsmBdS22OolbzNdmmxk2hgx9Spd9WDFxmwxw46I1YzYJ35Z3YgjWtZ
xVfUrmdnbCmSXjYi9NeA3kGL+adMXcLPxvjDWBqzUnxvXnxtmiJWXSuW1HafKRhr
kuJ5qkbngfyYgTK9wPJUsttssBK2bwdVrZGpbLfM8fGf6rDwOFz5kfAmwS013HRP
GIRkGB+tNUZSihBUcuw6ceJ401vD+0c+/OqN5t+op5O2/DwQmHAG+prtZiIuF7UO
yGMTgOE9SKRzSklB8jUd1smXjyc6ZCusb6s1QP8sMj9AmYPafWlG5qeX38RIG0QQ
juDW5uNuByKaOeLfWlhVXUjUIwq5MsmqkEhBmlTU1fStfPKII8c4RvGMLpO6ok3L
g/Dmc1jAabiOol8taBr2Y9OIrV6Mq7u3hG1J78gwXMFSYSykanMODyXao+1RPQXF
RznCZoeZuXXjXvnCSWDBO8FMGxRxzvSAkLK5haRmFLj8Tpjz97Zl2o6gsCOOaj9b
GaKG5xENkqy4SBfTVHmJjklQa7kOkQWPM+T9P9qNXPLe2uyTsLn7WtJXygc8CYEk
ULY76nGlM4m7Lsse9EwyY9P3x3H6Fa7xA/ojBvUaiu3xMtoSWdZCvbBc/7am1t1A
hZM8mGSvCj0DRqGJV+5ay/7SbVr41ftHdYVXBYGDEUFwgyhKhyQgBn5LFTWKSRVI
hxqTcyCl5RWDaFR2bnL/CwLklcRWkow7LPJOP1kNrHWewDz62hkeXDjt1ow5xkKz
PLQc6MEz8qW65oGwCkbvcWa3o8Opvdx4p1uICQxkwaOyJEhAXEDwBPNi3VJjtiZj
mz8DSWkgF+1+uHm2k3UojHxU7K8m5T2AHz3nUvCfnW6e/zYgDp41Gyj7xXw0Ei8o
wE6MCwGMZj6bauP9VWl1ovVrXSHR0xFrZavN0ktfMLLehnvmOltMf1XOwmPPiL4c
0aZvXd8C9w4m3J+3BFx21SxZ69KEaFU6TbnLh08ez91YP8tQvjwHEc9ZHMh7T8mc
JzYCd+5E+B3WK9sQtT4PrsKvwypPvVYxLN1gUUOJCpr6cDE3f4Qu6Wcn6PGXPdA3
SuoDfIhdY27g9EpiSLN+ZolRXo8WYGNt84gWtHc6ZoO9jVc1IHc89BNRk0Qvx1Gv
j/kmyCwlUzUpCHhkX+jISPCquMPrR/CAsDCE057mraSxo8AiYIa9AL3kMkW9WWav
OCBpzwMZwqayhpy71A87l0+qgBjXKt032gJj28OGMaWle6hUIk7snhzM5WaN9IZD
tnukF0YMTmVrpI/pOC4vJlFH3rdWzol+gP16BIvzXi6pOHd92O8ggoEcCIcvwDIR
QMAv4otfe2336TTr1+4xYuRhQnow6aOHYXwO8YeACVeDe+5WF90fL4nlYt8lK+eN
grOMJAWQ56/ogoaT6stv83e0rG2MygEuPS08H+Lgs6+ByZ0JwzWXjQnxjhiFo3lU
ZitKWLd8UfXlGVuWSUrCu54REfZiKDnYpP1S6+ov5H2uNwtAn51clc1pW3SeFQip
h0WJVHr+j4Vq/l+fC1T+HBHE8kLDFG4tyzRuIDIjqpn2CyjzdD/tu9XUr8w65L4h
9BjFlr5mz9q8s8DI1IPPW1PrVg1ZJ5WXwSuXXZFXINQScZH7wHXaoLIDbh4oeMCy
LAli1KT0Vlo2UtnuyQMx6WTWiWsaa2ZRVJ7lXdA1r9ecddtDI2ysaDVNAO0n8sXM
rUzxdugY/s2gZjgUuczkVODHjAHS138uRD53Til/rW0BA++yeZ8uIl1I8dWaHWt6
iLYXYeGzl2H3h6NVLeh3rxUP2LoXBwTaOcqkg7+rT3rKuj9XMUp41JeGijuE1B/E
0lrs4DI3E9d9yDM0GMVzh2A8E5nkTNhTYhn7IXIaV8FpQJq2SC/rpD+gVo81xAm7
SjzbZ2a4jWkt/dicj5Ycs6qQDkBg0Yggq/khJ02DC4lyMDzMVguQSuNQwbArusRv
le2DWBzKbB7EFTvAuv2kVMXbLQGqcNKvOZQ2bZQ9K3Qu5w+3i6aKC0ezBACYFcCk
EjiURnszZ4WXK4k/aHa+rYUfbkwG1xJM/CXzTffP0MhlsANv8q07xamlsduxFPEm
KbNWCdTkSkpQaVRutoXghJ43BBtRVqPK9rlSFkK9MQAC7qF2q2BkQbSxwoPwpyUD
33Zy62a+3471zrVl4kN/Te+hBKzbMn/T6k7/KdcXhu/OC/T+2YOFTFQUm2VoSeI2
tMDV5s5Lli3ysxrHjbb+SuSL3tf5V3CXNTKlQpqPjq+WudUhP+YPHIyRkhjcD2Wr
IpOHSs60woM4n3I2Zgf5G2gxMJLVa35NeSTOiUnQxSGugXYmQLtBaNTXeF+CaCQL
8mQGKesYgpAAR3PlulvK81I91rS/3o4P0xHCjC4CDQCVDfLLAXgTUPHhpxTwCQMz
HLFH5LXH7/g/GYxCEImQfvlMYeNKT6O/E2q2mj7sK68Q4fJLbmMbQdgS7/gK4fj1
Z8MET2IPt9KCi4rHAJqTkDcfmoy173wnGVz4HbrxgM3KYGl79UjPzvF+OvTJV642
YH6xYOtRXUDE4frVlUDFLjAKkr9W/wJyPn13H6cGkzCcVEZoTsw9oiIj87pEACQd
mu82tbFNOU+ZdIPt4xIF+R3pIIxIacKcVTxvTFiFf9vqCs940WOddfcuM77HXvOF
oRqej4PtiQob+6LCkpEC8HPMQZo2a/8f8G2hgvo3LTiMUqVwqvzVO/eRPfTOoPsL
wDds/wJpneY0K5znaGYMbLcRKdgoFCicHkLzeUNX7LqojgOT5v2UKZBw27e09pcA
xhu4oGWxJ73ErCBbKhnCCoa8VIJ+FVWx/i2mjRut3vu4KhRFiTBeg0ukW1TBQYXO
gDVCgaYDeiqg61CyIj5b6kbgYkzHky4xRLBQXV5g7D5YzdMllH3ooFfhRViyTHQ+
7GtXZMMvUWu0wy73pXzNwzQvlQerwQp8sKdxtE6raWi1S+Q/C8/K9aHassDWPkUJ
9wplS1mIdob3frlqzA1TGrKK0N/alaFGeT4Bio/vqMC8P/q0E9bBhJrrdcpPeNqf
ejJHjgSNOmZLaxc+uStC2/8qU5wtrZeq+gbp2oo0l/EovK2eI7C8vSoUnZrK1fwy
RcLzIu9CCRaQeh+aq8GHYSa3YUq3HxYT+4SowjpPiqEgIFbcxlX4IFj2MiweYmZC
SSruIz7r69EAMdo1xZmK510WPlOWUJPx/Mef4kEw9qYsK+YhPCjJ4+PXG5Cj19e9
theSf4NpL6d70fLDUe6PyiwRw8NlbA2G1mIJF95g20mG+TjLeLghDNl6D5d6S5VM
cs3o6ExQSjMYJnbYzdztGcTH6gZDuJIR9oqHWiHAqK8K1vNhLi40XORdWK6ucHBd
73ny3tUm5knLf2bToeZlCaLSGsvkvJXs/WI2y7eZ0ZWdqjfKQnavCE7+Rzi1PH8y
oGkQmoR0uRvmTaG7O9uWcBPqY+MqTpqfsSsvs2q8x+1MsDj2CI206o9P5wvc7q9t
8A+BpGGNGPruU32B90p7c0GiwY1GLIzQ81smpF5bkiDjhLC45tliZsOBPp8yfAPV
tYKqnCRO0i5FVRQnv5hQYkiGR3uErqn33rCC6rlNwNAlMFPvUWWh6Wev/v98G6G9
8nS9AvAf9niKbFOPwWgkZ8Xmo1G54zlDEg4H+F/nJjh1SP3RvdhHL/+RfzFf/yaO
igtW34XsOQAPYUtdCCo4DwvuNAsGsnfCWZ7CIZP4hadSIk+oscgjOOpg7PA77Q30
yE6B0jzIYtyGHSJCRO8DOX5bqPxBe+muCBsN0sEXdOI8h75AVF2jz8ancE4nLmwp
O4ibOpqqGPMYWNJSDkWt1/nReO3oNDhr2R64t/nG97WgTRgGWYMu8NzvinGYgWdZ
7fb6unJTGZTu6O2yQE8O8XvLd7MbW4GG90YLbVhWvwy70NboYoeYNvR3Hi7H3TmR
af6D4GhT8aQqsSdKVMXjsRHXG1PeHsFqAInkv8DyA3/KIpImbmKJPJLxKTus9KeV
VCtHwkkDu3xlLkBGdvpzbiVpICT9jp/D58PgkV4vG0dEmEhmFSXY4ubc44LOVDS2
VcY9GOeyt3bSZe9qYczJCLGgqK6rWrHilA0nH1skuHKylAPtUfm78L8LAnRB1ZIB
EQ2XKrZjng1Yj+K27II39PBrrbZsK7vGoITDHdTeCV/AXY52LVqBrjCAy84/V3h1
Cq/LXNbdZMaNDDFuu6BtbE3oIpOVraXBO9PO/f4/xhUSnV+/wGs0fEumb9Tf3vKD
oqsFEzKGtPUP8TDN+SFM+NqN04QInMEIDn7WT+gaEa6tCjAFLfJ8uu8RWP0EpIHA
YrWBjsy0nN8KVYty/eznnolWqORGcFDAPSZtAVCG7PZd7h34R8eCNFyU2XHrE9Af
MBP/50llIw86flUuVo/gOhsp4dHY7tofVaVbUtqr79YkYweD+emAvicwVphTfLWO
u95EeTPLZ3aZByNfl5rfS2pPI0vrvfuTSkv58+E8panus7rkpaOVp769AHzj79gk
vCU/I5h+wv4Raq7pWcKqY4lgGv4fiyySkaEYn2OgK5scmP41cIgdS8CTDgKJ/3aU
KbQukD+5eB2yRWgItx1Fkp7aO79RExjVKdY0p0cpF8M5BMRdy4TprMp17iKSePEn
86K76VI+7LZtXbcikTyGWkXJxuezs7FB2EaqZh0bbF80zEx6ddyAy4lUMzYJhjIq
Pk1nmYZxkN6GEFZGbjddgKiZ2+mRs7fLVN2h/JQ92iLORVb26El7FezxCcmhmwaj
fPhANHMaMzorOBADHuhezwRPNwNi0zBY9M0lO2+hJryKbEOnRFlFlYd3hpy19Vxn
ZTVocK59fOF8Ple0rbOuKp4Fu2xrfPBECy/yKXrKp9woRmUYwnfjpksgGo9y1s7/
/M89WwRUDKmIUoESH+oZU7+ITJYhhPoaFuAqSOh0NVtUh3LBR/rTcBzWoFy+0Hiw
nrH3psb30Wz2TQrwvUKSL5l4VT/q2H2ckeZsE1c8dwUJJ41gjI+5lY/uNQ4puMCK
RPTdIEvm7rchfvH3GQSi8urBBiRSjUOfnvrvKD9bXa8OSK/NQqsP6mVtGpiT6XSU
rJ46CN3kXBK3itmMzO1HTETGsamhElRDeA2TUtiXNWTC5erHsU8V5WsqruRE9bEF
GKRjpVe3NrOfC1aeKI4dheodGwGRBoag8oAs+2jqpdAipsYTAzEGjlUBv5r3XAFx
FaiXQ+pj9TQ/SMAvd0JXWd/iy8/0snAoh843yh39MHZfBeOL7sS8D+YWzwq571Co
wfgrHYqLMfF+gKNvKWhRaGbTsZ7bpj19n0roBkuVjnHlCHbffX3mw4MDtEuOFzaC
wIyaioM/6e1fm0TC8syzA9xlucscatemsF533NMHXjgSRaJkQTMOkmaAQmoMeh3O
Hj/HT9qH+hN/L9e53kIph0yu5sGhc7cBlsdinRfxfexrVVha0sna3Ni4lFr3kmu6
WE6kR2iO4X8uR0ZFJxc6ojxH95aSDq5z2LCWD0im/s2xb+aj1i8ZcfOxf+H2kLwX
vV3xGzktFUNjl0cSt4zIWBxm32dNKpRZejGSzOxROo8hKsE6LQF++phICWCpNiUX
tpqzwiXfACBz7R7fWt3fqeSxt7H38FxXzhr6NlAzaYPymfQv+No5XuReuXg/JvKj
YxOPY2n+z+vWkiTR4rep7ihYiOKLoFH3qUEuWn/acGKOchavcaUnmWZid+AMcgJj
tAYQtQ/Mu+yIYITWS82v7YirUe1F+dUPq1aOQudu2i+J2LV7e2/E6+dWgugkMbmw
BcWaBBt6sgW+77lXcrQC/BPA5NKRGyPnrk/1Jy1ycRQ=
`pragma protect end_protected
