// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 03:56:37 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kDePI5pwa0a2uTqijdh1gcGvPtXG/AjnC+CL7Hxj/wk4NSov5mAiZvMxhPh0jPgm
L+aNugWKurG24szxV2PSe9RY0rM5xPLFyThCC/kjbYaTD+viRInZ7Kph/D0AmaoU
JWmVAWgawf7rMgShuLub1vWKdaxptht/h8s4m815iJM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8400)
oAh2tR16uBIjCrceUdXj8vPYh16jcAkrideMRQY9TDYRH8A8cKvDQdPhwcISrYLP
pihYQ6LPov3QsWXrL0MNNjamlL1XA+zhgdM505IB561a6tQFzuqF+4NfST6lJ9r1
qbM1YOMspmVSouFcOT44msZKE5mYToOZ6IEmpqA+0rR1G/esMI/sC4wBGCefk8eU
pZaYcEUESyUGbTj8KRQUla7HLjTYqTia49XluZUwN2v7jQbCtb5mk6w/fA3NsbdE
aGf7x73bn8qD9HK0ra49XhC69rmXseiUtX0eSnY/dk0sWfFO0ywj7EO3WBMO91SM
AVhoFoKpHDVtsiJfIyhe/4tQ9u7an20bqKDXMG9Yo4Pe71lB5Pn6ZG8Hmrlqv9dA
z+eEewYB+A6TrZBgnE7LcsMT9yvBMGLHRq05uEUkayhXtEheRfHLkDgYQHZq+sF/
wQLZHU/wvz41bfVLcbDzBBSFPNTqasDpadzPm06IzTsqofzIMXXbLJ5lfICRMbFp
UGzrQBo9hGqK9en2ZmqCtUY4y8WL+PXQJRp764t3fHTog0dmWtjIBJ2GZ0tkdBMm
rK3zCyZJouqCRKekVkFZ2DqUEDK3G+WdbQ7mZWMEcORqGD91Lje3knnECPVJKpFS
5TTqk510gyPreUQ/utDdUrAwoKZk2rmXM3XY0jY2yIaaGwKUa+eN5jzuuZf9gg0X
SMwz9GISSjdaOuv5w4Tps+ABiNj94n3msRcW2MG/6mkBmPKg39oOUQngIQceDKqj
uJbrFO8qhmpIi/vdA5oqEkl8/9bxUim+/sSTNP/a+HmWZ+ZVpHE38QFh8VWAORqd
zc7I15di+zzKmP5mZFTwlRoIJ8aYEYe3K5RDTLZjAakiA6Fh3QtQzXJqNsg6N7Gl
noVwiRHDJkFEHwltg+2j1CbZbmTg+dFkkzC5pMzJYnx0e02AWNNQ883GxV5PVSkC
UcflIG92qZPDaBG0OFFca9U7WEm6WR+/6ayZgnO2y05sKvuQMn/T4zFFIwuc7Q9f
S8HWhv0qwj9qY8NZ6xDYrnuxyE6KRynaWonCD1dPRTxJKw/MiosnUEO3QsHBajFD
6W1Zm+8SWOWAdkX86Sjp9cQ6PAYeWRtQwAyYOnMLv6Hrp+JeFw/85VH2vmETwIfC
VaYVrkTMmqRL7UjCAAwVR7dkhaEI0BFoVo5alAENBYKljLdZpN2oKtfotLb3WHlv
2E8B4c79IeRSBhY6fbsfS6MK+ApJSSRYn8S3/r8DorKdAWnyXAG8aznyhVSaZq80
exUs+LyiabXBfN9U5Jo1ZzoeZriNI53aZmGGeUaI7gQd6pwy+1E15HsZlE8t7o94
0xlgKnWng/jOI7HX/XsXN4cViHoPFBugjXEMhGpvWrRiOpCGz29hgfVUfwo4VUIp
A3aPyLCUDJBkpF+ZjWZkpe5DXdb/FQMbv6W5eSjpZCmsENcdAagaXlJlo3RzdVEG
4n3qmJhQxo16+ZB7grILwaw7VRwcbBMuoBzEM3xtYrA9uB4CydV7tk/iPRD22VJG
d/ietZDCXD6RtK4g+vC9hDWhAziSAZqk12xov+6vQlVnC3WQxADoVjYE6ZSQtdxu
YJf4/vl155NnG7oGOG03iPCzcsRzyyP06QuDFZOuOK93yce1cFAwpd4abPGOhHy5
kQO4djeGbcsYVnNDY3ne2rSDmLwPAbDIOCbOtUxDtad3WfMfRKfQW/CYIn4MO6BW
bWKbtnP9LopyBoBG1wLYhCbpSGJmWAKQ+u6IOpzDO57GAR1Lrfiz+/OyQt8RMPP0
NXvrQ+LlnnO51RtEViVOrs8aUytnpFvtvQknAuH+YRUJVT00DD4EuVXWtQ4pf5Ba
pjv80jr2sw1/5W2NgmA0b2XEE9zQGP2FouIUY+L0+fqqYbq0+bgGyNCtoPufzzTp
J1f/fsAb7Qeis0mKrYsShAwzi90IxZrHokjuVrM0hEYfAj0JW+xQd1JkdrMFtsy3
Nycf7qewTjKzXEe39dFxhVkJ+X6PYtjmOTfFpK0EG2UgAaCGNBlHeF8rxRpoEfuI
O1e8UAXYc1Kk/tdIUkXKDUq2DoMsvUUZJK1JgCsSzAoluOUfrw0hVlNdve6h4z/x
ui15LvUTm0f/YSmZ1Q/iEzSPKqoYd1a9ctZ0EkHA3hAhSLAqPkUyhqbiCJhlLXJy
Vg+lcDIauM+FkJ0A9vTbzbvuDG0AZXmr5YESs3D3ivVOZlk94CTxLPr5JI2UWEqp
P5JiE2rxl0/7vMkoYd/ZujH6D783C13Gx9/RcBri4icwI9bHgWZlkh/cwW/3DDXQ
pQKYoHmjqMKOBE6OAi8Tu/eTSbVnUzUyRomLL0DeaysKBWLBWvEBIMmuBQGEYw5Q
Xdr+q7zn0iAHhLCXeI89fmHJb+WbXbGvf69+58wihsNsPlWyGGkcTyuMy4AS4+CM
WUb8wgTDwY4/vTvcXaAGxMvYn5Uly1SLTLfYjkJFEg7W6AAfMo2qEY+AfoJxFzSy
DdFkkSU6q5plhO6jEa5jrlUWs79MmvE6QvVQvwBswQCfp6U30zScufZZEu49wjh0
VIdcxpDAD6qYYI6Qe8zYKjmet3U1FQZI2zi89SbfbhQbJwNoHMToAWA3SX1FaDiP
1qKCHfHp3H31zF5lWXyQia5G6M24qy5LEEPlHk3ipdLK+rnR2mhIC/9tCM6Pr85r
71kv7AJRieHi/qWdDxhAP5ucZ/HvC9/ZPtfTW/zscdPY/Bu/Sej/lbls0yB/18yq
/CBI9asKlTU78WCJFzCQ//wzWJEYbVepAMgP8Utm/3Wc61D75hAbbNp925KbdVYr
7p+oRqX1dLLzzs7wgKHRKllbw73VDOmOb1MbJgxBp4iG7xV14yqEQY36Gg0eNSd4
/z1LJZEnWNfMyDbW9zXA7MRm5Oa9FwkUKQ0FjtpjKGQ76T3vY2ks3MSowTKafXN0
zAXosVIKqJYvKe6IbJsw1VTjwk04syDeabFkH84FoM8+GEGaQFsux5e+ca4l8DGF
CVICRWroR8z0NeV3GKEoVwju5yCUO5vVuwD8kS5tX4hbdvL+XzbKI+W1RsAkSrSe
nBMa8L/XEmPnhxakOauvWshVNPQOc3gWiqF2u5nIBHGWfEDh4FVW51HFjHDFJiDB
ryHezJhc2GuIrANwvf+McaQJktJBE4YTx39cT2UIH5jTIXa/B5DJZBq9ezO9867t
DZlfZa52Hy+pk5MfwhjARAmZbAgznORtfDn8F2VmWe2Looe2K6HrJLNfWlC9ZbCB
ttZci9zoAZsMn9lrwKt+ADIcgE/nF6inKqKCr+92Q8jtkIYogd73o63yS579hEKi
wXFlUJOIOJcX9X04oylwDY8Mjzr4LwgM2ZRPYCHblwC7qMOjiYgwTpIEG5t5eZQg
cFfczszueo4nXEn7AUWAFDvbePQID4IdYqJOc/0O7IDORKS47LRlwT306lHoZumq
vZkLSCy3vNPdjZvM27QXxBiy0MuzoZ3tpS2644M+MXJjWjiKyHEP3x4fOEGOtwKg
tSbUrzW+D23SkrqZP4wycbMzQ7Ypy18I9j/LITa3l5+qEHjejLOZfKvKRjdYBm5H
nH5GmiJlVInerv03Xb9LSErpaHY6PC0lmrXh3vcEB8/aYlHG0KhXCB4lj2nvi5Xj
swS8O/M2Yf/OKqXoVOtldgyFXF2kptIDIk83KdVZtrGodYjVo/U0etS6IsuPqe4A
W4ovmoklCBBf2aYQyjXaivg5oBtRjAkYKs2lbUd+rJe4mbazoSM+Fy8LklWq7N5Y
Nh1Q4R0btX3cusHA7h6cVnBJwt5af1+sgUIw5FXYEXUmlAvzg1XNdgiHTFC/5WIL
VjUwJYs5t4n2JGYNe8aVbINFiLi55+SEiWWAEP6i15jftr4XS8midFPMKiTGaL3s
fK/4wdAzBUMMuX7zbR87FC98t7kpCP5lTB7tBLVFBDlijMVmWhQv4VMwDhFO7X2v
EREoY2cinppLnGrTJpl/CEcS5kof/+R8Sc4SCrSI5jAloUarPA1C6KdjkKLdR8kY
qMd+gDNzbNSy2UR/I2/hCZBBHPs0pog8gXB0qJcua5S+PathlcfnLSbzLakbWloO
/agBGWklOs+eYJGdlSBd3jIaPW3WxzRDEEo9bjIw8Jp8ihzCus8uvI9nBtTThc2b
slJGl47O7JqtTwISePUOPbwRviUZnjPgsNpnRhUn/M81V56L/V+hJR/gtPv/YaP7
hN5MNjUtHTCN9o3txZh/Fv3si+OzmGDrxvJeoA4WZIpllNflUZMr0ToEzLrmBld/
v0Qe71G4YT25IDMB5vTQ3EhBcjotIIKV0tNqxD4A1DBsBg1dEDXiL/QSuGq9mPiP
4zUcK8aq+sK2EckIshdt9er2kfId/YGYzEZa2vXZ+o34VSuNtvBQEDpl406+xrVy
AwnVTZsz6R7sgKPtTkTMyKbWgyQRDCMxTAw81feUYyI3BjCc9kuEUgQn7dXsO4kR
dwl6DSwHObGtG+GbzsBXx2o7TSGOay/vm0FukY76wZ5qBE5BwedvH23ivFSFJVzl
4TKWOpCNJ7nzTNy/wwepNLfcwHGmTWR26bMoG9uBaKsVDesu37ObTe8KXFSlrCvv
LVNS75tVezD+uBZrQDVz/vI+gyLvQwaXY6oVMJ05kMdmm/T+f4fPt3XwqbprLsU6
y87BRVWtl/szLTbgFyFn2e7Uef3kiV3jYbuecOKD7AJsmpnuU+3/nJ1/aU/G+nPY
fHSs26EfPtJUUj9Wwucjmluem/ZScF0tRbBB2DY6PcZ266UDdquGeFMonRlHOqs3
81+yuqKGdLRGVZpIrUb51w4KpLgl+8kXd0WDYlPWOk/TWqvVEaF42nzQFTWElJ9m
fEYTe3Vfrfsq3JqJc5eESOHywsORexiAK6pTbiLTY7UgAIIbhDNmOlSw8cJ2Gkmr
nI9RmDMEnZv+Qme9WC+x622+OTj8JCESeLHNYdzfs6MS4unFl0Wb+VyGAK+e7XmA
ctbBM8zxq7Ma6Wt0Y0YOyRH5KQhayx4+czwydh+urMNQzKoQSuJgOjapZ53MXoRr
ValcPbm8SibfT4qB5Fa954dMUUpBsUX115G3yhNZpxEdsMhF6Dkj21w1bVkO5Wjs
mIUTev3okC28bkXrscHIzlT65cFuLFfud71nYg/fs/WfNvmbb/ik5iG5azFOrJs0
zKki/dzJP5dgX26edX3q1ePIOBpiA+PN5D9FrIfd4vH3csxBMdivWkQyTvisZ/NL
R6RcelOuetIG40rpci6I80WSH/Fb/G582MSs/aQO7Uw7OMZLDajYUomgtqRE+CdR
eCf1e3ZRIrEcha6TkStn0gIE7Kd0CRxP0q3PhZG01sUwK5J18ue9Llf5cdv6+Rf2
dVnJP9Al1VbTpONDLh2LPc/ZDuHoFvpDobSYU7LKP6WnthQ3tSirekSWt6L7i0jV
F4OBzfuWbzB8wMn+3Qf3WQ0NO1y5sMvRbzIjlt10UlgEXNLJPnv80HajVtX3WENz
lQz+prnE3DKpQ6noVc0bg2j4JfN9uzZko8ytxjYw1UXlZXB4CxAJnlRM82TI1L/l
pRCNHEEplehG+MTbVgZZF7lakoQ3xZUSuCReSSWyzDOSxoNZqCSlrW82gOwjaBBp
BSzqrgjiV+oLSgDU6aMEwL/ET+NlhF7e3hIijBCGnTNqm3K6FqLdK9PMigVAJsWx
QsmOoey28IGRVD2qwCJ9sQsvLN9gpdvoNSPSM+IWM5XE7bnsXKr28Cz6Z96o3buw
F8hjnIRYq3G+fMXBtR+KizxRemX1Eq0C2YPEdadaQWRCZg6kN8z1SZM4v/zd2KoW
zMuBb/6SJ9zB54sTY9fGuHz1ft0pXzip33eaCeNOUB30lEDKXA18ARMJLliBoOxP
f/YYImV/AgLKpknkaxgOkzfzidZiuVeLEaOp2u6Mnn/ILEW2t5HMACqOwCCUh/vJ
OlfY8zz2mFka03Lt+Ms2oV6WBXxCt4oLzjat/XTmaMTqUqSuXq0hNMp4z6WeP8ZN
iNHKC84if8OpAzKkgOk03cW8djWyLpKl/4G8VylrmNB8YhczDN0DWcQiFtg0LpRX
wXXufZcwsX/Eq+s6EIunTJAR6paJerRjPmfhiAi0H7ceejYOlaxDfsSwSqcTJL1W
81hRueW2k1Ia2reoTsT3gqWUjE/qWpJ+pD6SZ6s5cvjOSbRCKCaKJFsUEJ1V2ru1
Yh7XOYXYw4oZJyXpf98PJsx91KecrL/nZK9J+sfw7vJvjkb+xiBSetWXYDK9uJnF
+7SgYlWeE9Y6Or8jgm65Abiz2R5AcSrrjpAnansQJ/Eqbkog/voifl53KCE4b0Fg
9BNJaFV8yTw+v2zHVdqCST3gW+l6IdDY8hMnsSPMKeaIb+7OMGOOdLqOIaurMJJk
X3fG7gcYN2kObyJyQUP78BHPAB5UyFSgGtPZ7bKE1p9WVYgiXOSygJLlOPCie6gf
iN9HNGKKFoF0WtWPyKMfUBaQor6MeDbD6j6saBQh5M+wx7LwO4G+YTl4u2ndxSlL
9+XWAWt7v7uhMCX+Q2ZCdveCPX1Nu0REEeMg2byGhgvo2wMDwwoMjlUj9D7LtFvB
K5+fzpBfj1xovbK/Kk6zqCNZBDcQtKq+Cfxk4m7x4GmPg1zKzxg1I0XF0V3QmKis
SamQfh6eEPK6aEr1otVoF22hIyvlo62/w1GMgVcByw14O8O2CpRNjzS20gfZXFrz
+R4EzUHMqfwVxgzokGH+Fl+d5IwIeokejbqeCjJRySjnCwMs9YkGzcHiWgoPh+e1
VAOnugFvd4DyV3Epar3UgEtRyU3Xuv6onR4WMrQCvdJ0C5Zj81TpJw+cU1qAi+Ru
e5+1enUNE3TeIeL4LQxM2eoA67jYhjSucri1m2BE9vnlwLn+TN42gCj9jB/fgJva
TWsHXNenaOaKLXzRwEFCW+lKTT0x2h0uJJrXYeB8c1CBNs9NNZzUXkBkUbpJFTmZ
NkIt5kEzm5qmkhUo7CPgrnwJY3g/LbZLu4izjzXseeUs5/hEk6Dm6FOqvktLVGli
bb+0JXBJIZrrlINJ1j3IjyLNHN1TJb8KV8XrA3pLobg7jICprINxkPugkcgCzlvr
MZMgzdrAdaKeem8BhpFRakvebvF1E5b1zYl1/0i1taGSBssWTaFLHjTRtb/EbmL7
4ljzN9sOWP2ust4QK656854us2IcGWK+nggiuUBS4OhNR4fxb3GwPu1iguZp1h1D
EVRy4eMNPB2wffzoKzG6+t9l2uxhcTvqeG5+tHhJ3z5PmhLd0NdUDL/gEp9EubfT
zSAYp/9SyVKqtGylFpXHXAnTcuWMsJ3Z19Kj8UN7AO7TeCbvdo6lByxwrMC2DA2i
WVarsTyh58e8gRjriptYWV3M72WR8/zr+ap/wZLEzqSeZxfNkl1ML7hRJlaLnyJD
R59GH67ZvcjAa+f3ICOHpOeKuzulfL3tF9ngvZ2+muEsE2y4tQzPvHiRCMknx1mo
pTFQ2BLKzXKsKbuPPbY23KXfAJ8ZMf/URIN8xh6L21+QqS7TZXx8aUfDTkLD/b9B
gyaul661uGUKVrVnAUN9MRI7zCsF3OZxOzAEAebBlBjVI78WtL/0UnXQ3ia0XrRZ
n5tzC7NT04m2Kqqiqq5TWjDL3zPUtGy9hYpIHRNblUppVbrmtEFlNiB8PzMMWovL
LLVUwoMpvOsHg7wu91fhZBnMAAzNfKHDkYYD1uCbTVEw8MvOSfkRIEgKxmfotldc
8zelCgrLGUfhDVi8dKiJXQ0I5rgwj5QEzV2elT+uVhyoUuaTTx8DjBATyIXZYQT8
FjQGXkf/eNn/fu8Hc/MH6xkFc04VffyCP+Hjb0URSdQQ5qGo84ipztgj2fnIoj+f
4ZM6Ka3njW/tVAngZ7XWs+KVbFlu6RNfb2JDDFWE093+IHkUP5fpjMHZJ+DLUTo/
nt4s/+gsR2D7M4LB01SldB8WzUjAMuIKFT8Gnv7gg+jJgGta5p1U4o+LE0bQx+JZ
fQ1NvNh0QxHjS8mn5yPKS5zAfQn42DWm+zWqkKSoagJvgI9d8uxlXVwR42UqhCd7
GG+E6rGU7+R5N5uhKCtYbC2S6mFlxCM76UqeHJtXaSUXXk1mQkKmSQrkCxRvx5Cd
4dioDHhtd4Zx5f69C6rMpynYL6xtjkfG3M2HEXz9b10q/ebE9kmcDYqsrXIdzjqA
Lja8goXBDJFA8prhxe1Em9Lh7iHkE4zDXMKBjp4OKBHWAUfcVuUwdbpiHk7R3TIB
tnTGGehB+iwmj0f9QtuRaNjKKLuOHRZjGTbE6Bw9uaax1cyFLj9c9muidsNChJHQ
AOAsaOrdp4/mX2F1D+a15tg9DlSmoKFkfE2UyeSrocCpPHL8Ed1GFPCD0NDip1R2
wheSSZwueqUNEf+PR9lLtDPDhg54Ag5fzABY3Uvy1+4h7BbgVlQ9TwlZ4+fj5cCQ
G/FuuaTWU5SubRSEK0+dKE+oVuvhE3Tkin11Y+qlNawAEz1iIKissHi+xSEzUzwB
UOtKnRDePO1gbPQucrr/c7XDIxkOQzmVHtfj590uPfhzUBvG5sipK4ZxXvla/gYy
cCGAAALXLze+NMvHhDaN4n7+Y/nJrS6Vp3JD9B1siabmdrNbI/DD3sofB2ZiEy4N
UYfHhSIQo/RGevnuRNCQHk1rQNtlmRZOMmQbGmT1XTjqg2bergETdRUT4H02bH2n
EAge/fwxPq9wjPk9jazWXcD+nScopKHVVqSsfDON5UblTXRl2SbYxslknTzuWWWk
ixyUO9b/v/001QFXH/w82EnZCW8RFoOtiK/azU+riVGrGXrqAk92bfyeIB+evuwX
my0IRt40/vA6mh0wt4KcLpnPN/BtLfp3jlShck0NAJlMvgtt2+Er1FqgP8Gp6g5r
2LSBZCe1H9hoVN6xJRDIWux1zACy4YTNsmqB0XBtZrNS026r1FEWuZQ8rl7FjM0p
YyI5iX5a183a8oGUV8f2YKXSydvrwtjZ3MdKJRNajP9Mtk4lRpcxK6MMtXwVvoD/
2E01NB+zpltHbJDS7ImULFZ/+0KfkH73MkuHrUAb4Ve/0NGdXJdQBJ4k/r+3bFgV
Gt7ZB8jnDErzU6Kl0Tdc38+xGA/rC6NYwU5RsSdnmcm2ceYMLiiVF1LK5kxAKX+R
stG7dy2kX27XxWOzWJqbGo6YVik3/m4oWt5pOzvZ+9uDW3cEpNYcZA6gmXUsmD2F
hnCT/7LDWycOtpkr0yhDH+ltC/+sTsetBol7v7R9WTSYwiegRgrfaxBz6+habZeM
2d30my4P1IElqeTfiSz+w1qDGys6kG7d4JJ9vTbTRaAlvt7B3OqJmKPyg2j2/itp
9im6Ubp2UfypORaQu9ffGwZObzEArCTzNQui3nsPPSKwILUkkGTFh78Zc/E3ObVj
bTOrvIZGaxAGIb/lWamB1ghkE3njAh9VlVzSAbzR7r6EESNJiuz73eqGNd36RVDd
8lZCVqWodJF63x9tKBA1xzwh9TMU4FZXWdkJApPINSv2oHrY5UY95J2HyVJWVtgC
vZpjFC626VxnC1LCK9c+yHOysgjB8VCBqoO+cWhFijSrEyVTymE9HQjdwFKpDldY
wdh/lX7Zhhi6SBaGuNV1WodrTQ22RyWdnsWNaOLZ0n4yODrHYmo6/ek8FchPl1aL
uVEQev++r4ZplrCtPmoRy2Ljel6imQ/XmrvqCsEXb5k7EHzRQEpmNHqQ+6JNAAxb
RTeHcl3m9zL4XDaG8Pyvh1Ap5p7FfkKbQqA+y7nNfzMrH9tEGRBrVmuIwhGagOqm
WF88gmzIOnflH0oul9Pw/OmIKjvTb9deWBnN7W14t9gMELusZVwKPHaXL/HDVYnC
5oZP6xDHmK7scLRZgUNiR1is6EFxK/7PGOYT+LnsOX3KGz+VW1A+XzbwHgldqaAX
PSJ6eo3ziqHjdBiwGMWRzJbvwfgfYTyjZpDSBVWXlYjKXIPIfqZpdNXF1dYrj7q4
/k5OznTdc2cM8ke7ZBUOXr4MT/8EqrnZxcxOLBoYpGt5eg40701iICP82dqLU3I6
u44fdZmGmufrlVtdutqm569ZrRYGm3CLaItDBoBHMgO/dokAOVxNHTABReXLBhVm
S49ggiR6TlDxHK/uSX2im7QunIeyzkcVzkM9BM8PWgKS350tTyCdEm8Vl5OTbFb+
EOJTHcOrvhUmNM0QUQFVuH6j3DhgGuZhnOzw7l1fFKDTNbXfeaCVDb54kaofxIzJ
xg+uum7p1TLViTAy7r04YKp7imnay8D9Z4oC//IxTyBY+tiaUqqmQ7qXdOXFB1pq
IFMJ1Eyf33IuFHu4Vz+MeBserIYckrUHfuPfGlTPUtmzoUm20WgpfqdWdzoSYp9h
JKCnof0F4l8juhwTNO4ehK1PvmVyppr2zDWoTkjxX3LMiZKapWEaGIAeXGwGg7Pc
d42uWczM2+m4Vyw3RD+bnFpECoGc3B3Yf91Ma2YQ41djmyN4mKUydAS6ZfA8CA+q
CmB3lxx2SQ4ik3rMkv2e1c5P2hxWWeAxSmLCTkieksqoSdEEjlnsjh/XTahZlIlm
Z+QFzNoRu+h1C4Ez3pDZ5lilxGX+OeZXecEG1ieKvUC+boZP8DXPkd5pL7jmT6e5
aa2F9rN35v1+7thbBtM0X927iqrZstEfk1mZiFfcGfEqpajIhmMuVdI1mXjkoDzf
XJJnFRys4kSYksu3ghUqH3NJXLIbAiZBZ3YBtwfVR+5L2FPhAFT7orrdA2RsisiA
+EJpij39nwFr0dxRidyG6yECbKpgPENGp5b5bCK+hWgTaLy0O/n8wWEtOCS6ezHE
oM5djodMRsgSrJp7YbngoeHQRzfzsdz0BNnCy5+x6kc2d2s5xY4tRRc/BPMEsry/
A3eaHWDvaX/KIqeZYjuBYd1fdZ0PZbtb7wm1SdyEuVl+WJAGSjXzzb/tgCIin2bW
vN8mFd5IC92MFnpcYQO5kQEp4Uv0khd7TMLf768ZPEfFlZO9vXAydJ8pLMbAEdRG
oxLItpz00QWpWHnFnLuHRo0zKtm+2dNkNB6SPgevjwhkioFuI5K4kv92V1tpbdom
fNWInkND0A3pISGJWAsYYv4vj1Siz+2mBtu2a4EGRCOJcr2YGa07x9WOqW0o0Uqs
4fkTAbj42Tr98sd26Ww8AeWfPVs2LSXYVo+MBbU6MAIOLOe9dfmxHf2vXPpx1MEi
`pragma protect end_protected
