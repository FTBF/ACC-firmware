// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 03:56:34 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pxoZpgoPHIcCM3JQ37L0X3pDa43jWsvvLxUlhfRFgYZrd8hSqzHICmo4AuBs+oaX
ENBeJ2t8BBRhUI1c1kRkYIRX24PvpFYF7lkcYZQzYHdatjjjgaZ+tMt+b3Yi3dc3
NxXlOVhvvPLTmTv/ec7KSdzzp24i3ezbgEu3Mg9gseA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 176768)
BCO02r9GwVojP+sNaQDGU/yQp0YYYfyW7CnBn42VhLj4QwQLE+FvqDV6bZ4u07Jw
DgJ1iBwaBK8hF2TunxWNNcl/riJ2JFrd5/TjgOiWd2w+ZDnfaWN0BBv7ZPArfofh
AzB8qP6eJBhOUBEhJm/2uRS1sNfFDH8ewpTNrlg4Dab3et5URtwqy7MjosdpNF5o
RMji7MeyOY8gYU5N7/fAqk3UhoWXzMla5ow80ySLKWvN2Tgf28mBAa5Fjv4tQmkc
lQ3I+rWk1Gcw4GhAh3v4muPVs33RvTDCIe7MawnEpcdrx4kZCpU7eSKqfw32PWly
ieHXsV296NHbyj2e89TbI5eKnECgSklbFS8Yt/i/99iqGzYfUBztf5wxLIIJhd+W
Ak9T3eBz9RTMmhgIP2PGblbE/AIX2ReXmQ8+qyPmbPiu+RbBXrqRb/g6g4PJ/ux+
Sekex5Kz1Urj7Vt2PBI6XOvLUHd2pCVYh0BtWJI3iH0maGHf8crwQvM5i/K2NxX6
ROHrKeZnruobpoD+Det8wDGn6f+qK6mC2lmtD0Z43Vt70cT1HTDfJXoTfhrdoBoX
rY/x2ZJf8J9055qxKwDtCzWKJxVu9nAcVfkzJ3l7gB4+FpNciheSyHGXuGC0zqbH
aNCXKLwnu3+7Si4xe5TG/zL9XLBSxbPv24EagfBD6aNrnmIV7M690ZBKRNisdALl
7JjzHuLj3jNPYrOm01tksRPwYvilpHfM3twu8EgUJ9qN4xjnqrfTJEDjj3j2yJp5
HK9/DLhS4yiDyLbvP8S0FD7+F/T/uBwz0hmPhW+bVwrALb5owAc6UiCYl30k0jWr
QmTjQK4XYh38eqnB+rHAegBOEpLMtgypWw5TWCSW1YR9olfNRnVJsAJJUKA2N3OD
kBwDC28yI4kE2wC/Bfzorr7Jf5x4s3d/ymf2tv9FFi9R/37EP5hJgWKtidslHYJX
OOMXUUaEMcisFUiEuHatKD+7pAtI4LtLujmgEmZksD+hchtd2Xcmde6JFCNPLVXk
DShOvxtn/77XdsVlRaPwsx2n2lWvWMM+r/RBSunCkwXe26t5ycdtldtS+CqM6fEF
58Pp+kPohGqIzy1lNS3GW6cOQykd36fZmUgs/NE+TNksllFiCcVeaJfgvlLBw5Dy
qr3EoHxF/Mf6hsZAAaddd9SjqeP/VmBhPAwbqDm6Jq6dRPAV6ExoBs7aX5yrodbh
a7ifE3UGOGcc/5v06Q4ld37RcoHjbuh4AlpjL9thoVpyG/2xi2ytLlRSayIrSb7u
FQ5ovMkyd7DyboO4YiooCcRXjWH/KuJ68vgwzeH7LMebrtwOHAlewIUAVNmzMam9
qMNHbS1jcgWUF8w0z5E8jDrrde3leO06fr4VuBx01YcuUiKGebmO+I62I4IECTZ2
DGdNdNzNS30a7EnEisYFr6XL3TlTSm/1Vie8hAYjXG/5L5P41AaOe2bzEc82Wv23
HQWw/ZbwunzNVuBizQzbcBNjSVkIeFpYTcPaopr26Y8TuQjMJXGovNgDUYAiTpx2
XG0WUNPr79MPsfLQPp2dyohiZWPROjDLHQCaD81yBUO3Mrl5ahFO4+oO1wPnUzU/
twCgf70hEV4dPrgTZqbQlu303gsRMpRRPY1ocMHWmJgLQzWnR7TunsW721fQ8Ema
RoECIFp/Bat6WvwKbwyzRrl6euFvEFYabzrH8LwuoP7fMlT/yz992WyA9jLdXOmE
cbqWMJ+BGqZw0W7G/es5odDJus/3Bu9INNakll4jPal16F0eGe5dAfs1npUw+mud
E7iA9zekRmh62hXzqNLqvEX52DWt9jpOQpRablD9WUKvZ6K/2zfmSPzW578/mFWP
VLdw7YBNK6uBG8TGu//hnHGOOO02Qdei59bJus1tvJ/SQK+1S6ZVsAwThs/5mj9D
wesL/cQP5SwA0Tra7smruvdIHRpQZe7anKGRFifnkmlP1YqWCKwLZgr7hkXkmDcv
9fbC3Q7m3PNdjNbc6EFygAsPvjfH0ZOKFxKiLH/gzkIOxXp/QsfTpQppgyNf/uxh
ut3sl9poU9/aLO9oUnBpQjsRC7pAMRt19QZPVhywEDM4NI+mdb2PNIilT+ZsOpQy
uuIHAfN4Y9dxKE33UPmMmLlR2NDJpX8BIylm8oDRV31S65AmwmQoIvKe5uQoyM6F
7AzCe6h4m9VYllSSxGxUxyGZdx0+7qvrotyJ8SpFfcyacYAuIauPOrLrbw9y4Ec5
I2RiFeutl3HT3CeavvIz1MB54T31eBO2/2ylRobVA8NjQV0kri1b4LEesEysb0lJ
1iXd+jI3M7UfXebWO4DjBZmoGmmTkUG4r20zAHY+Adu+drS7RzouXMrHtwY9ubiZ
Cvait4tR+63QixmEyEdMn+OBGLABloZWjN+dpRe1cPAxF7CkLijR0w6g0KHH6gB5
B7Vjg6WXiS2SJRx5E/uL0ULrm+7rXwOa0oIZ4dFIRIstRTV/LPGrmwA4rmlD9Xtd
V1QBkuNKQvpbXbD5XU9mS53qpQxY7nyPOo/rKjKn3+zfmzfFFDqX8IYwsTPhDKCN
7NHoEcVU2abCGUvO6Obm+ix+DuqSCV3+dQGz9PMdBE8avZY9Pcq/Ax/lxjKOPAXF
lpY3wnVtDfUHbrseM+osZD8uwqxgvuwfSM+NOMGWPn2MD+BxsQOZ+z8h7a1dkEg+
SaIaulfuCA4mfwAD3c/6N6IygnGHhCGi51VANGKiZ8P4OjaRayEvqMBqVQosRpoz
+y24wKxM3ioKjEx3v9zE4plB956/TRGPAWj57jcVF6sN+I796Mx6/sLyu279LG4Q
GFA96ABsnpFCSn9dPudIYT5RHPWD5GCpznX+IiAUzNDUBgmGjjkMFuyhMVX09oTv
EY2Lp8ly3d0yONKv2EoPkKYoeOJ6NMt1FveaAZhCLldGmiN2dMGK4bzqM3Qux4t5
qouHH1wbp8S0tOZz8LLnZmUrh8qNFPN+lrZJzk1OATbsDMRUlRL36wV4jiKxZ2OV
fZD7aEFo4eQ8X4+5gdHoP8+84E/sCbnUntLf4vN8W1LH5zQeAmX+4UZwtRG5BQTt
UqvO8rh+RYK6M5Dr44Ih/yY5jYcex3eTU2G14KcoMx59Qu8GmLVb4OBCUggM4p+Z
R/BYfbcynU0HC/UvScCcSwNH0FuIUrOGaT4yAZJrliD4JTpFWtPljL3phZdqT+ak
cjLNcdZV0lbp++oOeTxC+a4fOmXzX2xhftY3++B1uuqavpoqA+o4CzrWTpEyppQj
BQQe73oWAjdFbSKvk8lC5zOM8voFGED7JMtlmWx0tV0dk3b9xHpRlwFC07UdccWE
LfpP7TXoBqqpZpN+x43JFm2G8ooA3HerArrEpiA9zJUzo/UqVSY4BU9/oFnb3SG/
/7erD1S/STCpwEc/ewWk0rqDnsP9gRH5pN92dw81L63QfgFt8JzETsJBTSLFJOuU
zPXMEaDo67JLzmj4t6ci0jHgEsvAINa1EaeG3iQVXzrerfDZknty568gEkbT08IN
wNbtRkuTlPWhgMFI7ZVcRY/3YEoXB/cQZovHDYwEx+61REkfgIBi3eksSvtQ7XVZ
5C20UV7mm3V+Yt8mPaVHJRcVK/c/osbQO0cLFmOEeMGKLFdAleDvWrwOb5JaDJ6D
ApNQmXfl2qhuh/FAN4eRQ7a+jrNolvF4u4+RqOMqSJAZN6w6A8NEO2PwSVWMQNs5
1ynmniab7Yn9D6kpQfPZQIPP9IZsBXsC6S7egJ2msKqY/Cc3updwbNEJHG4DYDis
fjaeyv8dCet+ruVL+XzLGUQZPruISaiUmeSvJP8uhh/kTWP5vovtygkL2CTvXitY
Vj5EleMaeDUMvyFiZihjaqZbFHd/+rbKXIg26aLf7QP88teRCOUycGdIFkr5g4TM
AFpoYcdEQ2b684WId1DTW3lMMz+SwSw8csjNvZo161bbphPm9kXJ0WsxNlgqAgLo
29cQWwdnpB+0cCf2BE36JYwSFlgmGBjnTuEObxPwfd3onpMsY0BLc4bkU97+nezP
Q9rC0TO5hWIN7nEUcVPK3uHnsNGKiEAY1VRLjUrD7l9fDeXhgO2HmoQnS92qSk9Q
Y9tdCU7SUB9l4CnsLjz26gWRtSwK2rzphd0bU6qDGwIe8avur/W7SU64PrEATVhW
nyJKciiCoF0uv/KPik7QyinGSu+jeSleKdvfhJXdDGABJCNePtSYp8v9DwjTOtDU
5LG6DXZ8Te5b/KUSjCXZwN7BVmWstggUveLD468IQtt68NUSXM4FuoJOgprLeeLm
4Yh+2f6HafoGe/WSesgecfVeFzojQf/jQdO3wYRl4x1hmP30iIQB6bSLu+LUgErb
Jvsw5y5Jk+UfISf5EMn1p4kMSfgII3nezTwvFWnkpPvpejaXiFolBV/0doiMZ8b1
c0BzuBbiU13PQFd1Xhy4SIXIDymOGvg0q8++2EFzVqxmid7hO8ydpCNdVlcTBuKt
bafbOza0377S7/DZ7HoqQ6fqgowiMhEG0HbJkas7IIteZ1McY1O8dhcFtttEN7Rv
hmz8/uSXubfeowywFnKZGL9pUBrOIa1qxe7y67lfo5F0YeDf5GgYlPPSfxXebcC1
8HpYjPKjjJgvzMj9HlyOUwjxxAYw2UDwQuV1eJI2CR70/vMFmmcXztdEtWA+6FL8
z1dyWndDLtxLreo4T7YO1kGtGg/sEexGsKlwz+c5cgyH5ZClkBHlqSj8Kd0f2Vs3
AETiRmBln1hrJz+TlQpa/vs3zSNxQoRqAneFnoeTPX5N1wflnhAmI9URAa25NdtG
Kng9QDbGCHa6yI5w3WUw5X5I6f3e1p67SYK4LC4W0PlZ5Omjsu+gJF/L24oFmpWJ
pCyX2AcUTqZO3gPkrs3YoIBMDVDeNR61UJVXGvjNC3kRFwMvEhu6s3SDGRZ5ieYC
kWmzl6sKz0e1jFRV97RNgjovplDPvy+xZNMweYCmFpv4sNoi0zp/HRCHU5DR4++I
2whfDrqV9H4zC5kzGeKRkwXaDfYhyuONcONDyMP81sKfFpj+0BY+n2esDIAn22T/
xsZl7xKbvap64J0WyMFVu0wwNz2ji9hia0MKa2FrgWwvlbsgjKsiO1GAS+fRorXg
jpZuhx21ngiYAvegkaEt+B0mqeqxb5wvR2s7BfRS26M/mI+ue8ZgTTg7S7lOuYkq
gFZ4X4xAuszsvEOgAobc8NMnQyRSmX1niTdQ1odIvZ3rrUwpBO2b+GeN4pIoMxA5
8mhtr0JzZwXf5hLRLe1HrH9BeIL+mM6yLXPsMvQ89pzU/47MzgEX4JGThUj9eZEs
pMF6/lpOev2mXhh5ZE7Og7YpHKHntVGEYE8A8AxtXlmixl6WVu64Oxr+luDzU9MA
b1Ks6pQXtz0YpXUIW6XmW5iGFglbJWscQG/4ZkjiTFiz4TEP9istG0nQ5agDNBYQ
OL+zceNoKsvC9mmEeNOAtmhPNxNIz80KXU0F4aOkZIGVmtlIT/R1yWgnJm7itaIS
v4gBDDZB23Gb9l65xupxZkkno1TYn72ntlcIXCjXGEzrM/X4hjFZloTD4yqU5vT9
edkVWJYXfTpfTL7GuDCnCEmuZeOh0b/WkvjOoYhZJNP+JnxQpgdwqMVQ7Y3U9yrQ
zX7hBwPYs5L424rpxmetm9pC+zdFVcvV2nqDtDbmFQcd3kL+KoJf1QZfS5qdKJEU
+fDts+nfwoSGMWprmaxMYYVg6cUhhnnsnlIQ6pNSe8diwUFqGWHUPS8AgKbvjatN
+89JSvbmg+a6xyO7bv0UGWKX0Ibe8L8MlBfjJkD2aaPf4HnXEoDQ66j2Y71BhoqV
/tH+xyrzb2r3LPN7AKNiZ9j5HGx5dTufTGmsqd2WO7lTRUlqHnBlqMey4kb8C8LH
fAsfWTcqKnBLJ4wjs6CttJxiL9yCGZEGUsHy5VyO88smzkCHSuFYqCKBTqm7lu8X
qDT9abkUdEowWMDcJs/NjIf2p4FyU0YF0J9K0TaY0Ob9nEFsXpQbai23e/7q456Z
qyinla0B/dVkhBoSVLt4YRgss8Qsm/LOmbCZI0wIdg6rL1ZqPRDReivo2eGYmV/5
6sT+Rtgh8nyDkSFI7o/+Q1jXefLVU0VfRUpuNM3kzP3GPVhL77n2vAUVxRHoeLRS
O1Osxj84xc0ABeOYXn/a0nbBiGrBEORI61Kwss4JuWO9Fy9wKCWgaLU0kG4MrLZo
QbP43/QQzjhslwlCkxyC7m4KEwb6CQ32liJrs77Vsd4D7ob+hgzikYopA+ki/nBh
Pp5ukca/ehVLdGkLcahChc+AP1Joo9ys18MmcCywpdpJvd1xySiLk2AjSx0ZS6Hd
S1r7kndZiQbI7hVLiiRAo0NrNa/sk27Soj622odzaWDuoVfVFunj2+OAJamZArx3
hcFqo0f9chcD7j34KG8tX5aXJcYCj62Yz8WbVgD0YA1Rj3NwzEyd21QRdeH3GMVa
wHItKAuOEwBtgmW26uzMBU3RR6ST37u6t1FUPhO/lMXk1gVKUmRZeQvStYRbl6UM
R+zgmCVDlRIfDWoPZTwCWRqpfIOVcjMXw7TttkdLmjmU1ZT3GPhB7aLPJnlXzC49
HcvBnx50IijSvIsaHSR9QrqgvserYWgajK4GZ+g0sicStRdZ4r+/DKpC77n479xu
BPWA81Vq0RtfplJeBuUrZZ0IbILffuetvauBNY2PA69UfpQ6ErwYI0Z0Ee9vk+Gy
LHx49feEkLyKlC1STO7RGGi0KztVgM/rWsR0Ail7jfYvRGWlOObVAHYQ33dcVsQi
gNOZIZ9P3UCwnbnvppGnPhJkuQQ8NBNJjpDdfO7looMyM8yXWkqR62Vhg8jKY4e1
37gBSxBPi3XtBRlpbLEExlho83MwcD6nvvwntlCQmIlbZAgbYL+tXAXSRfUj1duL
5Vnc37srTibEB7rl35HBSndS37sy3nULUYe3i376EED1dUe96TmlW540UKgvvpON
OfkI11/Cnlxm4fGfa881Gd09NeTr9B5/HGtPpGUKU7KLH1iR6ztL+gMy2PVa66Km
IFJRQdzLvhHBIOqlwmjF+6iS22eUnb9V5VHhKWgtSrYCtOyJgn/yporKwiKMi1aX
qricyB0JnGf5phsK1CTYXNoNnVkkCgvd5fRZoXwkHZ3tTVrYCZv4TpJIzNG4QdtK
LRm8/EjRCniMPz8yKgKdoocqk3dZZoO7GNaTd2o219zk3qdbQF+6l4g1fSJLfgra
5e1qUgiIwpShXSwz3tKKvwivVyGtf9zllos+i6vv5wEBev8ZVmt3a/aueju1N8a5
KSpukemNdIkhbUtYsxAMPelpS2R4UPyA/fzBus4YVxVCYsGw0ygOt7JLjsDFK5eK
0Ui2IgvwAfl0YmMRcqOmA/5eAU46x2qOJ7s6esCgTXLDB+VSHguPxx/KgClwRTIk
EiDFZ3fmf3VlPI/cpeFBG52U+Uuzj5V00t2533uyDaUo8izx43+Pd6FvOV9Igiqd
ijyXKjtt79SrDqKWQ8iiYtqpZHN3tdfzIn1jJYlLZC3l8qf+/eDMrP6k1PKs/OiY
N3PtusO2O8dE/cgsPr/UbikxOJPuo4D0qdn7uBPDofhVOUDG2rOOYZV14AuJtarT
LHzF4Ty8xshIGz8E3/AwzrblWPeeAsqJqY7pTfeViUIx8tDaVNiTcuvbgTLFQldP
VdiL3Pn58+kyjyVUMjtgilY3flW+MU//Vt6+UI43b0KRBrQLz/cFEMXipVdYrH95
F1dU+M4PTzKtUZv0ctMZsdm/b7UsLrVyKBI1Gf/QM5EXCCsbTUgYAXi3Xj1kTlWg
kEIiFAAmWqxPaiPmEtdJ3CZv5jZWC/Gd86pAWc2O0miCmQQtZxGWaJIT+wSHPXQ/
BrxQAXmmDUw5ayQLqhavHh+KI7BitDsPHpVmx0GvrrFxdNt4RYdBx3KRQwNfb5DE
FuMtnr2wgMX5K3v/261B7legqqJPnQ/eXVsLwxIpLtSykV3HztcGsvEuDApQqnJT
PZeP0dle4pUcSutiK0RMy4t7WpBKpLssy0+tB3rZsfjcck0ip/0zGaYDa3qRYjdl
ODowfjO7u4lS/P6KTc3v2OcZb8nSKgy6UQ7NrLtWwgalgWmSmIPnLktUwKA7YWko
Tgl3j0eKzqXFVUGgIjoz+gmly/MI/8JgTgmZcBZHpnZgkJ4UkdZF4T7wfosGqFWR
jM704fsAT2jJcoM3eoPMvXtKa3bs6p+0Bwyxi8zZ2d/s+JblNeoFJRVK2eUbRoq9
NLYon2supZF8P+NLsNlebatqGhDF94IBkRAQP+EMcKepWHMji2WHJzdXzTvbtAP9
tB1SBUTWxf3eRd6ijv7RIQnzejlKK/LxtJJ7cben4h2RMnkebQlrEb7k12R5cA4B
eXo9n88h6M8sgd0dddXbckJeXayD4KxnoWE0Ncw8ZPFoAkm3RKatjmpv2EJDWN3U
5Pt/EusknB2AWDAfPbOu1/EbUxrNYrZXw8kkjp4kcqvigmLTU0qbr/EExpY7NOuy
cmbnsQDLKw17P6jkbORkwC3lIUv2VMrWdt7Wd7KmBYsvyNUOsQXOBO2XdS6SLwil
TfVK3Ve6SrMrsMd4ps1qMwOac2yjO8j00bgSFrt6RAKmvOkOKRNHNQGJGhB6uX4P
K63yXzJ/nBwbx7uAkdJoyB++ULBl8OSgmuPh7WXKlBGk1lPzMBKFTMnt6z6Bmzqg
q4QrfIX3xeAABBNcZxkugjsakqxwFa8CrouiOFuFByrADzUBvlUfG7La/WF06RnL
83+cnMzbmDAtivLZPqxLlPkAbfZaVwVCXH8ak/D5GvKAUtF5jAozxwPJpmaykwLr
QCNsNmGYoPbUB8FzymkQORmicORpHfEoSNYDWPJwvptIMUyjS4088VbzyBhIvvfp
sppErmpQV2Db6F+EKC17W9bmx4rTUnQhLSuV3VAxBP7G0mo77pXXM4PDHREj9I/V
ai1imqGQmN1GGVFkx0AuXLFIVfRSfFWDrQlA/7OsfIZmxUmDE7aPMSXH/ZtqqqV9
nU4XxEcGMAz9dYLYhonVB0owQhiqIfAaUvyWhjMrgkrJlmqZplS191MmN/1slHh9
xmCT3iXkBgQn4ADiJd5ssnk+ff9Syyos0xtDVy0U0lb19vrWn8jsYoQqBBjCGSUe
y998SlpDIcYqrSpR3QhhpB16yFHxn0ZmP23kWHdcgcSx1WSDC8S9R5J9gt0WavW2
MdfKMKt87lUj2br672NTckUy4wFXPAsPyHF+ohUZ2zjRzfYuurRzm9BUkmPXUnxL
Uxn1HjzmHEYj/nWA53k2vo9erQS5PwrCCeFZlbv8hZYR4iNTdW1CzlGPWeKGQSnA
8mr4to5sXFTwDe8xIW7OmIbKw1gUWvn25TKqsadg4UwmPkuAmgyrDw+j0Cickk1q
4fmraXCYPGp61LJRnjZgFvItjdp/fujAqvK+AHtz+4Tl/tOIJqwGjTb4jG/p2epV
bYvNfl6RXpmaB1KdFieepekOpHNigDb/8Jvd0HNI0bDueuvamF0qF8Qmp0Q+64eH
dJIHdfvLj4kLBNuxLgpGkh6ye/ts9EnMYgPRO021S+8W55CjD7phMpGVacYkk3HB
2P0CPkjufCdPzJsfvsCNqGhY93x6EGWfivTfzX8b6q5DYiBeLOAq1kz+5X03ntMt
13qL5jWdi5RstbeT23VdNYAjHjuFMvfoP7ASzJqki4Z/yQyjZWGTUrTAPr64BZ2A
zZnjbpnObl0k8UyQS3+vw3W+2DiMXWAPXXGjJpjQOejvEgXMPnWBx3pd6tdMcg3W
CjPedn5OzRyfc5cyshh7zLDCNKMESDGBqLzomTJsE/AvMaYbBdZaaWrE/nh06Ifv
+qRCY9Gk0LYQKVy9FuhTaIaIJ36+qK1ZEZHt8zrycKUg8JWSnYP7gk3Wdd2VfQGk
KvXyYkec3TEgyjGf8CxYFxRE6ifUx2UvbooEQ4cdFZXfSeWz1E1J0Bgod4WPTXMa
ObF/i7SsXn9PaPN2ih/9ALvqMt/QR7uIrrLx/8nvdK5/+mM1tAnLdJf4tBO3Ji8g
F9vj4I9TPDWRQ+nYCc8tWRWkzRty8TIl4SnXK0eOvvMWCw+LaMJLUKr/PAG2QPWA
JrSlDKTUYaAF/5b3YABg8wmWUFRIaZ66AcD7kJ0Gi0TSY2Smm8oE8Qe+WokYP07V
1ubB6HncBckEeQOn9CPUdQdXpUuwd8lsM4kjwxbxmDRvET11A63MyC3JUTTzd6wX
TXNUfOrvfx/IHjAAtcLq0D7Uze88VbKzu6Qt+0DXFCAx4RJMPnYJ2ATm+gkaxbqo
APXBGSJYXRHp97uohfNfYOBy3HzJzEYKRir5+JFQGtc1A4/KLJHVtkqCpGVC5UoI
5gqZEqY4xdu6MXwJFNeyTT14cAqTstmbqggMECVw+PiZvxNaZpEMFCu4Bv1Ichue
obx60EZoIZriTCyZnrN2iGQWG4cFe0E8PFQ7r64KITt4QI5YqJTVsXewmRHlaoa+
JNm1oTeY3o82hEM3ielAGHk5xAS4obthM4svi3qwY+2GQXf6kIHXDFZzEt6ZxKXP
o4zGrBe/v86+KfPGuj/kzR5tqt/vv4WRWxscj8Pb+TBTsvWi6zPNgX05cIztTx8K
dXqK/PfZ+MR8qkY4wNjNW1mXSDo6V2oUycBpDzq114Xfdosf8HdRhH/cE4M9bGOb
KbjXeMIjfSaQgNwSJePbicly9gRVT4GeYnbxotVmyQYI5yF5cZnayuwNF5ro4uOd
UtchS9iTOJHrclrgJUo6i9yMea3xbrNjZFw9U04bA8aFsmooc4Lxh69VehKU5uhQ
294i0R8a+zDv4ke1fE4iLWZYgzHQXPyhHbAsRKdfpbWHbncB25yMvO8y0Fx4bKBC
xyiO/giXS7SByO+5p5nTS2+vbXI/PNMPVe6/KiOv62JFdf+a93EXstgsnxv9ZGkd
zvIdcQ6lXVArRwdou+/kVsi50Qlm6a92X8309rupdWbGoqEIwwmt+/8jcxm/iM8S
j5sTGoaICZEk0EBbqeAqhTPNjhhca/t6E3T+XDce8G+dNyc9kWpcuk3aCg/uxzux
ybHaxYB/M2sSIV87bVnJ6URfJxXWdZse0IKm3QgAst0sDCoQMb5cp2KuVcw2hTWa
0pAe0J4DxLZ/qlxDetONf6scz7LzkOOwLsBNkjtZsdxf75IKpdyUPhwmp0CLkUQk
WW3V3QJkd7mKT4WNggeuMmgCkSqVfOYLglEkjH/Y7ap/lxHrIQ9HKmzlqYrOeJHp
WU8H5ntvaslole+M17oPlToSs/wLEL9KXCYaH86q6KRY6lF0zLfARpM3dO8Zua1p
ejrziHNyN3ncOaUnecOemaTAeFuQxyKtMCXJkaZIS/HWtuUSo63Yep8T++1EBF2G
8W++0LnOD4Z7AO/UclK18DdQVy/9FyhWKfL5ivg7ezo5bQ/mT0cZ/3SX35JZNbDr
VpS1JNvA0oUx6awMGv23YTbD1S8yYWRfeOAM/Wm4BtbbZXgjCabFPtYvt7sEVsUK
AoJU5KxiSX3Q4fiYLfbvxhdOvQFaBG8jk+2RpPXoUCVL8yIXk2b1QLIvd1U1/2nc
aGX+l0a+4OWZrSC7H5nqpv/Jz03abRiYPTlFVLoVPYEOxVF6jBYbko/j45HzZ60m
rc9LthanRUnjxlSo52HDl0jCTbpztQzDGaGRsGe46bJ5mi2+wQEeRw50vCeakyVv
ZKAk5DIpkIRGxnIyHFUIOyP/oQ9wL4enRPwE3WaNdYGVo40ybVVwSt5+D9FHLhds
+sbrssLii3nGQT4tj9/kgGieTkexbLg+CxRmD9DgNdWGd/pTK3p6DIJOa46mDePL
qvl0wWOwdMxJETePJmsPF6BAJRuWq1+PKiH4qHhlnWJylCM6B0GU8ygmDVEUspVt
al1KnNplCvrsFOVYsE+blJPXfHRg1Ywt+5g5mYZj9brLYPXoAI/hN8CaPcKQCI2K
RpwJDpiaTyekh+S+uGOVHVe7XNp1EVMRcPp35nRg2AHO6bkVmczzs6r/wZgizD1o
gj14oC4BC3meliUTREj3CPHPk0kj/wh0jU7zAsacTBjQaZbh3wJVSdS7GOmInZGw
OkT8+TkSF+Y0pXlpiQAjqbZtg9KI591HqQ+7jooe5l1WxKfadvI0pkI0d30kLpCw
jTxTH9FdEgleSuasT9M32z8Ac9J0NTZ/NEyMY9TaoKNwxqt0tG9ngkxw56TtZUCe
FJjaIsgyu+TkX1JeEzLSkC7b5gz22IzdQ/ei4x5uksPQCIUHevDVNAHdiOVuUJ0a
+3djEtltrQ4b2oYbyACEa2NqIIu0uEclFteLp8RJ+OSlBabagKQKEnGdhUYGKqHa
Xt8CT60gfXFtpWNcbjkVuclmA5OAwm5We5UVkPOjV24WgVKacfE4hi9urhRzjK9E
efBAt8GQ3VxWcwyvVstk7jvjvwQqCjoOeB/mRrOG+VfMb9o4ZRTN2nfT7bjuqjx6
pRZ+zTnPqsSNRj7FoHmsbqSBh1vYtTYcP560oFT6ffxTKAY5w6yX0XBWEpXGvMTX
rBHBZT0kFNXuWjQZuSyjGFVHedAkErCdRadh2T9Z/78mcsMKM+05vKStmJ31cir3
jcrVn2/mVkzm4YA5HCdIGIPcAwi8/P58hlEJDI7xhDTxgCi63VPrZEiR2TXlFH41
1aQlY0ctlYB2XlWfD0AyH7dXGkK/DTWExQW+QIXwJB1wdHAccyLra5H8PdFR94al
CQgGt0AlOOJRiDlvhhI4ev/lGz5n+Yd7Uqp4GY3OVZvRvZvkKXe3zGhPo8r3C/Ji
30jjzLvD8IoYFTfE+tYHmgZvazboOaTd+tHFQtEKTUmP6bTaL4Tpm1mQJAtsHLpc
+2qGOWtHH1ByZPd8uM6Fr8QvAH2vnF4Zkn1nJuGfBOQDhribUxE/D8R0gXLY/YAi
axxxgHGrzoGpFaD2WKakuzKLQ+REk+GuP5O/D2vBObxz17SRC2CPH8yIFc4ndlgN
CGMkq7ZRxVVllcWvcQhELjBRdBNF2yqgXGFfuF0ncltMjXNNw0RhhWzD/HV3n08e
CPyKasDlCHISxbykGVFqWESNO544I0IvMr2TzWTbVzRwRh4VG+yDyBwCWaplDMMC
kqRQ+8nYExmjvXdTNClRyDA81xNtgxjce3ij8GkhxoxIA6J4w0raTSy9CGmTHPx2
bGtsxUk8yq1XcYbHOSYaYuIF+5iFBI20AiDHxIz0pZEjU/gu9bKP8ArZsQP/p/0r
bGEsYN0SaWap2fvnh/90etckyEXCbvtwo8rz3T6C2j1Wspy3vzZxQPMDVySpA6W9
l6kL1GzTU8jovKPkNNL6lKSGm1W7uPeVPFn7t2LuPiaABTCKOVu5Tabjwzc8KV1g
XlPrJD3VbUq+X0gwEhMiSLnX3LwYi3Ue4kCxhpY24Q2+TUiAtdlAmmkbhFsCxhCP
H8L7cSm2LL0xtvR5XNEazaNQaoWlxZdrGy2dN9eHLmxKBOJHSoRW5+2a4ynY3QVg
bOZYEbhn68nX2tMEKiwORsofOTU/FILnPfeq67DBygmuKeZKQGoWkQY08mJoB+Sr
hqAhD/2LSguc688piHLKKvgTQ/64gJ1+1Uds6A8+rMIbFeH27kDz3dwxslymCFqm
2m2lpk3CrPfplMJNXRVj13kqJM5c0pphCw60j+AnytnVl/OFo49bdDwq8o8Zl2Kn
ySn64RcDWvkXXN2q6CV/KNkDR0amknhgzGoqY7BBDcXDNuVp9QF5uYZKC3R9QNdF
PouyAB2YQJ40iaqTiXtnwSxR3VydBN49fjACKSuI7X6RxepcNBwuv6kC0uUvjuMN
xFgCKmeU3axrgdFuiBjVGHDOGh5ECZPzkUj0oFuzlZ9vsdLL1ilIjuMpCjMedcZm
x74bSFHUoaNB9W0OZZgXKWiMnjyHJ/CEoCsyA8WpTSrEpC40MOY12mk9q9wZ76PU
9e835bxLr1lR9gxUDdnytet1InF/5AQVelHDSmBCNNuN9PqaBa+N1S9gd4m2kfXj
rRuSPeZblDLNp8J8mqQKqfRDAZQYk+lgCu38i6+41xouyIcFa5t6phucbsUCNhn8
pKK0UuRLtq4/R5AQkWva5fKHk0UG1kJUHkLyRKZszokgy6r06hEf8/Sc3J0bvpcy
TxbNbZRaa6KdJyfQ8SzfVn2rJKgaSsbrPCEMaqetQGsQj9QARyaJ1TbAJG+A0vqA
kEjDTXZWdOaQlV3vtbFGItNuuT456coj8vQgretd7xengTdVn9acIX7IX7TqvKF4
R1luSjqiNg3ch1zdLNZEJtuhY6LSdFlxALUEjg9mB1CbYFELzo78ML4+2fiT2vT5
4fp4tMpFK+OILDp4WQe6Q0XwAk3Y28S/yPuDde2N5dQb5qYDpq4Xmw1HgAOfMM1y
rUJXLleNhgrmQT1nysLUrQbKG8bXbEw3CSxfEo7a/9dg0u+f5joztcFOvmREBUVU
nQgaqrKUvZ2YJmv7shZqkEuET83EO1UvlpZji4T47qDVsxv7pjDeImg+JnHfw6k2
NAgZw4c3E0ViZ2IMR87SnFvQFw/YfKlQxm16VBsBhgtDnTALsFX0Daz7qrG1BS5h
XvrnaEvV39GyN8zMDfWF3suo8j+b3Zeg5h1nCuqrC6w5xPjipyLRYemTsp0qjrgZ
B9Z/p7DY1EvkRXOQZ5pd7el6dauH9okGW8C3fTNGlY9Dfn+OSxGJwRKgrZI+lSBY
C5mWppME6RM+10evn2KN6rtmRPOSP2OGCe5/f+VieLVgXSU3RWzvzzLbOKS6RPBK
SxlPuYD6a3y/5RkSF4ZSAY0QUaqCfSWAWjgAS2zuGrkGe9a9chRkbudu9pUA0ncu
NpwsR2RhPQz1cgT4hREL3ORJYaaaoB6vPrP8US+C2NCsCTdZIwuZsT7ZTDPclK3A
SlcS8Tf/HmUebdijoKR8EJ3dqqlZXEg3ujdObz4JOpc1i8RNChkPzbHnpGsaP6Mv
PXIVoKWn2fX7e0/Rt99PjWkW5VEa6fA+sOZJNgTTqAE/ZyRfst5SnvzgRyJiCJBy
iL/5DFRA8t7fA/7ckYT3TzSxXQk5R7+mGkcwwOg4G7G34I4mLabAb1NhggkF99mv
4GtEJHlUBfNT3vX9PAmrooWy+ZzIwBwJc4MShClaJkZuLaaSCKkr9PBCBmD3viD4
i7d3YqDv8YGt4NzkYrStcGtglpR4pVqWLMIW5LviUp22Lh2hRH4W5mL2vwmQfO16
MJL2y67L3dRAk0j35bLidI51R835wnNHkYGuRqvHcwrfBdBkSsXPdOKdlZ24l8Fv
kvteEur67DdfXZVxsrE7PaDBvDyt1wZ12C49nzqE4dAN74gnkcG+S1KS6IyDxCeY
8jcyczXf6AgJAXrLV329C8tsy37BOzL68FvXJLNBJsqGGmMj7fT9biE+AG762NhZ
cioxR4TyirNL4jaCNt/gBlwi5RQyaKAbC09Kk9ifqYrwGQdHCAAsq+15VurmKL59
Y2UiZnBPuYLuAacB1EaJfxbEbM10iJ27J8v5VmWZAd+UM7QjnO3Kk7cIifn7Gpir
ZpI9JhvIKGmpnHOmt6K19Le59nbF0MHNCeF9JGMdH2TqiJqrVsU38mc+JqqhEj+z
7uBbeeif9sMZMLn77Nr28kQ//zg6dtKR9hdMYfvThrsIL4K9fu+y5/tZrcjw3QIM
chqdi/SlLB3I9T6EnpXoFAa1eRYj3M968e3DPAcusfCTPnywvooWcz3skqEuVQ7+
1t9YTlayFVSRIsY5ZFPTXP3mPZNNtMMaRgSJUU2mjQOEdcEgvVyvRcIGJlVCyRAX
yA9b72nZQVPT3ZIySrYqaF/hnL9sTWJjPacyACnVOdnZgqSB2ongyqZ43tZSt2SK
cNAgwJzePof2BkbjUn7b20dywAHhmqoJYPZilByewfSWkJvUMouKTLLO64i2XwAI
TAGZfJ9fYvGmdTAYUq9fE3/MgaHcM8DKK9eG9Bym+yEL3JxUdb7XH59bz6r5O6PE
Qc3by0PJ6htxgL76oeiCMKMwDx+JWAFondhaIxSgmmramh3HqscLhPhyS6IQkYBk
s+vjkPljR0buvfQ/Y+RJ2Yraz6sIshW/0TxsYHURgFEO8wjhxGf8HzjSvdQ3t5Qg
C8Q5uBpSswp/foNA73lxvlxy76qROHz87HD3JSf8kBUdPF6/06cjYqGVt8KyOPMH
+9EJ6nnNzmYv/v3HfTiUiJCY/PFXbwI+1ZWTlXdJ64S30/4jRn0qdl/1nV6kiB6a
Bi3xZmCx3n/jLM8jVcu3rXWoU5nfuQ1bvHfucQpyTObi27fYyXJBkCnkhCJyhkk0
P0RyOecOP7kIgqBL2KS6Mjs5G+S6txVDbGAkZ+OZVo7i3q3e9nKlng3Gud/nA22m
Lfg5lAqzR4Rl1qEqjw06e+8EhU1g5caY94GapPoWXpyhgeWssmwF477j2gRVueTf
36WqdvFwhQr4WjQNPYkDr7146fvrBUuCkbhit53CTUhVIAM5FYWxWQGWjCV57EnB
AH9R/acLAuBVWp8bjV56nfpma96aVY1N3qioTqJES4RcZZgY02AjFplRF1dVMQKl
G79MXPqBkl06EuXbEtYwPTpnqJgonD0tKHx6YZHOvTiqNTFr9ljHz3Z9Ikg3Drwk
xNtc1/b9jtgjC1rEY91U54luq2tsRQNwXZwr55gWwT4NvXXMxftC1n7Rs+IQX6sl
RzswKhoFiwrpoW8R6n79OZ8p2ln6/N3oatt5bYXL3BQplZPXnhLfdn+Lq0CAmHLq
kXLRJ9uXbW6+Yhl5q7+r37yb+HNhh6Oo/L9KU9ztL8Ep5vxqXdydKDJqfpoWW9nZ
bI5cM+zGCRKCJsHgD0jvMOJW8tJbvkGfjnrSn4BITq1bvK8EjytlZnL/ta2A00gM
MYE8kpdLH/xmDlRB1p/A2c2ql+rz2PEmIsHf9tOpl2t+39/UuC3v+/isLhcYCrlX
a32lP5v23/Q66HQ7dIq+xWxPDqHqhTiRaZyZwt/cI40lBixKUkjYTzHMfqw1qHdn
CFueYGeWPiDD0TzLEb9V3w+9BXjle40nee0ydZXeGY+K8ODGS3q7MV28tM9hoGmy
LU+PsnvvF3tkP9OtRwQ/rR4PIe7NJetNoYQDarFzmDwHv9Rn3Khb6WaIJad7H/3x
CpZ4IHHgin0rBH8qyVYD6eNjm2P2Zrg0oGdPFOk19C6VeObAzGaxVfaB6/UzNijj
Abw9UfgYKeB+r7GmRkx7KfJFynfkvYR+MkydNHZVk0rjkeHK+qmHOgR2VGa2fEP8
UBxIl2pOs03TcnFFqEzUsZbnhx2qEx2L4zIiX6itxBtZV4mYcjMW6fiV5VCBzzHb
oIDQfeXOjmpkjLTe38W2pHXkjnEYbTz0uAH8hMVuHUtMN9OPpI319ZO/e+eLPcwD
WlZXIl5soLVbAoU5yUWbBD+3A0ipGL6lkR1/xRn3uGy91vhEK5MwnzhhK/OuV+nM
BI2S129bpnfBl5atmI5ULS2GMYotvOveUzCYOlFX/SV5jEUK/xIBRBCBr7D04Q+H
gEC4zAj3Mbb/quze86e616FZ6plNCTq65aG/iBCkEBOPRE02zZkBwfOfI5EaSrvz
hA/yORuTrMti3rlWWupTNveRM0GL8eZEB3c9j/674ivrBJ9/l1xh7OUpCOXZtLkp
w3yeMFHedjxejD5gifx3I5NtDqCWnwA1GYoSgf5UHNeIASYG43yCvgZ0mAhw4BPK
H4YyKOayqBUqJMzIxokAwUn/G7TgqwxCKzWYr4b//bMn6QOWYqB1ikYGIpk2WBL0
iG8HXN51UFVYiL0HowD/y0OpHmLrjgwx2Jdm6E7Ip3Wpx2uY3hE3BTBmAqSVp4Ez
jCmG/F0i4riw4uaKj0wsAhVCuEbhz5MfoNj7zbJl5iRx5lwEmbBLl9egGokzha7P
CVQl/qIAoun5qTA86bPLws2j2r0HpUPIs9GP/pJiA26W8bCC2SwyiqhufXihMVsQ
fh9k9hz5hBMw122EPjkexpm0y4z+bKJQz3ut+x5MGxjTp6ToM6lpwiTXwlXdkH+p
8i666XsiVW/LRGlVLGIsdFRVftuiuadGVnwTNMf1JOMalZjKQs1h678v1HZRCTGK
gtnQAXjZeMmutOt86QJZ8b3L8pc7mttOpbYg4rQ0lPFNiAzIrD+8aiMDcR8nGzZ9
pxI3SptZPDzIFl7l95zk2rNZnoA3Zp1OOd29JyaFbLNrmhv9VWdEfPy+ufCGSanL
g4VKmfgcz8Azt0jbg4iDyX+DQ7C/FLToHjiCZuGkMN6FognyEYh6NoQ4cISVZKAn
ymk7cPp21j6SiokXH9ymkY+752ndxJXJ5YGGzOQay1XlZ3F8td52a6vz2opUdPQ4
qQEIsj//P1ow9OU8fmPDgMdNMxyY/8JyJ0EH7mh60/GAk0X84EGyiaRUZgUh6HkN
ysAqHO+wvYCSOZ7K2MHqRkwEwfrkP1LEg/S5AIUW+iOIH54tRmBwa62g7/pxeyVK
VKvdM4tO1m7c4iUIwRM53084Z4B+sVco2Lb+ThEKkrySrr1AwNQusVyTlHM0LbOH
Yy2tp6Rl7FQIqqNDK2pr4FYr1OhPXSxgseRI1GoS/Jf2JiwROcEiX9B0yqyBeFqN
5mxfFM/Bygk6TtrZ/XZDTweOvRlWP6eKMgan41c6XUMe6rVEGLi/xiy3T7UbLRaG
qHFM/rWfX+5PjBwltRCr1K27lJtt7k910L+OoDgdYQ/psFY1c9h1rT+XLNpynb1e
tNmkXpBo1fi9j5W3wHL5xWAns+YYQj+i+B01G/85ou3jO4Syd6C+h2nV2WFfOd/f
dNjOU4c6otj0zfM26OMWU7dS/OwqypLwEKDAbaFLOSbQjGKorzcriiGPwZ5bYStB
w6CeHRpkArenEine7Sujx8Orx0RxOF1e+I5mTgSKQp4iUK7WO+CbRepfVv60x5OX
jy0o4Q5NlPH/4IOsqM6EL3lY98smKImpl7EHS30/ZraCJ7Y0kNUQRUo1NsROPKSG
pSzgUD1spua/pnujJ332EKcM+fykWgL1rh7HcDd5h+zDiSNzF9nImUXyp1Ebj8RO
zR5Ns8Kr4kiQatnQLdZJTggPnvChh4MUYa6d4GNZxZkpfFdmt/8J2423OJcneXHn
EHUxekqU313hqen7Z39gGLlwFfgszhZCrC2r6D+EU6lTfCaT1P9cX+l+gJGH9AV1
KsaXt0u7RgvBp/txrylQrScXzPX/CpKT6NFL5jmoQhb5MciWz8ZZNsCvjOl/sbd7
x7jahkelOebnIrM8yOsP/TxT3xH2T4+AVtX2CI2U0uhyNzBtnPjLe2vfHBdGQV1i
Jd4AS9Hwv0V6pNogAYSGUTkJQ9Zn1q4V6slhE7DYgNzBy54WlwfNghn3Osha0uFn
LoYnBFwi7+tbnjdUWgjBux09ivwgC8ljKqoXNgXxWsoKjHS0cE7CTBbbrFkZaZtl
PDInMc2PVmMW7VmWdpMK2KaPAT7zCfMXf2yJUt5UgKN3FfxJsDBXyT1YuExbLTgs
WE0d9ZIdh4bu+dQSBtgOAFdD8EkUBw+Cq1W3IvsCOnW6xJqBNT718zba+uxr9Hw9
XNSzv1u1ab0PtdS+4McYj6VjCDwQXnftV32r4MzCOOafQ7gnAMVUxUAG0ab27Jyi
y/DQQ3R/ZZRyyBN/ot/CYYdvBh/quAkh4tZ0GjCAaG2+kFZ5qlpUGhvRAWQMs8n8
KMX4E2ArlzUFj9EgstZ/Ed46Zs90M98NNiE0aBbhjU/5kmFUfgAwBVFidEZM8Fsg
A20YmXHkG4BXlIePih68Cwd/TVhthAxMXOM2Bpa9LreEevopNwCzP9ub2iwFGBIQ
T0syyBtjAWVEQzwnVfagCUnMzHu/58x797pJbrgLCWWJ1vlZRGy5NKu5caQdO3rC
flVq++gcshTMdwxQyRJTSgN2CkSJVbwH50NtZyvV/Ed8D9ako7dftlCZNpsYutKX
3xadCDqRvvOt6tSqGYeczLDGClZsPim77EzcrLSS7Wve7Xth8f14YtpUJ6B+Dncl
NwtWn48JoHXOjlIleq+kP9fI2yDXC1yKILJVBfmrN4BtUnGILr2YGRIN2aOjMUhr
vRF78iLtb5dEO76rJBn6MBJG8LiezPJ9AZIBz0G+GuD0nIGBo27dQTTmwys/l8Kc
55Z9WtyPvBmaN94T4cNSiXFieBYf+meECTI8iUYeSmqwtlfn+GavF4HDGMHibz/3
0pCbRKsQCj6pUMX1sx9UFmPgTppFofIi6WX14xWr+sjtQpXs8cj0vaCMgkyRPWbo
XIxyNlelNiYjFEVHJvIdZEqvSzJZN8kgy3h5AS3rGWFkbLTbVQOoNokp9EjdpktB
twtgs3F3532VclcB+YVzb+mdPufMkZRXVm7/yUcdgoCe6/fGJceOr351xfkYhVt7
v8jNwn02bms3n0nO6AWjdG10Cg9iUONtfKdXoPc50grXO2Bwv3AU/BIQODLf8tPB
uwlJntCA3gEL4ZtOFb/AO9OVlhpPvBHy6zM9hz02YT38P1fp1AzWJvHB8Lsningd
/NJDF2MWGUR6bTKd8QwT8PTM4kQvAu5eYegMsKvJEuDS6LFqBuu2d+AQr/pZJ+TN
7Cz/zb1PTOxo39uFc1LMd7DmKxYQgWIml7OQ17xNzkN628sQ+QkdpzrYQlH9K5Lo
UEoE4mPlBqNMqVKDdAZs4FHh8Gdu/dILuL8Np9XWfWyPlv932pDv8D15GHlZDYGo
XOqFqBjlweQpVENs799m4TQ6zV0TLHkPNSHeiVp0eRG54M0TDe632kI6CHlw2LNT
K9qjYHg0AD9bEl19EDIrnkE3KoNWo61gq69FQat5wml1tkiSNQYpNe3B4qZs5mfb
hDjzhOdzjNoQdX+pFQsFbkqxOiGTAfiRlThWGBRvcHBwUJvnp9FK73STsFkYTh+Y
rCsOh++WSfRQHNPbyen46EQzNehs80oOwBqHuTTRN8zVLddjfcGzGBr0g1jJ0KIg
5ErIkdjxcetI6panZHIPyon1LdEnncpISlv8Ba8qSqE+ALZRqsIGfSr3FGgXY1cd
oKZdp2Jb2yVN+9PTW9ZcTxt99QkX78adMBJ+wp6S7x4Sc3i+XLBSOh/ddu3UVOLQ
IA+i1g0B0tUCU0yrOfxH8w2G/fdIpHpB6RSFPQS/Px6F750EX/bxYtxBvDEUND7l
EyDVh63vMcdRM6KZPaLs2VOVEot6FoJxyD7fqigXQM0Nrh7jUJMIDyrzbBwgOoZP
XK2QRxEZhILM9zzFQmTmo3MI485hSspyRVyTTUTTTkpzc17tnO6ZDDtp2vZgcK11
a6YNJDNKSjPkCTJ9mRHK1aeUz/W/gvuTde7lVCS3yhOdlQscfeyy2DQd58kd/BLm
FSGwaJT5YDioIBSCRnCuZK9DWBzB7RCYx982vKcwieLAbNxDoLRCuWFdET5b/B5M
BeznkifF4M6LZFT7tvZTnZF1+WLZ+bjXBl7uM861+CA5sXVJ8G97Nh7+l8310C4T
09ZVFs6Sary3E+aYQ5G7EaTORJ5KL8uqlOdMgRoEhjCvR33qsM3jKLvHEhSU69te
1nlxOboWj76bFp0NDvUofK3fKPgqFlrb3VgEOWMF53I8efaft5Y+wuE8WRDvc2oe
VY/xe8gg3WXHjgORGozBB9Q4vROKR5vPIMJ1hOITCEIk8kG6HD6COA5CeRM4b952
i6hN4E8UeK5XSaNISpw3sUrqhYC18YmPB4Q8M7iXCgHsmTCIOKB6d82UqGfC/27P
F+LWwTKrr2amem2lZhmDQTRrtlcM1JbEI4eaUgTIyGVp5QyEiTwUCRExu5Sm1flq
2mQpic8t0yzjwEYqzO14UvTUSMXhUXKgkJ2pkp4/BL0kCcIIvH+mdSRdyLy805/r
+vI7Zh8n2cyETqlMCep1EgBPnwuwpOgbW38OHTgsG3wOMq76Ck7hWXtO3jaUGCDf
8L+bvnv3wu/Pp2QVKQf2P3Eye7bBp91Bk+6d8qW5GxLZwUBF/KQ+nDviXvv19kae
zyobFMNR5PUhurifF3on9BEc0IEPFarSpTS0sme4dVzv4y3rh9SvUdystjCOO0C9
6wPZJ09bogAg1DXzbEfGBY3lpKgdBczJPAWF6e0Netk62CvH3tq3/mjNP6AyVSvA
BmS+PgH7CqJXf4vh9uMB0Oj3v/v+uj87Bd4WVJ/rjGZIcAmKKY7RLP7RyC/NYM/V
uASpht8WBppjMOoy1y/51zbvK+4apZolfUxzK5jgzUNHe63oUGX9G61fI8KHXRAU
UWeD6S64qLxGWkPPq252xURGlEoDGnXtJ6cCzr7vrKaJaCIX76oiT64qy0VH0e6b
4J3t8M8MCOhgUxre/mcaEBlMHHD3OvGeNeSd2uFideESTxwwoxZIg1fujmMXXNMU
Hq4AfewZneuiQbskpVULGrXRXQyiNqI8g175D9Eg2cCJv9wfvM4aQaZfiGPqkLLH
XSktLyIwesBS6uDW9hYDSSoWM2n2xdmMcu8Yqw5LlCWN1n3ZG7uigvHxhNoMNbbI
GBakQvVoV2v0e7k3WdODtHl/WbfLsv7KDtBqupeVtRAG7CsEhZrP9Ehp6IEZZKfM
wModUkufLlJDwKK6IidWaoH9FCHDTgu0N/c23Kmh07xGhq4cDpw5dA80bLk2SYNO
iJs4ib4wEsqX7vrr/v6jIwDJJY2BUhvUidcCxetSVqhz2pAU338ykD8FRIg53ws1
/6cxns2KBFcTLVyKg3iXGeEGIrmdJBfbh8ic0Z5BJv3CnkaOlEs/3KFPsFSml4f0
/UXnIkvqhyw9tSzStd8iCpg5WIKD3NQNHDGs4MB2CgGVXXTB7fuSqUzy7tQQUz2p
K4tiP6ii7aUNOb6MG3Qq3QkyV4BPzb9HTSZ3Fkg+Zm6HGTwf1BX0c77zgyX5J4Zr
rbBqV4wC5cMnUPluDOFysPyQBcbBuKbcDvBf0otcll8x4M47XYaEyH6L2QeYJyDG
WGY8wUkqrVE8EHUyrsFAMpb8EEPqTdmzH2SDe2eYVWvsMq9d8S4F2ZEU/Mg2D4yj
tXchg28fR0AueVazZiFm/u02Kt7R1EUpJTaq6f5ZZX/XbOsrxZjqsBi7JDady2cR
F/7CZTx3arb7t2/5LCsp7m54sox3V0n1FfdTSLRxWmROU3/U71Nw5nkNCU5Jt8jI
uki3Dc+5qk7bSiIk1Rav1F2Daaw7Z/iUSNfdp/hoyXxlW0l/zX7Db0PSuGjqW1ZK
zfZIqkGlbwqemy4cNIjrmUqNIFK9jZp1L1LQiJzLWjFHF7PyTX/9A/D0xUdAigd1
yIkFQyt9PtWuKGG9uTqH3O91r1HUK1xry0sDqRrfsY/lWYz8/gH/0kjjvecBKw5n
7y7MpWVmwzVTTQGYRICTrKPY5mpDtDQDPLPgB6Sg+7ixiPRBOCSLQTSbbuc38Xt0
6m8gmJgzA4uPBZLEAyZBA+GTruSfUGj5I9/U1XtYpzuaiPscKxlDqfX774THolQH
WX6r4h4IIwJaZ5lxpK4eNw6+6SRmWq1980EvqL6NXmh6fTPhe4UNH8UcKpae42Za
h92qJLImKypdy5gYEHUFXIbw4OT3HpuL9uTTPUNVdXUO72c5g94UZN4CF2uFuZiU
PGt4xNPDqwanP8qYeUIaUkizi/lzZlZe1c717EM64OIt8ivoCSZ1SYoX+Es9oaC4
i22VnyxpoPBHia6RdrGfxcWul7omO7Eiqg9ikYLJl9SkeNM2k+sXkkkMcAsfUgAh
SeUumAUGayAaJXn7qYAT3BbBhHH/y6SZyi6rcYJIgh5xayBssyY73h/JDamTxtdr
0GNkqcfYgxRBwptXcxBoBH7u4SUEE1OFwfCORlTgnVsPiIGR8T22N+J259eXpv/l
xo5pzFVJHUVKUZ2K/bZsdoCMPIOuJ6t9sNcoXub7utf9AXEHl+sQa67SWrY4NjUT
6much8HNLB2wmEd2zwtnBVrU6auaNZlpVznKtZmO05Yo7VQspz5SZqQd7Wyt8Nn5
K9JAHLSGPWN9Wy7lGKhMQIXLLy/34HfV8SSrL6VVCzB4479VABXtazv2zuPkAc+i
QF5mDgqlylFfX5KdrhEPrpLwvA9470s+Xye+xPXpE5FLGiPKM3VMpTGGXq7BCdXe
GtHQmhRQktpztgP8x9ht0O3zuBGLL5hZTQH6vQgJIR+SZjhEJ18cL3Y+jDsv2onG
FfCHAKCcKy+9khzk53WTV979bNIij3kNLiaw07QFtxJE1lgcz5SzInRgPWK6bwp4
w/Nu4f9HxpASOOaw9earLHObad/ochtsPQ4eUGUmilibppv6q4D6shPFTYQzDCRI
dLKWI7cVFR7GTNHaHj2xUdLb9x0JBRD5zXLIsWcXIUlkp22c7ocEphXgvHgssWjC
PNG595HSk1HCePgSHsl2zbix56WfJ3JWA5Whbb+AIMGXZgytnnACLFzfxDxE5TeH
UPejWVn/S2ZuPp1JatkZLhrpx2qgOore1B6TCvfu+jJMaLYe2paRQr0sjBGqVv1p
ToQ0MkCPK7TeBg+Q9hu6UdYZl3ZzcbpR6VrElp98s/a8YcIJzjd6kf3Lg0Q8Ap/d
xwRcifDlYK62lH8T2QlKJ4VlknVAj2aLD2m2wg4RcL0Dkwrm8o2c/l43loEELzFA
kNKJLfWKv1qBtbvSweAiZRl6g1djqizuuODq0rmFtIZ8Cg6ZAjuGYgy+/c0VVbz0
KjjWQwL4AtjZFH1QW/b6pcg3PEmW86ecesk6bvR+Gvkr4jNso8JObBfucZ8MeNRG
1Y/y8VRW+h3GYTRQww5oV1Z5ef32Gs2bXxxTIIg2bo7+Qk/7VYEfI9dQShllT+kd
alw1pGeHZfJiy2ml1aa6/ZiibQE2CzjS1lK//Yr2aLLtXU5EYJXA6ANrIPpF0+vy
yBlf2poABDhC0vp43Cw2efmXYxkv3qV/KQncP+uQO6EkEtTD6fUjUO/+To2unhWO
3/7vKNTSxnRMqf/i8zzFTGANfL6JwJPuxoGxUB8ljiYBuav8KwUApPRfH4GWE4XJ
Z/DKDy6Tojpho4vnF0hnLCwalH4opNi4/+uvONmRGExVVcTg1F3pL5XVUuyCyEM1
WJoSHaJAelezTYl8w9wPdj5kr3QZVgWpmTxQUGRj7haUM7x57TVhz+euHta25QoH
zu4lwQxvKBSnCS2M2ex3VFAS80N1gdVMudsGiInNQtStz2+bpYEU9+6Qs9DNai3u
Dgr89XNuNWx3yx7livYFIu7/2fxPLYGEOPetH/f95QpPe03cQJdOOfJIahWIQT9S
ufmuJJSlcnSdMtmiSvchWsfv0YoDEBDil8YhQyMCbPpbG6wC1yskIMzx6efOmG18
UximwFXptyqk3S4TSeMXyGd4cA8g4sFF7l0T9ktWVLJl9yLFvjwiwJZJh7unh7Qp
0dOxzR8f75aWfC6MClHPJiqHk7m7TTOVKqqbYxMfMIwuwhA/K4/hxVtr+p6lLzLe
xcO9OFBNt/9NfCMoMk8Vx6bClRekhhvhNjYlQfolT5unWimT+ihxZXOaJngJHmXN
ecm+ha6qqv8wu5g290AlxbYuqo3Eqqn1R2vCDlD8/W6Ks9EA2iclLzX2W4clPM/D
LymlH2PDqarA48uJxmvE/L8Ahi7PY+Zhm8VdcLtzogcQ1v7Ibr08/oxkkjpxxdHU
wyY0CmluI3g9bj/Ef+Z7rlOFtjh5jgWiUx0Wfl+9k/gdfXo4/1ChHSmGI0YJOpXr
6vBH6z6XJX6g8Yp5e7TUmZPmwCd2zUOXeGzXmpz0UortziOFwNi2IJEyIFK+Jznf
5j5EObF5oZLPYy5jbNojXs020vrGg+Y9ubBbyGH4f3b8G72Ub5TwvjqFC36JsuS1
2qypib7FhrqOoXNCyAMAmjV5AxFzOloWvORMcAS9iWFYnBMzZyPqT7aNIiCafv73
cCkTbNTgBFA2/I5Y2V/jg0GWNNAK1HUxHjgpRqjYnadDzMsrjDXFhD0MnOFjvHBw
ZJK9vOzik1KSAfa3CvClNHK8y4jqFxIw8FGaQ6X2Qf5ipEWziXu6ujgn6XJrF0tk
BajxzuW55na/WmezF/jDGKaAHlogO2A5HxikalbuniJQoThfpMn1rIPudvmHbsab
fpzZpFe5nO27YKrwWb8WUrqzy2KtpZPO+hXjFW/RT6SeIRVVEs+hYA48KjYUI2G7
cAiphSnciw4jJ0Xaaa+xU0o3PCysIeeLf+LqZkvPnYdFgqdHGX4BjFyZjqWKxHTc
dsX+6ISOc+7e/vuc7qezssvxNHEGr/pxzWGEC4ytkH9Gzmr1QmJgeZOqkEBxCi5X
mEwTOibOc6DFalQd/f6LNbGmKrRS6QbzWmOExk8eIxVBseVioy/88jXBIwRZuxWD
odIXh7W7eqLATxCaIfRrya5u7wuOMvjR8mNbQPGAwwzvxyFjzuRKiToy5HLXLSop
Mpwu+s//lLOT3I49OtOa7gkBPkx2OFWqCXxuc3Cik35VVg9JPbYJtRNJLGivOC1R
BCmF4olzYby7AwY1Afb7dO5FXwMA2Xi/c1GosKnbBr0j40aw+mYM+Ni3QYtQpVLh
P/6eaGxhAmtzLCqNFvgGUxPtbqE2uuHPiXV0+75wxr0b+DN07Mt0NzwdrVS9HlRb
nsTnkcdTFaW87r5fYlCAZckPDwWtIW1hqFm2z97OMCWSDfiYDAEEpGm4GB+Bk/uX
F7WFHAvq3ykjHNF5jTSxaXy4BOe/hGLYBubgoQb29tKoCNgPi9DvUpg4WxtJE/RI
4kpq1UEebSLqdVzhECqPezLH8EM8G0faDifJYW6Nv7toAzi15UxURM3sKZGKwE07
xn/hiZhwwhenpH+T0iGvHn4aF+sx9vve5Ccr74rYtHWTfpBqG7dVo3ADox0hWB5B
U0elvvkCWPkOwXubeKbVaeCFv9o7KftphwnJDylXJUwIUmFm5M/63ghKNwxRc0k7
yVb33X8aDtCv6lhvjkQu44S5XwwRovHPzvrGaMyufVRcivKgsJXgPd75Nd4ovDy+
0WPiwqQqKpScvQ+Nb5pRW4R2/3uGXKJcm+bj4kiNTfLiDo+k56eKsqX81jSh123V
f9zBe9tMyU6GcOrGhO1AyhmlzVOTWh2Jz7JBj2GlVOx0UfUh2dMSDLds7K//rG+O
dqt2Y5SPnVOdAstbLIbFyzOp4iLsZQpAY42I6myGRQ7o8f8XSyrjSSyAZbDyOGc0
EMKNEUbwCEuYdzFaEVdUnKCQq/UGuS/to9D9N2jg7WdxbuvIO6Pcj5efVkVdli1O
+ZAWTT7VN6Sz6l+/xVi0+GsCM8J2gN54TGNqAGCskmVxZ3RikkkZyqU2pEuqGOr4
FZjFdNQJ2gWBtZ+ybEtDIog7hGW/UigcEeOL+kh+jmofUAX92QLBBYL/YQEICcFc
wlkv8sdY0NB0oCeJYl0lVvI6flEr2EJ2pfUTA02cqBFTiELIZVE4T4tSks1OgjVU
kFslyR4YL1EIB200SnbovX+5qgVQcs8dgrND5SXi94mPrSIUlXqbOT5vQzhQ9i7S
+LAE4qyZHokqJAV6Wskbb/+BAw3NJW0Z6HtKEGi+2geg5b4B+5IX2yFK6Fm0hKVl
CG9b/iFYpFoOmqIAMjYJIhhU8Y9y0baKE4F9ciyHqMQzkPYCt3GvA1Wmr51R5LL4
giaMWWEw67JzKDPC3qVzbHOH5j0rkuOV2Vd6vjkMQ9tFUyZ7tO2Oa7+GAtqts+tC
KyTUUbE4deBa+TJCbI2DwEKdoAluRvRw586FM5FZmxXERT1MPZC8kIb5/6IYbDyp
UmAkYtl55pK24lD6nwREMraTID0sLnFKVitLc6i8mz7Z6mAKgrow/1ccwpGQqb/l
pZY8U+vRdcy/srMd7i+2F24+Ov4qOR7jqlYiXgxc2gbEHEaR5iedCCoJVX79FZfg
iJLotDl7TkZl60KYs7Jf0iSSKjsMrfZmTNaNSB4p7Qa4kEm99dmWhgoqStf71oeF
gy+WssL7rBC8Hzb8XJ+8mSAhNOsdjmvMEtdYHuGdm3wkmMx37PcMNUjPEmwITsI2
cox2B2/mtXm7KnAPrdlAiHf9Jukk9dVabbu9jp/Yzyc2HlPAkUPgw9boOUTE84RF
Z1hLexcJQC1DcyvTPoC61zVoirAvzAVOCwL9jykmGOWX4f7Obba+iG5dFYjDC8um
MI6IV/v8phjGA/kWJN/isrMJ90fn4jnXlHeLQXfKq+yk0a4Brjbr7oeG+GuBR79K
3atGUoguwW9g6RMAC5H28T+JckgltBj2oYmH34z8YhVXClian6sG+r8bfdTfKopY
r9infAsM0X9jMooMbS/P595vzyYP9HzXKEyg3T4OM6P6/jTZpzMSTEv7tQG9q+ot
SjiAM5Evq6s8jLxS789CMv9cnWZVHAAkpy96OXTCdl7mMvyDolhijBM1+1ZXvMK8
LHaxHborsdhzRxxKDA5PmeIb9IKKqsoy9Bbflzf3SNkxhsRl+8paQgGrrOCZyfTj
2jeEH7nbewwcdaSTTExjTvE9Q/Fx2afOoTzjFgbPZWP7qN9vhgvJca3sO/ZZKuft
R+VOoSMQk+0JTAQLgnR58P07OqfZBSD0K6UilbYvccrrh5PrMSy93bH5+AJLRkhm
8c8oUUZWPYtK8yRCU0AlN7/j0XOCMdoeVCtj6Y+ZUnYxE17ab7ovkd4I2QKWB1zh
8z7NcNBi/bZty6Ygt0jwHe530SuVJNHnZCRoS4F3smIc6dc3hY3ar8s+Wd/8DiCE
5DRSP6MB24NNXK2PN6iREsjwSiCLHfhbXD1nk/ERMFMXJEb5GUvIs0F3AQvA/4Uj
ldfcpxmwD+mBBHUnAWEoVbVs7KxJBb0HBgcRnLhD5e9dgVdW/UieC/5BCS7C/89Q
qt3b0SmCey4ehrn66T4z0Zb+axJgCj6C0sco++r6VwYIyqp24d5qpA+dR0nLsF67
aXFx4bUC8bTzKgPhPLb23iq+eiVEjOqAmH3wTGAOg0Bub2kUsAiHcpvntZm4RqKa
8NOA3GFFAASy0JCJWgmutnEFlJy0F6rd6wsIKQhGnqHSCq+KFJXbnzzClnJX6rzX
LnkJFaGM3EBXlspb9aWbWpIOW6aqYj3A+F5HmIeCOhGTD83OpYKDbmaKn9StmzlM
dIOib1jx3/hBj76V+2/ca/qHl7wemUvc2ycc2C4GSwQ8kEHTgI6hZ5sneM/M3Ynh
A7iUayw/gYzy2nBwCUmd/e9JRniIPSwYCFUmbK/J8z8MQhyxH6en82X0OuCHH36h
LZqg+b49PPMz5x/qzUvEVoVAcddVDb/r3qhB3Ht7d6EuRlAnozyd9aW8UWS4MtWv
LivBpSVlleV4TVgmn13zJX6l4ZpdpZE3t/4PwtkETJHUVo9L9RjqvEr5v+dgKv/A
NGgRL7WKLgw1k4GBcwlzT5gygmLEcESEN5UJVnvmagQ8T0RrbrV8ZbFOYxqStmVG
MiGrvhNW6OjF34B7/OVjt+RQKeZdH5vppenWjHgnFLJfnzxLt8L/Mo+dVGDV4b5i
/zsfWY3bqmHPiVA+mQVSukEcadHxUAp72MNACrZ10g8i2dGn/zKZj+X/eluSp9Sn
/yqMdRNW88L0vukxbzA7UBXOCrduXy3gVdSZbXge23hlMbkMpcos+sYk99JGYWOQ
1BZKSM8q8AZ55j7pCsGZ0OaqclyAi6SvlwcEEzIIwtYyFukx6dSSFJz74EiNwXpt
TqWK2vNHbk0XVBq2SbJLiJnf7ssd8i2OkfYYxP3RcDENHbLOgFBe4Vxp+8OgZlF7
LVuRanMIbVi8DLlOvC0et5PZywRcj3yZXaUP5IfDbfvdYBKcp1lJ5sLG5SVBqdWT
7236QyWkneGean1jZ4UUpeuobCCDTdzoCwnof2vCQq6etqmCK5P5FmGu+yit1Q2y
8jXsYGSmZRfG0UB+rLuYTjJARWum+puy4qgSt8hG0zEm3fuftj6fFwj6a9EjYybz
4J1xoWprTjvQgmhgaydGVO4sAIu/UimRWtz7xVQXlIlv/arX6gcQJaIvI/uunbOs
CBa/95SNskY7aWFMnA2z4ePTvQ0zqEViToPL8aIXkUF1TF7Uf/t7D5Fb2sL9EoDR
wua7RWL1obuamHLzRD8kyHgtEZZRkG0DYOHB+djuDDrQcrJ+cJ4WE3MbKyAcQGyl
LyOI1MP6apSg1dS+w/p96nP2//JoKJjLPrd0Og5ukPGyF9qe8FEUwch4YINRYkHT
yP4fG4KvdukYnnEAo5ML356RCkyIykkJnwXuyW58v7Gu+jHVfvS+g6kbZ3/8NveJ
M8KU5PF2Sa6cWcanrIgNfkb/XL7M2vJ1WWIOTVMUPCQoAJg9Qta23bObwvjlTs/D
0hys0tRJ6IWme5dsZMJ3kgZXob30bmFNbo11GQWyBBTho6RzaOUjzRWOd4ZZbRZk
f5SYmPMKG3RAhYVFo752+wBUsLUapH52AAKtFZ/oRri5bILF4IhxvOBN5oL56DAB
RA/YXxMsiLn88fF+50d1N6ww6zo3MZQsV+m++XBOGb0FggPie4fHNOjZzRryAqmJ
a8VZHMYcS+Z5uUFBxDXiQS0hq1tn2oP+Gqu+eTarOC8ca1ipR0DiWuZ9TMe+WSMt
XtwL448IcVXmvJZDaKaM4n8SbT7LqEc0rRfdlj0L2XzDjjyh9KJG1n9+5WJSsAxt
Y2xCyr87dlzWPN+weu10MGnt0sXn2eRWIPK9KXCOxY6FGin7ouyK9wZwLQ0zykYH
G8IjIf+vKUW76UK4W3DF+2yi71k5IWmtH9fZP3Z8QfkldBNsnh157P6YKB23UmMx
k/N4DJomGy7kqhGu1OTzNUt455SZQJDnzBz7tUiElmo1Z3CXGIDMsfF3KuOlb7Xr
1gfrI32xNTPhjY1p+10qNDAMiUZkY0OvlKn7cwlqYFvEVy/7NHezRGqqKfatKrFx
wNcv9YwvroRwYAfn5xzuyUMU0BPBgd4sdLe4fTKND/RNmVzhqS7hxwpSOEnusMR6
6YoVcRSz+qdpVFTRHmS8v2aYHy9pGB9mYYlM4ln4Bgh1nmtIVw72Uh2FrUbjqEht
FMoRPBJ1eoK7huImgSzbWYp78rqBtSKji6jYruEG9gZFyRh77DHubHoC8GsmLdHb
qQdsDWN+1yhx1KFX3g9zLttr4xUZTcNxBjn92LqUgR/3IsI5OsEuyswYFKTUGepO
wSkY99OAHwL/4FdK/HSi29isqFPs/m26IZt+ZJ8gCopOfETfsEG8tyQacyYuDYNe
gtplcNMXbf2RHlvcIe6g6X3sviQjmhSJq1KGlvPyMLzPVVSzTngaPGZ7Uu/1dkCk
ZrTYV+gi8JFMINDc0l3+i6oLf84C816TxGsMU3ds/BhdGYoUd0Gbi0ZqBt8AYei4
NkycLvxQlnhxD9z5+V3ovjuDT3WJcC3Sjg4KUVVCqKz2KEFJ7O/dyMKReRksH52B
DZr799Fm5ZMJ2cIjfDsJVmoTLviWTn6bjvulQAsfnZmHPTfMYwb7aCM2uo2EmpCd
ModaXu4v3D/kWQ5CQASn/RKJuyTMFmfWbvCOArpXeugOSnwRUwGgf0Rlb9kA/w2I
t9IVgilxJWIyP57/P1SKMJWim6f6sf3re3Tezcc66Lorx0P/EXP1xPnWlzi7T2xd
8WzQ51uyge/yjYpLUuoyLxroTvJ7IkElpI2egMLubq8naHoUhnY6FJZ+1it7OmL+
m5zIaSsbAgE1ktlhWrAybAgYehBrLBLl1x0Y9wwpVOcoRqrVfnOrNlzIfOBwfeE7
D6xFpHBN5ZTyVHd+NEeYq3wATKkeJq4AMnj/OWAA/HZ3AyRiCWHSGuIhtaZFJHbB
SMAO3uvzF91JSLpv03ARjm39nw8b7m4BRlZjbGKNqN2yFw+sEAiCCcXlTIbayogC
ggVDHRFF/U/C0SdVyB2Y2p89dkygIrSqOuX7aPO878tPrelQMUa2DPyvjG52IB+P
itBryyWU6u/hpPaEs4cPwMr+MWYHDzPE52K8pnuKVV1ktaFGENE4PMHiNiDBwOel
GtvOdQRdRIQjNpEJdXjaVJAdxqwZJq+VSTQ1cNRO8MaY51Gt5ctRRRSQEwrC6dVl
r2wsahuP23xNDiwI5IdnR/a8sEXUb7CmtiH6+h1bfCrsA7+TKWjkGvnqgfNWVrAe
7LvbIu29cB6Y3b8KqjnDdH0iuSIMPcXtaezOyVNKjeE5Hi4lYoisrCXedjn/HC9I
Io+Q3OZ1Z0JKd3Hx7kjTI7FHXzjenziwZ7xaotplCiMZuPg1aHRci6Pc7Eq/ZTpj
SFSUbT/EPPXxvcuyoblpG2yBUhCSA4Pcsqtwkbey9PM84xJkRn9b7bTucvpxVsnM
VCFjLYeT5cruIt+ybvXZPNigZzrww0yZrcmmyDG9egGAQaVqDftWFV0gfH4kBdgr
jOTDV7Ja3TTNkai5h9cm//yNtXbesrYfFFBvM282+rCIxM16wQr/XeNP2HmUoHFg
MQwzzeeEYiVuuqZWsd5fe3jiMderWdFSh3uiNT5oU/zsUYTs0xJBhHJkc2KWA0kn
GXKiLNUeXbi2AlaFwh29K2tGMTx7PycXaN02oYb42La5MCCP50vIaKKOvXJxmDqi
3MN/Fkvw8Bgz+j95DWe+yivZm90If95l9b78XE0BrM19OimTw+JS8frxxodd5qo8
zlb5FXdl/rFx+5Kb8fJHRgKGcduCeO6ZaL8S6PFBtG8IEwEJ1RpispXitJErcTvm
9s9sdhohAzKgoTsBkB+xzSSaJk4ONhgRVValkf2aXIV85cuCVbnikSlzomSipNlv
v/b3P/Qu9hGKmn75YoXwRiXGt+wCvNpEpoq3yeEFBXbuyzKK7402+dpJO7tRc5eh
rTy+nN3heLHTt3mZ31zbLjy6B6zxqv9oERCsdQMR73VvqW8JvfQhGFQejTtPbGUN
yebElZxcFEHyJjm+QVeT/POGe1tlkPWAVoFpQrI5lFSOcbKvpcOirFs7NiUl+1wv
2rRAPIXigv8Ehv6qn+ceOwqX0RHa31gn0yxz9SflX0cPWNsWief/5woL4ql7NGQ6
tUopje34ByCrzeUq0kNbeuf19upukl2oo4kpE3pF/3NpkwHvLrtzJyeNt7IDo5or
/Akol4+34OtKU/WEuutDENQDZxNR5SUzpZPOFBKftKLd8MotarxDn4Us4xaaU19E
4Ut0ao1r+BjuQpNLZ2lqrk3y3dCo9QTVITrq+xwRUCdFp45W3q4QAabA3yWvvGn5
70Z1ZVGx7bjMZsPVylPoT+q8trmvEyPLAWqhdI5QOZtYava+8Pqghrh03OnkF480
VvSfPEh5kMGH+pEio8IXezSHuuOvhFU/bBYCJIdhK5OeWKDFjf1jbVNRZvnIizER
0+FdfyAE/G0kso7IhQtPnbVhYqU7cipDAifmcwwXS7sWuBTZbpAYTjHeXtmorFdy
EJoOXQuiQpbi8JVB6UM0FVSFmoUzCedtU9ddHL0u6KcgZU3j6lpSv0hB06fbndfy
udxBuS6+S/9JXgmm+hPOUx9sbyNMLnx7ADAsLrgAnfEBrVJRNdSs5V50a55Mvryf
LTCrub6mLukmSsmMJXRQ7OL23NH+z79RVVw++63bl0FBQc5L9UawjSbaJNmxa/vc
EYtIxyyaqWUxscyezQwZYclHvSlxvdWo8BZsdU+AHn/MFiaPlbiLxkjBI3x3Ub/g
ctvcORqDhgM1cTtfI8uXrAB+T6VU6MFYhmWdaQ9MjcGOBe/5a4Kw0Ho3FXh9wkMj
3e16DMrHjnciZ7OqS1W8OMeKXAdl2qt0S1ZxkhsRmyapQxKmXKA6xVHm/t9YaJED
CiQ4We6BBLg2EVdwcNYzG3LsfJANag0gQ5MYbWFxrEBztXE8epYDM5KmnpKnRjlc
g3vMK5uhtDnRDOhdFy0km385Zng7yeBAm1EMqPexmaNgdb+yktkJ/THlzEy9UTol
yGJ1+5Eh9C2l/OBy1YHja3goPxFrAPE2Tx1Zxp8FnRLV+2RPkfnEfT3rLGX6Sl+5
zv6/sWmtXk32vbmwQ2z+9Cj2TIgBA3NLiYJsPJJmqjRRH54lbmETeNe48KGjEBfN
EVeXt+zHWz4/8YbGA1mXBXdnTgrm8mlFvpCd5ZWXxqjTPPvzHE8/ci9x+h8z4z2+
9hokIvP9jdEGQ8Z+ExohEgdbubIp+Ter2e82Bi+NMtCRYoRjy30KpBb75sRTaoAd
rAQsAQ72rEtHi5DEsS7cI4mkLAfTLh4xpZNbiekeaHTKn4+2DlyPwrPgI3DgGsD5
XL9OoPXpJN4rN+GpE4sauINLbcypFgSkBirYyPBvSPyUXbInjFvoFhP09UW6cLPX
stX2Q/E9Ow8150/E5tnwqLHoNZVopltCIIUs8amAUHcZAMo3I0+ixUNPJhUw0lBw
cZAGTs8NgnARFe5Hz2xSXyWODT7hENCkljxsH7VOe5TiswAd2Mdi7bMYc/18Ae32
To+wi9ANdj/F6dc9rDisByKKAwtjRkncMZuckKpGAyn8w48jSyUggjwmOjwu94l/
uGvFrZbd7Jlwcx2gS+qjN9La4WrflY1rKaoXwyK4N710m6mI0X7hTugAbxgDmBkF
XhOJkHz11JN6pQKgEokS5C9oh5ysOLQvzYt5qDowlMqVfcK3pegMUURsrMto7ufp
HBwd/EJRj+ld45YCqZM3p+jhzxvOS2XIhkXzEcz+WFatdsA36vBdgPYbFZixKED3
PhnNyztK3Q4LCXVxPlTOUSEf6WTZ5FNSAnU4p5kWQm0TInEUMLaDFEpqfYNFmhdz
vc7FirKvSLzS8lRIHpGe9gAAuPa5jgj/IMVFi0Ol3tKfzRBavrs42ZSgjSG5NNjH
Czl5mvwFSmunUwpUNkoZvV62LxlQO2UY1taze4p84jIxWSQdzVhIFSEg0a4JpLWA
riiY80SZfxYUP+WgsoTKq5mv/iQkBVV1+n7ZjeDpnSk4FU5klGQMzGKUYgk5YsYA
2fvqGmVLFpQ1QASOjSoQEx1Gb91Kcs4YX498yXpH+j+r3Lo3am8Zn2/6QIusjWG5
6sCY8Ik1LBCXcOJ2J3o+vpIbfo0Vz9JwlZBNvQN1sPfJyZkku4Vv5YHEEBfyxZdC
ncTSF3Y7fl7MXGuPdDMLRfrwR5TU8ix86UyThHjbGDxM09Y0rdRhL7/oMFj0PJBO
jXDegJUxyGVXm+OKYl1JDu1dUblxxrl5ooCkz6ql+atBfm7nBRthp7heI0RB3iMQ
nHYJICzliafqChI/iXE053/l2Uivi3kG2gI9AyDN2TXaOBNNTse7PiooXRRNSYlR
lFlX8mAntkrBj/demBOigTEk+E44mfYUm4h00NSMPIF5W/QVdI3i97iSXCrACNav
sg67eu9mxO7tDtok/du8B9JETEf1Oib+QZy+rIsiEX/mGolM+CxtpSdb4Q+sJEFI
pOoMMz0H7OhoSbm07fmPCZqpEbSgtrjXAY/z324d6gFI72ypOnOoNzJdkjXYnzdl
M1tvlnywIMteuboI2eNeOkOSJdHsWUvSpVqNzJ8/8NOT3GIMhlr/WaM9eu2irZgm
MgBj2MHBv9ZmMdQ1kGCOrqNIx97kMdkuC7Je+W574+D4GxOEOB9hK3uENimGymh1
hbnIS+NYx0k+gDJhJDL4xSNMqb6hH0amIoB619+8ki8YLCs8A6OaZdqB9zLXdB3H
5qnfUPBmmD6j5mhuwAiI8dTCeOsu+3NjjygTVHqUSJyprCRy1S13EJjCVvy9ElAt
jLJohI/u9hMQ1cwMnigA8UP12oNEGxlLXqf6753VlOC3Gf+M2fXOVqs2D5hljFEc
0ZlTu0AGdZNux1uw4+amHnR7CGdphrJKbwhwbdpPAiOvl4b7RDaegaBYg6JNXI/D
qEgvFN/SKrM46f7mZT0HCseIsalQa5qGy6eeKlCvcW7xkjL1wg6YEMh7JliuI2D0
jXcXs+m6x0kKeuURmpEbFRJsFQi5sNkqh7qxvBqv6C6Yk4IITYr4iWf0thr9Lxl8
8d/mY6WJy9vk4Tre4Ezoc/uws1izQ3TpPhs/YV5juHpfYxXUdGnc3kH4kNCEa5gs
yWd+3mjFwSJVVZKi0eNDHMB18ApqEYNtruxIyI/igGSW22PKEO8c0w5KbV3kFrAI
SvYhKR8kNRzhfLww3y3YRoZT1PjJsQ672sshLejgfe1xc8M4MLP/WSRdH8E3s0Tk
a1OYFh2dIdllq0nBgqOkcboDK0Y7akGsLbcTO9vHAI/jvn/2VTwjGjREHv01b3Hi
FJtlTlNOvNel0Lag9XW8HRz8N1fRycArvkbW71gcR1rCfBpSJnQAPAMnv7OsR6hx
H99vHPohhMFmuY6TCZbGu9qiLi/Jq9OoWxN79umNe0HWxMfB1My9BcGJzWRbl+Dk
5hk0pXJF+qkrYKE+4l5em3Zja+cUZ64HVbWqmLYBU2VtiRZe8ZC21nhV6+txTk/m
a3xCNvnelYLHv9NWQofOyv8coQBUPxCGzX1vSwyR82hBdns3wwvjN7pzqzPmvLsR
4VHuP57Q6HouSg4ZYXM/1oCxUavcXjIcv4BLl36/TwWjj3MmLKt17UthBmucoR7Q
A1rXvoVHZVnNPKLflSulHTl+sVduUSw6ayO19FAxPnOdsO6UDHRfYWXi0Kvd2uW1
F/yo5nAW+eEjI8ChC/c77NZkARY74fL3kPReWagLlCEyWOfIwYOu1AdQmaDCcUNc
mJbhtVGu5EA/9YkrZtbIUHE0VB1bVa4n+XIuPdQUxreEKMverlI4YccUw3C+LBz5
wZ+9mHw5JAWNzdlG7jvAZV2lIZQChUwZcn0rnjQ+X50JjlYYpMRRFg1+xYMCkD5U
Z1iys0ZWlmJxoFsUzzkCSxvlQmq1BasvqwsE1MqSpeUtEwp/TmTsBUnakvRc68L2
RY0MYx0eTUa9OtEiTApucboD7z9EWsBDYPj/GG7JEqIvKOrehpshacdiOgNOh0Tn
6Sxmo9rg5o3a19pPmuK26C3M0q50J+OJoNLKlK/m9TYqdNrJZGZwIwJnPoIAYTQi
VEwey5wBpLjWZITwAUZ+HEgpQ7YatXQ4vx+9EMlnEknbVhj1HpZVKc482713EQj4
0p6X82tk5Q0VyyXJsB3GylyoC//I/t+6cZ1ngicVvi3X9WeHx8X9XtTkW8aAZRve
ubLL2YOi/uLjQs+7lwADdAZEqVBquUo/deajb5mb82QycLqJn4RX69vHr7SD6Dvd
oKJl55EtrlWWIv0St2yJwwdjIXD1d6ghwrsrsdmsJYDhhErEPOVgiSyeDjITtSIL
+U0CQZ6nVIPI1XS3+uMTFoTthuT6mSSHoito+bKX2ChFvIjbSscrlsXTOpIQOMwJ
G/h//7HWPK0W2XfdZ5RttKOdVo3XMGHACcFsv539Nx9kVjrOwdLTjJZnbTxr0Nc7
6Ynw5jlHjyLIw9lvxfldvL4gqjWqXugbIkPTmwQNpdXFO2/wYMQOjFXiHBVBI7j+
teQUD35bf3bb4yOM4dFGDk1+mgBLmv76bTPlufVTJaf2Pym8xaOss0RUrr0TAJll
8IPEnZDXaXH6GctEywbFzcRDsKIk2sxBVwOQF90Qt9ui4oeulfPgt1AdYmiyrK+P
+yp0gEHj+yGslh6jlxHfamCqFSrg3rGSwswzERr36j6zszpdHoHrKMn6WB2VV4Rw
uZ8kNaUhsnhXqCJM+/VTSMXgAzGUWZGYbKJBZg25dZFryO6ZbAoXldmsFhp0nBX8
CbirZkCe13jlxVsBxD1+pwYTerjewXY6LV2HVqcW2LhB8ErR9eqDQwfgCCJdAtvN
1zz2oOMMgZHAOBeSsuduVHmkbfML5zzlLdJY4pI3vL7+TM+LeJu9WS9+PLZbXGgK
AER6NHvOITqHpNbiL36brzxPlNrbQW0Z0ruzzi427+N4CwIMPqo29EN2sFYz2TpZ
nh516jVGaItbdoJOyWr0Ofrhe4b/iyC1jWowC7DYl7oRGc/tH+LJhSWdOh0XGbK/
nvkQgBunf8YwkjSTI2YhTHLwa+1Ya4L5dBk3ox0s3n7T20wAjxG+HJ5P6EUNvC2D
iOApWTHFT+pSBfqhXdUP2J0sHVMiyp7B7LiO9JXxktkBrE3UQWLdX6nhgkAI25te
sHrqdtA0qkpFAnMeOwLr3C3uTZlmaLV5jpEY56IVRj4f9JtWeEbTX079QZwr5665
5RTHxD24TUxRXXUpyjsSfS58P6wibz+D5wO9uG+4BPd3AjsuyGKMA0DBZ9ZyoJ0E
scpuxKoUeoMyqgY7pTeNOEhVUu+Rcth9a9+lGVT+3w2mp6qgHcpgSec0NhoRMN7z
X2SZ72ONiCjv9UEBQJ48wKWpYEjiL83xzGnb5cS7jadSxOa+6QKME7HIdCige0tx
NEP5R+dwlRr6nDEh+RXwHjXothnHIVU91N1PHTZH1OMvZKg+YxBpLKYL2aScqRzZ
rh6cwH+5s1wMp3oo6m4wK9ZTgRCRrI01TeBqf5RI9Md0cHaeU5JM/p6p1qadfMdz
AZnrRuB689635wiOG/hmElQt5rpUZ8Vt8/r0Csc1kmdVZxEFYL6zyAz31+VQiEkx
tK0WdrRUjMzyNnlu0R0HVYd4RKX3xAHJSZ1sEx+6hb+qFzFMm1ni8zYNCyngvTj/
haqyyxz3Jq+7ESvrwneGDncLdzvEaexzrz2cEeQnBqUcTrAUrTthmKRnYV54jQ9m
yZ0hT490GNyor9fUptoV93cdRpj317NsaIJe+tcTHS8pJYQZriIzToOmiRDjBUYc
7S3L5e/DboSCGKxuyU0J9cHDRmq9HxNwDAXe+w4ZxWqhwN+vYvPHmYpwDrXU0eEg
8gehZezyV4BqrxJ7bf97BRtxy1FQSpw7+XHcbshPP88G3LMll1dgNzqTI2XqZR6F
wXab6sM5MHgRLW2HsDyA3TpzrVeOi5l8K5zF8IOJfUKks8Kw3W0Tefq12rqkpPZm
zciup/ogPG7p8xR3NbRWpb+nMuB6GMCX/zHbTbrXJQf12Sv8eM9cakJnVN8isSy3
a6kyPXkYuStik0U1RQCeCtHUqVaSE6Sr5lPB7WTnwCqjrKpw57PQu/tAaxA4wec9
CeD3baH19Ren2dB+LDZ3o1kjpqqkokNuYbZhFXj2ha1NdHm9Rpb/9ZH5d5dbQ8Gi
wgubb+sp0oAEAM6pzkuMjXa+4TiifjTzRmMAfosHVRjlQY+7A8DyHDisi8cpXg2V
yrdUsondE1kRBsr8YPtuzstq73my1GDIglauD6XtT4AGKDuxbBlzuCN/SRV4sG8M
fXvMn+wNJrBF2asXJhiXFijHczdbkiSt3H0+6aCGwgkP86WTTIxiYcuMg+BLFLqf
v0j8IhNhjR4/DnbKLlSnJP2w3K/tcPKQ4g0M8GqglTJ/aH+O8H0z5IV2IjHBwYlI
i9L60FZXwM22HoKFnJXM6pJPE5KzwhYKzWYcq0nzQIX9NS5ENQlEGRokIbJqKPYp
fPZY+wxI3ppJG3+aaa1pDRpa4jYy/VVLa4rJV6WHjSe1QbY1s4VxDfu22tTdhNmS
F0A1SnRUbPqXnqK4zZYoRT/8wpNjN2Ct4/4JK+JYFOD3ajQ7C05oip6OTlYU45Ih
nZZbW3/YTbDzshATlVPSwWgDSehez5iil97F9+DzqrBqzXA0rDiUfwU3v3DCVOIl
Tf/qTnuvUtPnq3daeHo4ii0ZTN+yM/57bd/7WeyOTTe6d5MmdWnCAdRbNHEtDoqV
3lwe9/wwj5oftGkHFSP8lfDwjzB4/1a7ia1TWbpjbM6bR0VsAaZhFB4MBJvrgzyG
q8sVdaq4ox+Vy41eO0J8EMoY1LBce76MWscnbuQY1nlTfsxB10Pb08ULAwSyeS0l
uL6RtWuhYVqtraXXxemDai/zp83gN+PmYIz4JLSEOQD3WxGzd/Z/cteVyyK9FQrc
eXfMmBvrX0RveZEb814xHgKpLwTN5nzSn7Nh+IP+TlrxYLkW6hs+K7j+hzEK2mvr
wNT2oIo5IgLoU6pvC6qsrQN9LlXc7J7K4Sq/YMOW4xAdUitp/jrS1wd/cmxGCDBk
t+VXzD1PXzX9ge7BA1Z7WjlskNeNHhJUmug+IBwbGvwQE+P5VXbH+0NeYNMzAgSg
SgX+IgVfIsK6QeTkWeFcqPaKhu/keQUbzqqEumc3qapfhYXipEQtBBL6mAIY9kzm
W+zHjBAJ2vhp9Gge/QHFa65pG41ZzXl6apcbh/yf4X12ulla7KVV3SnNhoSPRYVy
phdfjLcCBiLG/4LKLjWBKETV3ro5EqiG+epQYCRm1108UXsSDpDLDpzNhOaemfMG
Zle7Sx7hMtY3NgfMZEg55vshgS64tT9gxT+YBjJPICkcqxJCG6cM/YICkQKj5x6E
KdRycl1hrjT19XWKMurscXmcN8QHNfpEmKbx//19H5hM8AFJDxzyCb1YfpHg8m76
VkwVbmN1vktbeD/HofOD83fe6aBCK8e+k0hlUumxppGN+I1SqPJfxW+3OOxwoQoV
YyR051Lp2kH86ZM652MeBl6t8Fijla5Ir1+ifLY3Dcqiy7rkyNackfPTRBgHeAGr
A07dd+P3BngmrT1e0agicixiUSZZtj/b7/+uXPK0CubkmNaeJnhAavbBAfquwzUV
zdiaLCzETOgYS2EwQjDXV27I4rGkOuq+NOvx47FiIVZ+4tPuzJCd6Mpo1sKb860/
56t0opWm5UuQWrS3wDz4uz3oUOyDaEUHcNUPvU3lrHBtkH50J+AQDTOoIJJ7xjW6
mE3yMNty6eEax3mvTklpkXhp6y8QRBP3onSEq6KKaDXy8E+hafuNSAdkzFvO8IRY
CKJ/qUmTAv6H3DOuzhoxHpsberT6i9St/LYCgESzsqvigSwTZMxREdPULCkekJ+a
lv3U22Bm1BCXG5fXCc3BprfOhyV4/Zwtko52+Otg5qAdaPRzwqPqh5RyWerNiGjQ
nelkMdONyJCa0eTeyko1JsSPT4sZbONAc7sFrloWQcGQ6yBrciLtqUjPeWCFatMy
Qu52lTFHtDPbyouEDrq3Q+WAqsJmyv+HNq1EJY0bwnTzS8np/5hiWF9OKQfaRXhv
Gdx5wnHpdmZmHYJWYnxWJlDdZSftaWoVhOnsJxZ5ynAnvplYhm9KUNahnaEY1MAZ
u1/1lgEZJdJqJTpy64yyazuwatnczPkRp/tfQ5dBa/H6ZTfrWDkvaNSY5DFkqiun
qDfdFUdmVk43xiRkDwcGhgyavCfwpGNU3/B+6LbnMbTZSaofDWTLVYS/AXPi0k/V
GFoAyjUDjqgy5Qrdt0wt/tIvi7sU4Q3E1ujeZwzIsk6LOqP+61Ju8MbGlZdqVoLO
LA6dVM8iIzurYNlDi+PX9DOrKlWoSuREK6dxTlqV1vykR6is0Ty/H6IzJT4+w6/a
nObDYTnKtbS6RsQHl3vQKRq4BOMB+X5PYNSW6CIXvz2S7MhIeGB5hgbgFqeEgofm
jeeL5hAQGxHj+7GsBUKkQLuPtbiPzWr3UiNj0Yxr9qvRogOacMIadVfDDjFk1vG8
tTDLRA6UcdmeCFrALE53wPFtbKNHQ9zzFpNDv0QNxCo0HNPf8iCBsDKyy3TrOJd7
R7221oVi55rrfLhqTohQleZCYfNspStR/XIETsH6rljGxjkIlCdGN9wA4+QdD+5+
jy6Q4TGDVpyGiaDNPxLVmd/0ab/PEuX5b67XijQI6ysc3/ANW0QY0sddt3ITdabH
e8C/GjA3EXwKocxHzdACBqYV6RdBNVhpWJltAXg4w5KpfDCZ9Z+T75IhNMZqarjC
fkWDRX8X/LbteEaUirnZpBYqxOX40IwjRoP5fPceyPSUqkgGnScihD+nF38R9jTR
bd6kkmt96rZfW31j+O2ABQ1dfQx3GXkZlx9nXTAQ53VhA02cSYWs6Evm366Y+wvS
ay0wPPZMMjuZknL9iDpyELaZBr1KDhC4Bs5xB3aquXJ0nIdcVSk8/Wy4B1E7dKIH
2nPXRD7Yhz0Lsc7xsjhBtjI2ySHu0AXywjDnUWWyf+dY5FD4alZ3Gezrv8risBT1
DsKgNgTYFY/naXzbErbu9PCUiJWU9+6xQ8cMdQhFU3x2wV778szn8R9CZCn70Ro4
hocSy1je7dBZQpnSgJ+AwF9ZeBtDsb3BbQ/yAl4QY6DV2aAtltjqokj5fQZvBwwG
X/EjVhdiVbMXhZOx25GymJ6l5EV2bp43Wpe3Q6+GV0JHvm0KdFFaE3NAu/81BxWl
UQ0BWDbYisd+Y3nz+SaMJTZf4Y9eDuBh6av+VZWael4bRm1inbVtyRSjmanhc6NJ
xBK59VWskTpBeFJdepURI92rnmXoUIGjgrDI0WN3zAmbkhdG1MiN8YORnrfkj42K
2H4TEO//FXQPpWOqTPb2SjoBAR/eX49OJ7belblZY/X2r85zYgRb0dwep1X/cKBu
OnTnfUE5MILON0LNhA6upwQQF3b8Eg7ogs0ou7TP0P1wxefxvX0+CwrAMiv+8jTQ
d8BE99NcTTLF210FXlEXVyNWHTz3XYIrRivO2khUVt/jpypXNgHKSvtidZgY9F9U
kOUyFbwV2+anBnOqpGhfRX4ZIu+Xh0L2hEttGvzbbvXh5S3IbDuA797SIvZongaa
UicUS9EudhRQpguOIUt78BmiB6QBCemLefyO1lqEfV/ranpkY/8jxC7DLCm+YGC6
CGRRRjedyQphP+blcMI339gzRO7lnpYxkaVs9xNCWwKIvklygg6UYNGgq+F7zLPh
kksO7woo2wfyTHAlZcGGq0b5k8MARAxzthlxAz3fcZK/k5aLtYlHCdhYGRPnsORu
sYHodlcwa1pdQ4vyrBcr/Z4BnH1tnLph6nYXnfSDsHkNOTlZlBvaa3AbXzKSNoRC
h8Ky5eN/HtDdhR2qAogyo9BNIBQ2Td+dN9ehXJ7aXPY/cstLXdgt2AmxHujjp8VE
aGpLhELLjIpuM0VHHxOGqM51Xz2uCwEswFzZaOGjF1tZzTEK0uScMhxNhW9Ag8XH
0Igl93sayhdnODXp5JKyR3klvtX53F3W1vrXlRcZS19LOLObLhnZcfzYaZzXLcb2
SwkbH5UPKg59DpG5Xa8GNwLn6YlpiH868CGlfMUyOgdNU17jVbl37RKKEgEtvPO/
LpFSwzNNLXAKDTjlcJaB8EVOKRd+pnEjyx9zu2gaHsMrGXHR6Fkx0vXq2GbNysOr
q6eBIi1GQxk07dlDLKlYM246srhQdHE+k/kCy3fjUrnTh5ryFtdMtCFjKBBww08t
CuVS/Y72l/QBe9JGzFcCbYmFX8YC9T7s9Hx0E5SYgIBNWKMqEif/wbiZ7EqONGgG
rUjBp5kMwOSQwYAD2jgHJmdd1TQ6NFAAlK8qKu0isNLEX0i8pHDsDe3Yw+gRyX64
PmdcePHsro2jROem4gYkbUgjOvE+RUY33RXglyXDaT9+a5UAFSWky42ApY6G0BH/
OTt+OCO89IHFpLOclGMYA6fn37/cICYM/ME2M4ffXK4S3w3KUjky2WTjLkp4eFgu
UBfW20DYTHrH/3hDWVPvnsfe/EAsUJdYZpAlGcUvdOI8JsBdKX7jhQ9QMqWBv2Cp
3eKa8n+pLl7jUzC3eSm4ISeUkdYI/+d2pJOOYKyKOz960Mj4RI5KPq5qrahwbevp
T7QMYWDZVPVbzk5BK4jGsq3xR1gbVZVlvoOPyn+YJMBMnO1z69djIxl/EMBI8Znu
/kpvofnC6CGHwvZctjQp+QHzlBhYqPE0EvIixaCRFL12/DRjw23VM/HaXmnycsST
bD6qVqh2uAyswUI/aE/2nxrblhEmKgEinHsraA2fDp7fQXSc6qydSEvgiTeBTNMK
tuGFriZrzRxKyARu+NYg+FzuRY8IPUZTYi0Vr1DbPxvQ4rN1I7e6IgiqgP66mfGn
SzuXWfSlNu4T1aSBvzn3LGWkpZRy/B0dwMT0/RyIhIq8tZUN+/mG+VMWM1F3VNgq
CwFBSmziNGbZ0nxMWvgjebR+rLe0AJneBQ3anwM5Iwoqh7KSZYrfbxln3QbyAYxx
BO4gZLKBIwv80Kk989iXP2m4OiOLQC6BrBfB5btV3USTuuxPXr0F4Pfq1z/1tlRl
pi8Z25BxbAvqpA/2cxuWP7V2GCd1FJZ2evpjcGqtiifFTjfOQ19KxgH3QR2FBaOC
gNdW3WMY05/gA/kbfepJCCA81FvG5u9JU6TCo55dC8x8ufT87J78ySIwrHPaFqGG
HIUDlJg+WFwasg0d49gsfEmyejd51ZKO/PQWK+xYAiBbD/a/VPBbhA+g837mHFaq
7JqKWDvwYqdzBIGOQ8fLKPWN/SMk46JjAB2CfcRQKxMBQazshdfAnEntRuQHp9Dm
7ZdaTH1sGY4vMqrztd20OuCMU7vjB/yDHMRf7JkiG5ijGP9mGKVw1MXxuEa6Km/M
0OuaScHFLUn5nx3N+GtrJ/HWlCF4UqRoPdnDkYXVQFpQ8xykoePvZTUE8mENPYLe
Rf48qf5swFsgZkQJnt5FLYrKFq9u92OYS9eDlm6L4Ux0/0efFI5DUba+b7F9TYtq
3dbIkR7hwqER8NAkQcwM1h+eSe+77LJmJerxpPmr2oXdLGUI/9YIP07OcNsBXZQM
EY4vSZdO/V8xp1CM/6yndoS9uD+v4IoY13rdZ8D1H6lJLxWFL213VuFQgbVdM2m9
8QurtGsSiL3cJ3Vb+rSzqRtOtf6bFccFwcYecgUyFo4kxp+jAvo9fxyZ5sp5wdHi
WGVX80GFViDI/MyR5dftn2yrRDvVTXoQ9QtgmPYHZpU+RsvLSYuQUqKI6b3GdZFy
oDaBcBWNI5xjQGy28mZDfdNKK62Zni87seyEHd8VOQoNjcgAlnMJL3QLOWJMtQ0U
6AwNWXfW3QHCYCKWvJDAXKVBqdr2Icrs53dIaE2yKIRC9+R97VaIB28wcIzHC7xT
0f0eQDVxYkqzHCBhrdnLaPHRzcWCWGjnzQ/eb0pBCjckourH7B29lp7Ghs01jkYo
ec5jiKFV0prVzKRnIy2NVqP826A4oqaE3LeSbipCdXHsYSUPwyXamJNI2L9lFtqZ
ooVWc1iAzI04xrvFONz8gCkzr4MHpLzQcO+V6LGdB6pJfMUq5bj8ZmtYnk4YF7+F
W2JLROvZ+bGxS/YnmUHHx4LP4gfYq7jtywzt2YUiNVpcgPuMaA2FJg5io6Nkx6sv
6OoS58CwZvyVqW3T6IG0Z3pKpT4esQChFn5f575kxOh8Erbh9KZCM9p131eQ1QS6
rFrJ6T0txAK14Ss7gdy8DGXQQatyHAWC0dNqTkZdP96sqkbDsDXXqdlwO8kuuie8
PPQnDgbsslNKx1S6Wv2lIVBOil6IM7pGwSGk6udogFzYZTKUHYcdd+XuffvsYE4P
4A/IV+iRNjfdwhUbTeOJrLsavXf6emCSGyxtYmTXPWQ7QUImzai7+1dV/7/+V9Jp
IAGsCyapfkVJaG3SCzLcQbKpOi/R/yJ4OIngEbHj/turWfzvW+J8pPvtM0eYAYi7
0mFS01pn8PdYtB+fWt1PHvBiGATy0LBXleHwOBDt05ubbX5nME3aE5scquRQ9R/P
5flhmEOTIql6Vvquvn+T9NSYFU13/EP0eBZwK72n+fkz4QvBZHPAajGT/HJ5dYUZ
SAJ9kzHftZMGgBWTKMrD/EKgUmR7f/7ZonzO/1GCxL6syas8V7FqBKegK8r97Kud
V8QCWNfr1PDbNVyb39qddkA7eg/viajvnFIoaF4dtKsY6Djx9FofrQlIZ/o4if1t
gVndV2O3wD/XbrDC2BQb3O58gK37T1zLxzxKOT0i9eGwHwWHe/hbKLrnVPtoOy2R
+eH6gP/n4j3UuDSnLdIVZkHg6LDePWD5rF8y1StYl+090Fxzd8bjeCoKcHY08qWc
Yv1gOeIwOkhIXD3PzlC4/T84c9z7w2llUBVKLFI/qBgkSuUmXgrg4TI/Ftic+uRb
q7rjG3KBtu6dkbkaKxskFF3rkrjZPD5+OY+GJQCCUAOycUP1fcjFRMcGnpP7BGxI
G+cTR6VrWaZtg97YFMgEogLIxK869WaZik855Axcm0FroHVogN8yBlua6e5w6VjX
3LGrQO1u/WkVbNFl3atfEv2Osoo2OJHvxPVXOeTvnmpf+xy4m9elTlJXrm/zWec2
BBLfvK/jITGaCtKbWW2rKwrzXVA1i1Nro/hFcquqNgOSQluDhHUvMvywN4qPboWA
3UcS7fWJxp5CA4YjiqnnVk568J7cSaUw7kGhQpx6bP3ggnH5nlanALyS7BicB6Pd
YzzKWOU/obzQ64CvVZgHxBIjx8FZvyBo+HbFRW8KnbUROFpMm8T3dz7HBD/gqOwN
Defl/yuSm0QmQT8gle+hfu3xa0Jqhou9sEglMAow2KSRqnRGCh1y4H4WM50G2u51
zEawMh8fELOndHAht3X5yR2a7KxHi053nkPzKjWLrPvv403f1VZLj52xboBJZyJh
OEsuXTZlMOq5R2hbH60LHK7yU+04H1aJBpWGWbf8eyYvHwIHJ56iGKSHzdRqCo9N
ZkYYa41/yji2EipIWI40VUGPgx9Qbtbga3tGqYSEfOd8hK3hCAjPDUV5AyAaNeKa
6dvCt6wSAWeipjYxYXFZDoed+ppmqo+ulPMVdwIqVKLSUMJeyNkiRVmNCuSRXepr
6WDoAFAaA2wgDO2hRTfZ2RabKaSSQeGmTx3EIgQYkbawibyd7PIfeEd4Ibif6gVa
IzoxzD0iGkx8cy4zqKJiiDh5iL2EhNlKDx8DPZM5fyokCGzw3k5Q07Fr/Bw21pwB
xUBY0gb0DIrpRBMhbjdhWnqrUWl93FoTW1WCE475eqGdOyEAJ5XsnlCYd/IiCC3g
DMCb2QLnwk+N9GJ1Arnk05CwJZQctUyS3sA2wZTkZ/PpukSU++Iv0IPPcDj3SXnd
btqv1epNwCv2mSC3FUJd+TY8x0+CbWOM/nPT11QZnaXzlFXaozClbiWgfLONK4zy
gQSZ8sW5unrDboxgXtEr+/J0y3FSg+WaVlz19LtleLi7gRahfFnF6VYSPiX2PT0A
YzB4RQr0xVObFTbHYWfAloEso4HKC4weQhn0Mhmp4WGqtt1NF6Lv2LDy0HeUz+mq
vuaBjmAoAfUiRKlgfpWfzElpF1eVLFSBFszRekNKXi49GCUWUqZyQa9q2DiLZmFf
j663zhQtc6sRnFMzs0AV8ynfQSYTYQeRX55wXHazGpgUtnZXUotmeKsTALG4/eJA
t4bhq1PSyE185umVAcB3nu/+MZTBDAIUZZK0smXVBEZWmD3cJuMfWmfiq2fm77AZ
BhBPV1dodErO2AVMJYmwnhgzGq8+Q0mdkmbHB6IsCZyjif+2uc98KFK/6aDEotyy
GTzY/H2lUGbQZBoA0ehgsz6poznhAqLg3s8trn9lJXZj3bY5Fg9I3qRAO3vuMaxB
AGFareQGr9HGzAlk/m8hhZgOR9eR5MLjStMpd7Hh8qW9UgdSFr1+hzouUQczNfob
R394XhuQXJXz59wqmOwWzPIJrnKu4pYaOXFdPW2vfJfxh/KSUCxw2z5FuFJFsNt7
UaX8Hdene169k4jymT589ZfE+LkM/qNdY6Z1wO44GBSmdA7e/YnycZKiGJeOBgcE
JUrgrl5IMfkZ3UysqPQu4ncotPA+WRfRr9uWtBOzygp8HAl453Uqgxpx3HBFHsK+
CpZI5PHub1PXZdgMdjMyHc7orxuB0ndqLrKhWJUKas6hSAuvq/8jKD0sAtuzLLur
JJhBhbkkM/I8HnshrSXcVZd1yQinihkcQIjDJg7EzELtUIymNDelZE9OZ6ftRmny
k47PWkOo8fALBJMazVuf5HhhaEv8eRSFwprTBUkpdyTe7785VFK6yRIB1HXIUVnx
+AMp7KVPoK5XwkOKTklR+etbQ5bY3vEf6zSumUzAdorMbFiqbDbhDqlMy7ZeC2A1
Y6spGIQ6HxqBmZweNqiM5N1/NSc26aTHK0ejyUQWI+3JBylOOtU9P9/DO3vZBowl
iDgQ3q/x9LBECDAb3ND3g6svaIMgrt4Bh13hfBJX0A3h4yOAmd+2svBIN8s6iikY
W8STgZaAjpE4v7KymG+q5KkJqYNjxz2bmRBAYj5El82hQTjrgzxX7Xyv2cBsxcLT
yM+QkmKiMo222BDfosOIbc6UcgjB8drSUvrnuOOiLq5oEbbmZ48AYSg4i+MgP6kH
2O0Hnb8wig7G8u9erO9nhlVvOyn7M4wCl9/6F3klVazg7Ofmxb2xWtQlBvBYMnxL
L00wCHSA4bdajTBX8C9KUWjqMg8rsQQp3nTIB5gLADBSHZ3deq25/aNIrl3or5Jb
HQKofF/NjjC0vDh+uWhiDBSmBVBA13WI3vMqfcGE7jX01rbKJ2nc1GrzL71lpMoT
J/ChwxkiUHc9LCD10eeewjKLS8K/p2DizggM1fTV1loGPrJy1gqeGGPfF+THap9I
Tv9J/f+KLClOQDpHrY/ZnsztU1SwLX3Cnsea6thoJ0c47IN6F61BF+vBMbB1mxYx
N0f/d2tnmNDmCKENOIme/oZAaY2SxP50QLV5qG8p+vZ68DMTGtOzgSDw6I21infG
M6lKE56fyPy0fR1hlSV6EsYmk3Jt+yFERlkO4Lf/6zf9yb1Fy5M+uN2EOzUjDI7g
aF/Pydy84AeU+IccDH+dHx+gEatQA09D2gEM3T+AROFLzSJHvlMUX1dnuXY2VQuT
220WQ3EQLqmKygU/6RBJgZvgnFESea8xGqWEO0dbKauITvyHqNNHsghJ3UqePdTa
hNYT/WrxTcS1faXLC0LYi+wnwGujRiiPjai/lpOQISs7M+abzp2pNQ+dqcSs82RP
Oypq97UxRjrwOA60MjiimSjAjIJFEOv5g1ifcCUPHUC9Rym60QbbhEgS9qO9EqvE
E8T1MKjLIaO+VTKonaca6eETp1Q5eWuoEZE/RTZ5jjReF7FVn9+qQvEQUXYg6+xp
newmF6Kl+u5XsGqmSr/Ef0hrmIf3HFyFyWDUad/cAiH7cRoKupHJUnN6T4dwX0bg
N6gtmnBu87bloiOgeWZsH5G9+n4f696vOf3L7bczMopUkdzZUwxvPftdg74ja3Bx
qJajZKJfvheXfpA/lBxDDUYkyfdSO4MzAQb4IbtTKeo1PDyZzv+8tDxS5bA17Kr3
p4jEoDEBXKxiP419MKmiRfWvkn8AkBYbgSF6kNjH1B3b5axcc5Kea8tJhKs2YpuA
UlQawdWtQTzq/VzLY2Xppzu9q7wrytWbpWe3nU1pBIdOYpDQRpPtfmeLa5kcKxPi
5qchHba7zQksTNvU0rBqrXrBo3hWJt5aZVxvpOYZ2QP7uXCDVj/BQp2E8WnQBDTX
+6mCwgJHrFaHRLsx0nh1SKcqGM3hwRSy8Mh0HPh3QuQfQSvD7qIbRZz6SYR0pgxV
YojybwfE5hSsUOZcFWDJAHVaPr4xPYuCeIJuus+krfk5I2G6a2nGvbqJXyz2t0Dj
xHwlNLPagv55EMYhY1OVbdIBL6p++CHjzM+03u65/cLk90qrJhjT1axx/fMzD5R7
VzMb5wpT2k7N3ZylYOHMrtxhXR+zmjWwocZ0afvKvq/roSS4uSJt/ByVeljLrByF
ET+SsMN4tTPrX5fy5jyelP9EpG9e/yddlDpPN7GAX0ib5RSI7tQIjT8uZTSgfSp5
stjojumpKG9Natx2RPjgz/VI/7Y6kEwPDdZzXv3I1avj9H2BvJTVmLf0zrENQao7
Ph7YZEXa+H+mx1EMOlaoEcwKtWs7XijNhN6lixJTOp4ijTeEGxZbtAAmYZbeD1T4
ZZ5KqTfdX83dm4/VJTOwlft5vTUHZe6ep5SKqIvw0kuur9CYy/8Fa4r3GODsi58q
cF7WyW1M9+nogngJFtv3SgQi7bBYIJ35//KikeoGp77a3shfPwpYhneg1CZklKcZ
ejBGSZlAnGF2BkNpPqpCo5lD0uWJv5qulWFWagNAoxW87i5FejIFVskm8XvjmsSL
TGoKcu3Ob2XV44MxYUikr+9nrIr23aZ8OSIiV8lDDu7bxcyfMht9++SqgpMjeP03
pAtC8CHsyUAI+bE6BEbdReH4Yf5Aw8b0jNIUtPDulfaiKRIuNwQ/KW1CIdpKq8+Q
sWTQi1zWQT2rlg3ybzAqTWADaxaMk0GH9JAevAkQMzEUGByKgXUHn1hlo/sdiqCC
ChIMNZ5BQoJMYXXLL2R/vdu1wnO+MjrEJ4XxnaEs1xubleVA+uRr6SpxB+lc9Iuc
/UkDCir4UzDeNM03AxShr0qYAepy/5vZl3Vtdj180QNcfx6pcJS63S6/19mU8aG/
pargXhkcEqAHqMjUPXHqHoY251hCTpp6ZHb2PB3IPW0BApl2jSfWyiDlonoHHdKl
vCH/OE4DfHwtqEOrlcfh2CNIakKoWHfeFY3YWMrlccxRcIofHwR/+E7M5aov46G9
+A9yNgZBjPJKRYzjkgzgptyZs044bfM4qZpU4pFWETug/bBdNvZhrZ54YTYd2UYy
QTIEs6DEdEOs76FCHfUAP7e135HNJGKhnVuLi2MhTmoqM/dE5mByfb9JmTr9xNlx
TVE/pf7m2kQkLNcrfK6ETJTuta8coCYBqVACHBPcwAuzu68gR4EI3mgT7pi0IGIG
bjYWIkA+I+zeV+tSRICZzSWbveePQj5lkRhJk4ofzO+MosMZl9hdLk2PmVoP9TAe
/0WuIcj/uytiwQnInJIova2DiBCOnmOS+3n1Z7e41PLHnIOQDH8f1Ax4syRPhbOM
0tm9rKgMQ76lYdVA9mhl+u83bOjEWwAH0ilQEmIRovfRvzACGke/6wdgt8SFp6jq
W9dsRCKTToWbFkcEaWlxuifGCwVzvwVEZ2ufDFTbrgr0kwCZALA1tznHdn4b4z8M
JwuNdnnnISqCiGkW92d/IkvIqAOXqhFjowIIvY+AU6BaPHvAloJH/gmBepEF0fdC
Gxiw0RptKdmb77oyg3TIhxleyr3gdmA5KjgwNEXRaSOxEqQcAiX8uS0dHHeE8ul7
Tnr8Hau12mHY70Mg01KxFJS0RkYXFiPtu8OsMJeL/jQGxP91GkffBpoWEBHqUZbc
haxW4PP3l434KHNsNExjEeU1gDbnHU3I7GTKP0VJtzXvT89dsESaqiSD0EKPcLAE
E8g4copRcZ7dkvNf+uufihiKTwH5KtRiZISuJ02L7jYZQvDOZvpLPxTDwp35MGJq
r040GMmZaRmcwuYUmH4GRl2ti9cJW5WbflTik3M1PVjmVMW42tsmWVkLTEnuoJOk
/okHpWkj1upbiE8zC0e5v+UC+WPiBoNrFQfSfmObha4U40cG0PFo0T2YaOKIftmE
0keUoxO/m65/g+dcDlMIIJigq1SDwicoicnSpbLhw2kT+pz65P7zlWdpZJg8fpwH
jeqhqKBGjvOEl98QS2uF72ZSRZXRfbJwyhdqZLC4z8x795XsaWv0WcUFlOXZkIcW
6H0gp2sRs0FwshPsxG5yQaOyxTCxu7h5UIIzVA+uG17IV/1dXWH4pDlxXkPZvWWA
1wtsHC1DHrSLdRZp/m1+RgPFE5t7HoosThZkKOb2EnWh/4JRUixOAMXjzxLQ09Bk
rDkUgmLdtQXcKs9fVIhrSt5Lfyb1LACIgC57O81sHaCoxYO1HIN0UE6+KDAuSQqM
tev4Lm2dM8ACbK6v9veNLKSNbSLzKxBtPdnngHi79o4wOdejHKWwAd6TNLocsV8m
C34VRXsDF1Iq4Jrx85Q+2LDlz21yO9ZObaZfz9vfkOhIcrnD6saK4HdbtfyKd/SF
H7B4Q1diE0k6kTFEMAFZymK7GiDwoYPuRukNMYl+x+TgdFbsqEYtYBI9iBQYwlR+
Eak9caE0c4aMCnGrDFpFu9GDjqLGnQiLw2/jNMr3WFWouCcL1ZcF6/fI9lgdJQzh
pgHYgIBsWZB82Ztr+SxxPYZC5+WOeuelIDxtaycl2YcFZJr4R/YBwkVmofekyTON
u7GUZkYfegefopHVOGYcnannQQU0qe3g4rFegt0SNNOrmrGxY7KXjMUvb3iQLeF3
uDqvKLw9M7vEFpVTNMoDRC7q4tAHhn5xE8TbXh70ljGDAKlz++aft70GPhbdOqKl
ItYdKPac7UrBfPYbA9U71nLCxPdu+9ZGyWqG31HzwIu12ZyWUZsqgP/08P7c2f4e
9YO26whTLofPlRQiSHAW8ahkh7I8GhA1Io3/sF+yz6TfHoyewwtd5GXZsv/24b9f
usBkbYvVletIxjkBt5eT0nGkPEa5l2cp9plRlUod0T5SKXVHNLLbsSzcxn2eF8TD
FI6+g3LJ1RTzcTrplVSi+hEpAI6/YQ++7ER7DsX1RzulQw5pdW7zaiO3s+fZ555V
Y6D6Jho6dYwtkQV/KCzhB4++QSbHNZFqLls8nyyVZL8frCDPR3gW/B41vy5QR3qh
DH5Az2CH5zjc4yQoa8gBnGs8MBzTyXH0QHvkGNm6A+dUHDI8cfGZ3RXAESuO7wz7
MT8nqrTM4IFo3boo9tYEoM4SfnLzLh+lmHnN+QReAzuZAl7WGLLspdPU8sUApt41
Mn9FxoxVX+Oat7NzmNvJlJa5Llz9vJCpxfqVWADbqMbKw3o/tw0/qsrDAcu4Ayy8
f+QIVQ0O1M+3aJ1P3WbhXvxqDQ8RQqKDWQiFmqpuUGwyTwLq/kkLZRWDKmzg5Sfd
q8u5K3AVsVABpG0icSW84Tod6f5IdgFgcSsRSP8hJmRco+dPODV8HBn8aJjU0EKJ
5RbaIP+viKrD0nSFVuiiXMKvwFRadAIBafYqzr+JJhXiD6T2A8kH/RfDTTrG9I2F
UuK5cS/8tzejWJeJO45Zb9Lv+Ck7FjKeS180SwzVxJAo9RJX0MiiX8zZvM4K5Q4B
N65g0/SvF0AmfKP/Ggl3SnN9xqOmPRSo0wbxSLdaQjpL23W1HS/Hnu01kz7rH3zL
YkoJkoyKs75/NZG1km28u/Qo3hHRf/dTkLw7/xwHIRoQxBqYk2wQc3l5dyESr6Vl
nWh6QUQDAdTUQin8e3rglcz4GyunUwakQpZcr4LWqwwA9X+LKEcW69jz7ONXJtmq
2mj5T9gQpDcHZYHaqny8pMa7+vhuxCzo6uSy0qhYXf1HYE2+EFF9f4H9mPOB8++p
rhOXbWQy+yKHIc1mOiFMaUXl6NQZjTflcCjtmDcM0p3z0+kWQr/ckYzomeBtaGS9
68TKZ7UZWlDb9MsTGQ+KGUzifFsPUAycbSbsTKAjOVLhonifN7z5q2OB0rj6SXnm
Ivh5vJl4RsiYwFQzc+FlsE3MnGtPlrqbWgZu0Jdg0dT42U0v7V0ZOOJttnQNkc6C
9h+mEP3XIFJmq51h6o3FFM9K69wupSvFFraePagi6AoNAj+l3aTGgswTDHnYlvZO
y/+7gSkJp2wmsOCR5oKAG6+duMgnXLWyritLBuzgrYHxhuCqXvhsCCztbvSKLiMg
e2XJxS+W/E/gtESmnPq3bWgP3QDqeS9blNf3H0JStcancr6sqzjTv5ZKiryfIaMA
9N4wisL5wyti4HZn0kVRuyqCg92Y7jMzoJo3z1fJckgIDmH0FG0MJfm81t2fy4RC
S6L7+TJuxNEghlnKZ7Yq2fHe/+wF6TqLDN63SDY2f2C3hPn2SL4U4iG5h4KXgRsL
3iuaFM49CC8pOi+nkkUNPriDL/c08SL7LM3pBcRO5LlU07qLGt1BVh4HAv0JQuXH
GTo2Y3twprLlRat1xlLBDBddkcAX4T+ZiqCNa3yEdaBMt4e7O9mrYAISENMHrP+6
W5ACILNwoRy+yyWQA9QKAFIxVofCKAkzHu/8++WfPBccXPWdHy1CfiQZK14VFRu3
82zEBziiTgv4wJ6nLyodRkraO9pBSwKpooZ0p7k6xoX5wCkRDJCuVTyy2ivutkT5
MNW3K2WnBfbpiHNEA0eC/2/EltDamPk4ez3r7A0FWgg4xMo8l14CBLnFovFvQEMB
zrk4WYM5n/jjNa7yoaJV17H44FBwA0k3I9f5cEJCFP44Kx3zkNFHc9b8BNZvZ6Kj
ljm4H6KJqAykZJNbLrJqO5CieMxxVxjiXITh0g1XJDcPLoLojH2tW+K4EAPANBaS
FOkGILn2sUF1Xz7JSawvVSofGvewtJ+xkK/MXBuj1eaiM45DYEG8GwindNtaibjC
cXWH/oK8FiLSQ7EiL7XiyQ/uxX6wx0K9Je4Qksw6iuuBWIAFbbz5xoAdmpRMckrx
hHApAPmPo1W6iyikN22rjwrbsoO9QsKcBhHx4gW/TZE7748WqDxsUgH5SSENbjwA
BdXLlaKMKEON6UpVpZOfYOJT/TBSw+K+OU7vsSWBlJQ0FtXTXhqoHyURRtgwDREW
1QGB26TObzn4RquBwN5fsXE2SVUZ5Itz3PdY6wafh2WiLUJ0ftZAh/7YQGq+A0E4
ZzZY35lTYIIjYnhsT9Kawk9BEujX44UbicezgqGUF93hzp187Oj9vXnIoSGOx7Y0
gTvyP5AwPaTG4s+tQxvnrwitDxveHelz0fmcj+A7JOyiGpXFP2zIkReNnzlMLfuu
wGOmEo03mvTMeAeW/fq7LDbHEICotAcR1bfBu63w99pVG5zzHD3SzLRs1m5G5SiM
OezVkKA1l4tzqM600Af8BNeHdQb936wreAxqKbcnTCOgM2x7T0cm6WkgaZf9yVxu
WZwmpVvMU/E3d8Ax+DkHwfKH330xLnSOnw7YRHzRHr6y6E7x8y52njJAFrj5nmlU
68zqbEqwGI6WNFsvSq/WYyK1i1o8afy2u8XTdWCTGX008Ybyb3nWL7P5bkv4EqYc
G35DGGywpdbdLjFa7naM8WGtxIH6pIgECqhAerwxHWMCykIm4iEFcAX69dvIE4Kh
M1xL2diFKoQyHDhzIa6mkF1rSXX2xFnDzCiRVnB7YmbeTil3MxOXZzDT/5dfWrKW
LnBQlELZquRGOfpqDnVBq1kVCQUl2iR4ComEX3yDyKYpiBnq+MO66DejkuhC+3Ft
yiQEBtBa8I0Zl+/is3kGisEl4vMfGhqFndV/F6HlkqTfnipZGk/zYqRNIWHDSJTj
g3NCR1J4Nm2AvgGs+SZf1I5AVX8wUlkRQdV5BVJsH185gChBIBqq4j/aa7dASt47
y/JQn8eSQEL6+4er7pv/Rxdso3ceDK4hZgT7ajK233rJ+ow7o2okP0kdDN4mx4Ia
vFR/LihJ8jd8w8fpDc0aOZkqaBjNJpYDkfzBchuKmaekjc12oBSHThtiJt5tnRUg
G1qdV0dPgS8dUGtPjEioKxycbTDZCq2nESq2xOFoRRAFUAGU3lLVwRaMqY0OCvF7
NomhVT/N58SmI1FrS2hO36/KkjTBRU316M2sfcwMtLTQQ/2MmjzEzd6r0TnZ9OWZ
tYr0sdSCeqMrMKKxU70eve+bklasw3cRVcQn2zrW7q24ed+tQJlSS9HcocbPk4tl
n4W3WZIxhGI/2VlKhvxwfBcCDYgIOJ023+cPGbTiMr9J0O77aDo6i33bq9XmjIaI
B9MP0HIkQSIqMfxGBp2uV9tJ1r/pmqHtTjsJXIrOUSgGUp02PKcaoQOn8QkPMgO4
BxWHWvkzTDWvEiJ/SH5Ezsc7mR94EgIA+HRpK0fcB22Leb+dJJhALHq9mIuGX7U9
Hu2KTyM7kYL2CQ7lPuRCLma9eSB65Ps3+nNSiImLZxkqtawrt3WKqVi5yZuUS1GN
TrL3yALcJqp2k/PCtl9BiEBn0RREohERox24UGwRgQDUjo6vAAecyokyttWSgCTF
dHdmRHVbh0VsW/ExHpYFWNGQ+smdJLTdtGdEnDM3gPCtkfqwwKIiTqeBI+OlLh19
2Fi/F1ebuRK609Yiw2AUzYVOoiqzXARz6sfsVXW9op+OfUDwBGOWjc5UJAT9MnR2
wfQZaxgRJqtWtvg4pPUI5yKxL2nVwh6v6JvtE4hBq2aCDnlY6J5uuel8Cdv83bCb
s8/671DFzwMMoGx2rEOoYp2BnwH4l/Ww72+w4Ej2Q4rnFKOkpR6re9O7YskEdzc6
qsQ7YwQled5TCQ46OBU0sSEXrGKjFH4wydT+5JbkYw3ZwW0Ki5+fqGTB297ao+BJ
6mvas/FUW7Tqc06L7RfJk0P5Mk6NhFL/GcelIDFjz8ZMbm7KJ9E2idbbu9gFnjcr
5VQzw0yOMZQvF+OycxuH5cH2pVJkgoZny1nTOP3fwElDgnO5zBUWzn/yzSzzk2Ex
TK9Sz47Hq+ZRVKisfUTmBjDx+WnMUvUAhKmhP9tS7E91Vr0oTlksPCVcWUpX5iQV
vBJ98Ag2gZ4Q6aT1hs8aPpMQysr0XlFS6Ivd6ZzT5grc+YSqZO1HwlS4aX/qG65f
4UG3er3jltPoAedI79JjhJYXHBeqtLuteTVzQ8tSTBjDeURDECToRQF8Yol8e0hm
9ChB1kDZRC95Th+PYoXbSy7wcAD49/9ozqPHTypKvqK/h7rXiVPfCo6EUNoYG1oQ
1uDbH+tFRrv2M6oVem2+ZC06RJcvS9HW1PFA995qKEJ5dqjbiy41gcSQXhBC4xHt
DxPHziTf3xzNHsCzP1vGabxUGRGSUaNqOHDCrD5unA8okMuCKHVQQsWvUrxPxeof
1R8rCc4Do1JU4fN/jyntJRSC56jgyznNcIEdm5Nreh88oOARIC4MKFspjHr8Tyso
JH+coqLEse76EKHpsoDO+zaoktzDWsFrNWcluhmEWXUP0MyuqZMZsoXN6YUIn2wp
ZjABKtXBzT7M5A9upJqxidpZc9Q8dNUWPkN7Fot16bT9rMSHb/VFGn6HidDzBYgq
W14nm31dzXBSleTFhcWL+lg/L0ZGMbcARTJCmxc63pxDqSir/dURv7eNho4YH+d8
oRyYkWVp2lhOfVg2nV5+rxK6OvWVnuc+pEw0CALIDLHjdzF67d3iVWh7DSW1fnFQ
rEZrjdbfYq7tW7DpUuZRLhdYbWAjAznQDjxw12mxV1ac5+hYSd0VOY3nwT+7wpbe
5yIpf0eB8M60pST6R4s6B3FU0f/kU9ck4xkj7opC8Kc2+xMwBoahG95ZusfSp0Ru
Rp0Iwow63fhLunxAzTURO08M1Q2tz1VghVEQ1hUV8xeo0UkZVG4qd09yVt4uNFJg
Y227XyV4oIYWtGcco3qTk9iI0PJsn9tA3se24m98Y3bRVDMEY7clwppEx4W5/ybZ
zLdcqJFz75ruDMNKKg9GSAqCoXGZv1UESr1Gi0qeL/l++9cOp+ug5mM1FjflQT0A
fsiJV5MjjZ7TVqN127NrpwsvtO5xDpFj//X4D+2GfR9fiCSlF61uU8YOxVOXN81Q
rxxIz4wWZrOu/YaEPwEqJLGvoF0tCEEHs481Ed3Cv94SxcDEbf+Mksz+dp32NUne
OFDOD6XcEs9oJcq6TaS8fzV1mdZYLETAyJa0OPRxsiw9kOU6VKmgY0r1l9RQN5Ub
1imBNZKpqee9S1YmZTv/vqsB0hOM117AvU5sGo7cKUWIrfoPC4VpwytFXTjgQsdt
WA/Y2t6RyugVI2tEh5as7QN/UGmqeMPXA92cH6TF8fWPLPS/ut1mGN0ZGGH4Xefs
aOaIt8WWbeTmIc07dRp4xIenffxSWRLgurUWlXusMWmvXTk1q//HPF4MELXqHm+/
9lyHPY3qeWhfbZfE7Hg6544VQN37qm3/2voXFzWrPRvZqupVoaSkqvAAgjjemjl4
LLVABy6u7IZVOsOYnh3mLPs1xSQ+bVp+LhtISjgXhW1Yy+SwQkGe5yMVVAUS7/Tr
aQGk7DAAVj2qL0OJt+l5pnDMkFwY8Qlz/kZof4ZrWbRjbeNqUsT6b7G/YolZTLym
y8tiaKWSxHdWdjJRST5lDvv3v7YiiLEeVPMaQPSuT6oX2kfESieKFxAL9XNmh2Hx
LXEJYBfUPj9jmjkDKbO80mxAXlJTh2RZL3YrYldbPorHI/41p4EWVc5+twW1BtXe
qL4il+1xTrD2qLbYMEzvARGDyFHKdy4e9P8hnjS+frg/Wjh853L4HJOT2ijBBoPB
COwgDiQgIPBB0XshMtNZf2DAhq25xtd1eHne/u6A4vIZMsdAUSyM0TePfherkrsJ
/0yqaqZEqLz95lqHrwOI48i1VGUpcEo0F1F8QmxG23Io0HQfrfO5mgOBLh7/XPLZ
r3AKlJpUcidQYET33rmV3DJf4hGERKHgoyri39pJDv/Sa2gP+XNIst6ldenb2M5J
7haTBppUchyrpPvsDUQEIWL6nLoPlB5GuxmeajB78nCTMzubFRxeUB+C5SMeaue1
sfNeGr5vFkEEhFw8rkljFpGtisG56E6SD25nx8wTpoSmOckL0/knJS+/4qgaInyd
hvypHCO1A86jVySOuw0TKKcTG/Y013Pli0N2Kj9Ihh1YqH/GyZtnX7ZgFYU4W7RF
IDTOFYIMaFl1Vyez6aqT6qVH7FPrdhmtiUj6zOzpKyqr3AvePxYam0QpfyacT/h2
6VeVGZJ7iA4Lu0GcVndiTsq/3o/Nf60KqloCn7zrk8l+4egLyL32qrr9TKBuYeMz
vcziEMP0HNCSNb+smodr3JkJ3XhTI7OqFlrvs5fJNkfZc/qZb7st82htQ3KrBbX0
SpN9FbXEzOd4iOomz53g0MjtCF7M+Ns98CtB27a9emqy+qEN+mUle1twsslUG5VI
HgE+N4P1Koa3BHCTvTyLl7miwSmaL+dDbUma55G8DdHASv+CvuBdQV/LwUI+WoWN
P5XZPZGB9SkOXXHnpDEHYvtVFM4Ihq8/7FpPZZKuOr92U+FYlRFve8Be4zZtKE5e
BS1fwqmF+XTRThVAu/1rSu4w3LUXYW3oizL9mJZMk18xYdIAd/kP90o/liNqQj2Q
zhfeOMfG2X4WD8oKff8s8O9EQWJeABfINaD5XpD81S4sO/D7nXvRqiksxBqPdtBK
nLSlamKtwtUSkqmpe6SphFN8Zj2TYVMVd74B96/v1MdazcEnafyRYjyFRb+mgFTI
6yKj5iTCQXOARKsNUwea7C95c7DVKEUDkT351juG7qR/4Gq2f8n06i1blqpLBQqx
jo0VDckD0U/ksCzt8/9SnNmbQyOgJs4Bm+XSOU+0PFnHfJ8ov4JGwkCtzfDHjyUs
dWijQEnBeww1awvhS5BhMTUkg/R5JiwpqybplVR4oUWRnD942EuXE/WZkVPtLC6p
tzT7zTV18eEEvIue+1P5olMR9xQvrCaQ9QghkSxeNSygwRVlDDhzaNzjAcPLeH+z
Qe/pELxZ2X6b4LPyCnXtQt5yymt5O/Bf+nZaw4ck+EPmMBw4uxXFbGw2hKw1lZ1m
cWuHL/9Nr7GKHukjUZsExuXhQu8abGiqBATXV6LOCSJvbl61bWRRoIjZ4XyExk8U
VflBU4Jzr5JvIF5q+doywQhJqyH4csxPDMD8NQPuyY9ZUbRpyMIXU2eZm2XT3O4n
m2s3LljoDTAFL1Q6gOGz2rVMgydr1MjWL7WJkAhd+XT23VtvoVhtfyd7UQVc4izg
lZr0Kygv/Tq6Ai819S83sEcGKJP1tAFqriU/pCcoyZtBnau4tg0MjdaTzhDjkEKM
T09VJg9nXgQzfaDch/xbOHPrVcigqIwLXzdrBEAC+jAN4PhqCgE83JsHkhZ56I1r
J3u/UtUUUyxLSZ8yPOSHetw9yaQEJTYeGGvC42qyOWcNVeHlpyASGX6vf1Yh2ZHS
s8/Zy+Ivz5VrvQkonRFetVzAwKbQOi2gutrt8Xu0uHq3KdymdBztX9Zc2Bdj6awz
pNM4QBOwVthdsso5xVjG6V2zxQiz8rDaJzycLpiGCyNMPiWMk6bi/oL0EP5c2DRr
0KMoG/ztNn/ZB0wedgALYDYSC+UhoQGuuayPDta9SXT4tVMKD4QhikSKJvbnH12M
Mgfguv5FI98nY4+qEQ+6CptPGdiNOZSr7g5JYJsne38LhGdG9RL9dNls0XZv6A0I
dS6FJyDY6Nz7YHdNBhKxTiS3PRi+yw5kh4N/CRSCfDboUiyF1MovoPIOKjqHEZev
2DH0kkT6u6uvoFgMMaXsZwJ9w0HtnphmAkFXhuUL3XWX1otUrMYrLWa4+y3uaHLZ
u+0S0HC/KaMbGpppNlRiFSrX+5aOgFO0rR3I7aKQ8Oj6OolrWTlOF5ZAMU0CBtyf
NPOt6uUWGVBsIzqTMVEsd2s9FeazPmuKODAIf5XNKba9JclbFQlDquPX+tUluWJ+
xgvU75MPmmtwZ9P2B5FxTVPfd1hS5CvwbCPS8FYn26B8/qGTL4xGpYrMcFjSeWtx
ajFZ/hb7Hz8JjR/hGtgnemab2DK0H8FmPEyFsrhsECia1UIdXArOtD9tPhvxLp+b
+z+aeg4702bJsOJFgiojwwuRvxqOUGh3Oaa5i3hn0qMKJYIQ7NcbYV62u8tdl/dB
bOR/aO5OtNR4INxFYjY+/3+FDM0cS7SEjLRtkHNets0GxtY43Eq/k4QTZb52SIUW
bXlRZNZssZ7GP76aeey3IVyAa3jUrrLSALvGG9AZ/3WY6NTdKBxDyhpq6G9/NNGf
X3Du4D3y9013XAcx58sbBHh1vRMOF7VimT8JDnXmbnhtnb2m6xqd9JqID6z9JCZE
td6mTDdprIKiRsX8GIWHxPqnzm2IJbiLdFmpdQ6D0K8ECtPoSbATwY53cMnfJYFU
JJVywCkCxTQeQLA3NGcpZ380s9dBM/0d5S6NfWuqqmTFZ903m5rMwaky79ypjjwF
JuRkSSRlWZpfort51lXYdl5HHeyG3REx1islGjfu15plPCQD8gORx9XKVAbHemGS
OwFecI8KzgQNKDA2lzHTBEX9Oq6QlqiaFctDMA4MRm684ZBu02oO45tr0SvQ2MQW
wNQGb5yXYu233ntr0mJRXKulpujBAWQNM1TD9aSJMetogyYk/SicIs1rdcU2eC78
/MLNQ/ZXqZb74GdOyVyi/ZgLRb/riMfQt+o2lEBsi2ImkkomfBlMkvliVFpaqZEN
A91b9TrDLDd9AZy8XBaDLEe8thFhF3P30SVu7Aud3GS+592egixZ4JBX6ENa8vam
Pkjv14lu9+TfKgakzSCEENLXmGfBjZod3OomuTNjbrBUvg5ODsdx5RH7Wz/caXun
bpB+TuMp7xF6k2sR0n18eNuOTrM/K8JwzRScWYRoGxWCu4w6w3E+eeOk4Fgoebe/
So67LpQGEZyHw97x7xeHypjs3tMUVZzrdfPqllLWdVe5z95nDoJ4NHy+SH3nHOw9
iXkbPLLnHIVAFgsOy0Qw9KvvfYWf0o2Ba8Ct8OVnhHfWesRpwyUidFdMnUVmi2W5
Kt1DhsqymlukpJx08k9dsoHv2TQiAR0Zv/Sb4k4v8PMxZT6b+y4oXO9bffkRMMz1
YQ/7ux60uj7cQBUQuplZuA9nl8c1k5Oc9vvuckmlh7Qz92thdZfdNCvlqvUtnzWz
3TrtlmZbmahnnwiyww6qzgu1sdErzS0Md7XraR83OU33nK3iDy1d/rVFqNmNgKU4
fCEq4vGxYaSPeHmD7elSoWs6S0mQ2OAk3OKFbc3apvMeOqr1bylPByfmEVfi1e/f
ZcX7i5UtoPin8eMdKxDHV1lenhofJ9XC+L7jzblNg69NP9Z3HyNFLzKG8cWhwlNw
mDjKrimcfD4aH0lCVrNl67W77jJhBl+0WRbIHk2gPxj0WIkeOQ0xqgoVyFrRpdDI
Nw2vIs9yJygIQ5NRrWRIiGuAlRBmc7iMYDR7Mxg/iPuULGS4ltTbkbrUT/DmhDYh
IdZ/SZRkj1httphDOE67c9Sj0CwOVbHl//NVtCoDC9tACuMe6bGnh1PqcFuZw6bk
eNWOcwmEw8uEucCga9gForvcev1Kif4p/K00OSAsX0BCQa5MtIAw+L5BcSIj0JWs
p+5QDqP+6vGlNElVq5dxAjsJpjkBmtO2Dk2tK+7jQyKMmMhvmPIashRIG+gh31JH
E63QSfKlkE76YGeDig0Wvt4rH6MeLUn0s8C0HctQT0oE4OoguBh6uigiQ39jIsdQ
Q0YtwZgWCeW654nxsby8fCcMQxh4tkk7VyyjCRjMWTbmJziGW4yTbFrdeOE2F+qV
rAFaR+34ca2quFb1eaS6oz7EhRxZc8pAIvnW5x+V+gmb+glLlhwuDopBqq1O2PAt
Y/Bdo05XxByxVsJuqctRTsfbLtu2HD18Lx6KyjpmW6RlveT7cADp6Mz9XntwEfQf
VnrfcQ/leFbPSekC/peQ1Srm04vR3CJGU1OJvAmQdUHyKBYinmf82o0cxi9ZxaYI
gRldp0zOSEc363ORj11wcYKB1iiv1P4r5rdwaxbfgM53ZOMoyVsy6gVH/+eGBPeC
7G75jASksBEwtsPxj03KHha2PdxlUvAkX9bwW+z7xGlGYRIZeTYsBdq6vgFRFWZS
+ozg0P4FoT2/XfRp5qrpTPSKWeR6DkQJnvB2I54ujxLByLc1n49shXV6ek9e5P81
Oh3BhgOK+ku5vDUJ7p0GvB7YR6Zy/VNBaaSLMuLU8ZLbBJ7vsRJTXvcEX3DLq75V
+0HTRnFWsx8cup4Xq9seiUoz+K+3KNCclDaCJBSakLksDRS2Ch1X9mxE7s6o/frl
E4cWDSSngQEdWjMi/NEW26xnnaEHqaQPexRDoYLDLl2PaaOkuY9r4AzVZb2ijLaw
Srkk32X9ntf1a3EJwoq3kUmkmqKVZQzLt9vtBPCL/y/hyeboAN0n9ChYafcxC4On
a0d+jJ0K3CwxjVfg6B+hE87DaiZFMEH/njIyYDPv1XlxaJhOLFxZQtTSh5+7P1tb
NrHAPYqvpMfeou8ZOm4e5resbY6chmToflhjLLFm3DgHPfccLsA+p4usdoeDKi38
2mVA3CnlGH5IjCdEASDvAlvCmW8p2DGi5kxuV6cMbrIfhXE4vcm/iUtioN+lKVOc
G2WByNYlUSAkKtzFIysVHO6DH0B67VBwNUjHYMUi4jFdouFocfAuxBW1RQ/ycIyR
nu2uTUAZ5e0ZCfuZC+UjSGMoZgZ3CGzYDn5oc3muUB6IMNCykQcR+T8i++1l5Agh
Fxj1Q3rrNd0Py1X3mmjHxS3ZPkV99UN0gsVsJ1Iwh9/hTP8uYIkTqUOtmTJ9HGA5
cSpXhQzPO696GZZTaUHSred0PegSHWxkboBpK/3/BlHFb4yoXE/Dljw4pnt+Lu/8
oqmBPwELJiVjU4s5cQ6Vv/Tn1/HDtBtpU2DgeZa7G768M/dHwkNlyOtsoorEQBAX
XgNKhTyBcgGaVyllaps92HmpQ3KEY14kBjKL47sf4jmWFpyA9ISSXhd7ndbiJJEW
7m7hXCD4H3hlBcZyCB3JivQE069vxHhZ7S2kZmoZ94saUhJxJL0p99y580lssjFG
HzkU/qKIg6ZENxTYwO1AbBsr65jq2rgVnFE/Xgk02/CyncA+0KNaMOKeh+y7d/Wl
GIdzoiPtA1xK2yIAiBI2Ssz9oCnSmpGlM62xIZ/R+QTT/fP1Vyf1KdvChDcg1VQq
tHC9fx7t83GXOxoYtsyCna/JepEKKd5SLTThktx3nZHmEYWIX5l/kt6G12pVzBbJ
V473GQP9pgU+O+KosYrvoT0f0fdjBn+cQJl//0Og2oz4gHRVl16HHF0A1ROywGMF
v+4rNVFoUL9PfiQHgA986Ww0vtJPUy0ssGklG10yl3mn61JmZIxhx7bLOSGPADEG
SDY0LD15sABHKGZSRoouo1bqZKfhQgJPc1bzg7yBEOi9O2GuHrpUT0dunH+04Pbd
ql3UVPCx1Uyk0EiVptJI0V9N3H5IE/ksqmJQ8OMkThbkA/2nCOBr7rR37T/eH5E7
wphVKguMIvzBCibaj0Pv6VSOKthPhPT5UfIW9Zao3R++gUoqh8E0iHed7nS7JcXC
dVtmByGcOSnUzshu5X97cYQ5VrmIcykHR/Lf9l2PH2HsZMbiuScYiahLGuNk83ie
62UbWh10IJN4eo0UR4CdA9fvDfMxYuu8776KJyEbmt57bKWXpM5+YbFG21Hkd9YX
AQXwgP3YyQeFptG3bHp6ySl3DIefNdNQjNZcCSms2U3/ajh40T1KmSxlwjPxB8dM
duA+25AqUYuIibrSPRlWQtf73OGYoya4H6QVGZYxif/I2TCPOaS0JtsMTwdV2wcm
NAwSC3tfdelDs+wgKOWUQqT4msnSpRFL9UCo0+9BRRa/E3EqKAdN7JVXJWU5ADve
J1Gx18AHgYn9x23i+SmJasTYJJlGEqd0+YS+jTlUFCGPbvZ0vbeXk2LJ9QZoiHwu
+3ztPg11j3y7N2StlHS0JmHYiLY1yPIi2q/+XpeSu5x2INJYP6H+DAd7+3D9VxNx
XAlH9E3/cErCEpBYPe9oBiDll54REhYRgafNkb9iCLyv3NhTLAGiLtfJAUTV/ohF
RKuHTEEXIXQYUcA0qBUAPWBS9PQwzl5jWLVWUQpwiKQcwbuNZ18oVI6nkWJ3xUXc
c7lsZecVpOcUwtwZ8rV0IYaaupg1jNlaI9GtJruE/TmSBFEechUqvZtPK4AScaSG
UNFb9POBrFs9kLTZErKI7I/vIueNYjhBfe28h8aCa3HYUUfOe29hurfO0EjEX1LU
E607CkrrulPANIsqk92B2khfmz7I8SbFWeiqR5hiEYtztvH8PJTuNoSThg6nWj6T
q/b/bZajvkykQdxwQsDLl8xOm2LXjD5YnHfgHPDXJQ16BHAZMsvSP+mkBD0iMPtq
/ML0h6nGNH0L9XJtqGUNyMPok+p2ZoF2GOOniWBCQ4DvZgQHEvnbcaTIOrg7LDP6
M1qnb4xDoQHlQ5tlDRu+tJ8BN/Dq/sgQ5Rs5oNJGNahel2e13+afadKEhBThyYoo
d/Pf7Onm93cxw5EUjrBkjlO9QYHYEz666SOixo+wCN6+RGYinD2FrLZerzUN384W
dpWL2ahIy6S5xho9rUiWOFyS6xHzINRZ71WLdIRnOmP/nap8XB1A0mnsAdGB0T/6
JuXNi+eTd00zniHT81yV4wkDiFihO3z1MmAXsGyeUskFqJqidaU1XFaEko7qk+sq
ierr2lJf8jHNC+AO06KVb04cNvex2AH4VTMbIqJS2rLkR7BUNQVslyiFPBX7pNOs
dIVSpZoTSYy3crIRwTKzEX9liwVuVJYJmIYF8RYwbavOBF8+gCe7LUyCXGljB6Kb
V163sgJpCR1cZqr+78Ttrcd/uKqw3xtgpsQvrMca0hLQfLGRP/EAlhNnlGOEvG/M
cvojhsCNGz0Yi3zooQMgb24IclZZjWz+jyyYbb+F50LXVxtcjlZNbRfY0LU+AYxU
E1QSg+CnAJL3V8/+l7N/8mxg53szZYDrtocPKLCmY4/JR2C5bZVbfnXqxwN2C6Yf
GxSm9LyUIRDQ/IiKw6TJFGzbZBKH8G+yOVhRsw3wW5BOTdQ3oom54oBDw8XZSwtF
SMkUrhKPjqEoPlyr7/MXc5i3dLNLV2OGFQcJ2kjvP/hLrZHkFfS/h4hUEqRXGb4d
G1yXRXTFLdS3I9eJuT6JNvmy2ue9smFoWNXh3a/cXWCsaQhMA6v+lKYbi+Mi44rj
HxyAIgqW+i29N++rm2qaa59PSvw3I1TZSAhMol3hpFHILMamHSbGrrDQsRMG+cnd
XTLGypfEF+UGk2GyTaD1beCdNpRaNwgIbydpUis2KuH6w+VC6kv1Ll4l7sNF3VUW
g/p8KDFz4wR89nMwTfuyQj4dWnLf5efxqE5Qn+Jtc5xU52gXtfJgbmbCadg401zO
X0Baqa4KmLQvYUjuIJVY7jK4aOeBDp0xIrtdWSHyi63FafFMoUKXll0f0vYjqJ7C
cX0bzEE+hqog44YHYbXGJ7G9NSYcrPZaLKVPcWIFvhCCidL5nAWIcYBZP5qtIeqx
U6wjWJPuy7433nzCfv/dKwQLropVjHKyPheH4wvI3BumuKpqLjyzbh3hELlgkmen
xPS50ir9rcMOxDR51uNj9DXA+iWQBypMsjqmZlZM5vuoYpE58ecqVRtD0djxZjli
w1kSv+w1mGr0Ur+BHMBPyCQuncmF64rTkcW9MUVDgcLUGxxvYr4A1rzDhc8SyvgR
qWv/jiw7zslmEtcQZUdRaAYgiRTvnkpgFthPYTrLSXzQbx/9scG49rbr39KN1+C7
TgfjiXjud494VKYgAM8oeY6IF8NQPUV52acCCOo30sD61Sxb4Z7paAMJFpPQqmk2
+ymb49irEO8ffujIut7cw2NyrHuzhRY+ZsWurw4Rt7q2YFavKrFo8/Z1wy4iPIlF
8X1SZe0yeAvMlmmgzYQMnhDZzhxLVCf4RR5z+E0rSy2BZnl1rQSxhZeYYu+r1dsj
yH0tTFwx3GRIVIHUK6/d63TETIuGEugTy79A0ubKqgOD29fHfAZjBXVyDd6uFUrs
6AVhpv9ntNtj+0mMeo5fJIqbsezJ6IK1wlyivzcRggAGohIbmP7/tbwoXSj7D30f
1EdDSQ6k6qIL28bG+pDnDyyri8WUCeisSetm6yCDE3yND25JhKSc8oDCV1b9kb9X
NRWig8KZHLQJKLrQEBdx6MAJ6pw+30PJt8XQtnmDOrM4Z0VNHUiPp64ym/6IZt1A
NmrraHPkmRRaDm+3jBvE2swEpojMqzoTDPCE51SRqmxdub12oe9BDrddVM1V6Aua
IOeB33qnBwyhM535JbL8XqY5nqVFfQIV9Q3nBObvnyEwIg+kDXjuZv5iPFwFpfbu
J658yG80y4yGMf0AWTCDIRISgiQNDiolaSKvLwk3Hdc2aj7kR7gs/45xpk9N+56H
rJKXe0qTF2pAR0VVAPETNiGsW3OAcyeE9AtFAvPb592tlZmupLz0Hw2gkNpma5aQ
/WRlCKVyXXu8fKLRKmM41InsJ1eyGfM673Z+Oih4BJGFhIZ9G1Qk9ZqE2LJgdDz3
YsBXDdBsGHbvMVbhdExNlABXLUi/Tgtn/GykUnkkbIPjjkt+IFetsyTX2F2tmg10
Zgd4JS9UVFVrnmXjDzw7qqJ/c+o7BIeGROFvVYbw5Vkujh1BGiNc5XE7Un3BMHMf
cUx6jnIRc8oJljNYzzxdRhqVJq1S+SrFS9JLTl6qO9jNp/BHwarvL5/rQyLdVJI8
dTSNhqI4DLKbUX4gpiH7AG/0vrN/JgTwDHXvgfmiuUOLgsK3I0GOwlfS6Hv2MP4o
F75VzVRP9pckwtIFaUClSocr7d3d9FXqnoemULhEZI/tW6X/FUhEHBSPCQexI8hu
4qiNrUG3wSzO2kxhKhFmN08qh8XDrgpDoqQFa6YgAsbz161A9SzPxx6i5akvFQ0u
W05V06jWw3oqCO1g64YyA/mIpyQvDeARLrRQYfUi96kuMlJcd4NlGp6X6DPBealv
pw4j+cTv2o7sqxvh8u6flWCoPHc35YCSq81T8cDP7GHOBbOmj6SYapxMGQygiqG7
qnh38fr4aJDBE8xBmaAN0DQKaINSh/eMu77+xGuYo6RkXXXaqJoTBpx3tQjjJucS
kqlANS3tMf+nj0zUZGZ1IsccS4ichet8Bf63uA8TEEKVD9Qp/R4HPIQXf1eot24x
mRXY0stKs4Dp4xrUwZJfGAGwbxo2qvcSLZmhMuZdDd2mfDgbP98ZqNtMjUOdSKf/
yvl8GPV0j3KhIrU3TkMMKR1j1OMad5YBjySIRpEoNYDoeRHpk3r+ZiOGV8Ox6u/F
e02X6dzTKKIGQgTbkWdozKyl8tiNlq3bmipL9dTyB327P4SbnoFwvw4A/yNeZ8PE
LoeeSNURkBZ7hAGpe6Uea5thmxzBbfMeydu8yMei22/5OVlBnPR4L4uuipfhTYqV
8N/bdGPkPVUJDplyv4XFaJmrXJagaeIr6DvsTAy6vO31UeWdbGN47VCzzBl6BP9m
VjhP1Hzd14s9gBIK3TvUcH5r50WgcZ1ZEtD9HlhkRhWvuHXomTrcL1hF1uKgEUsD
6FXHwl5SPh6cRXR0Rys4aXOBmoyk0DEwPBYwsPCts7XpojemsLx99znEHdY89KaR
6AJVuzYFy/Y9yjpQb9i9LZucNZ520JkupJ1zAaPpNbRpZFm5JRU5yqZ82HAifo5L
DFoPT6D4Ehc6vk/bpOE3bqHzCggNxG7hGbOS9qjSVLHO9bXx2sPKLUiQh4IiSoAS
K9fI4wVt8TmRGoT1KpgPvagrN+3sEGv0QcDr2qoCMzbtKcw9rdURN4qM4BzDpJxE
vn28Vp5U3Ucq3npIJ7dacKz6BmnyZ7M9mjt7WN5zBqC4U+E4WCxC56OC5BFjqcds
L4Ow1K88ePtD1xzBh6bNqGNYyfwAaC8rwqCG/D9iIUSXgDGAqoz8YOsYhf9UV765
eS8/sgn0W/SVgXY6dr0Xug4gTAXZkmofKugarN/Y1PqZBdxpF8q9mJ0Ns0pdUgo6
HTykWQs1ggQv+hx7U+G6h5fIXkOsWvX3ch/ZoIdfuEsPqaJfdexiGYGqeG/PceAW
ho70HDL2m8U9aNzkp3S80v5i+2YdkoNP+xNHkLZ0Aeak1iVQ5jl9wsUW73VM89M4
jCW+OOZs34/o3n6dp75SRRu/rqDOrGEymSLTFsOFS6pnD5Ldyim9PtGUh0Rs1XtI
hzQkYWi+Dxv6aFMxyc0EISyX5YHD+LXpI6SdvOnHTDRyKPz2XhZopnceIv9/w48R
v6+JVWZ4V2RSYsT+oMu8wVqSlV86E2+J51+fbsGv1CltgSR+MfUEtdA/x5sVAfcF
LJPMWv8Zecm5H5sXpnx78416VfU+MdH8rrhcVYUIxImzcSYvsZgHF16Gk/y6Pw0w
X3gLXsqpqDyR/oOvSs7+JJ7GZS+KmweF2zgFKLseK5S1Sl8GUHw0K6r3Er35Fkyf
xQL3EayPvDnckDGdOzpooPNKIP0Acjzwzegbxf6NHge0BpWGELsil+KIxq6Polep
bPle9oA5KtrlFLj2fnMpgR/Z1UCfC49W6u2dIFCgQpJVMCamddvTUB0vfSYb4h8c
wT6N2dRHwE6rSR69wy5r9nvJWHF0EXVqjpRSn1atLTrETg347EA54qspVxMXdXon
4EYHsYVrapl2yDskaCYNz9HxyAwuoNYR1HEFdktPjeu71hv01FCfOf3HTYccilHu
r1oALSxs+ASNOz50rSMrESQT7SeZIHupGOoYRnDKRCG+/xdypkwWGqavTcfKFOJj
T/FDhskAKuuPjlCvjit9hTslnR7nySLNd5v3kDusJXFcziuOexYf7kpn2v7gcPlf
6qBEf4eywoWExKadFIr2HYPGKaP15mBcAsQxr/47bTGCZ7CDm/Ms/LtNeWHLauyf
xBDTNqMdAIMLPeqdI86Iz5VrQRSCcqg5hKHTErCITe0wqRUbrOiM4xyuX+Uvtg9y
cjrRBe9qhn9vfdyOB8kvKvvbJHEmbuOiqxAZckPAB5NzgfAq3bZd40PE6aXjedGJ
z/y9ZCwj27ZRvg8gt2uK4ZiL7YVuWGaSNtsHqJpwBOtCqKrZcMkEQ1SO31u5Ywq9
9Djapx03S+8/TNcSRTwPka0XhEqcyyB6z2JxyXvkBGHAo+lmweAip2S58DLsUqME
KGo2xe3ueuO1E6FZiothrRriU1diLhP7E4KvqSlq3QjvyYnGY5g/IGlDK27z6UKY
+5oHHXP0rtj0zxkvcKqXq4WVJq/JXHByz1qdgh0tM1z8YWAkbXQVbdLmLasSLJ4o
T05EKTQXSF9B3So4KXGcCcIuNJH8FOb1MasgVXbCcAd6v4GebZAIhf+qsphNbCLV
QOmnkxRhyFBRq/be/s6whpQahCACPlj3VTZlxgzYDDyVWFiWC4dXkZK3/xG4+hUx
gMQT7gerOOEM6Hg0lH9fanGJ92x/pHukjzh3oGTNfBc3pTQpCSL3FRq2nxvQ5nXT
r9v6HurTV6ea4o9z8lGShjIu786S53Ov5G4EPwiuY6SIbwpdCx2XlhcryfsTlj8N
9FL+OCWqiZo8l0dIf2cR1E4gRLfhe+joxYVju9Ba9AC2UvkpHr27Wt8k90T/mM3N
t8B+pCXs4OeS8DLkHW3hL2ZkL+epDjysxp6FM3Kxq0HCpwAxKBEBRn0+bHqjEGUk
GlDZJcvyyFoFmoLoIa1nj6Xx5i6wg6mQTK/0susI39qQrA3sQA7UXdHtFsv2qqCY
PYwf7Cwd2lPRAyRzuQM9NQJkg4N1z0k958LTHbxp7h2eTI4A7CAgj/hyq7ok0Dc9
SUhZxSCF9Fm2hOXj5Y5CAVfjFwgcQ2lqX8AbgBkwsIPT+LvhMbLeU+4ULWi/AqwZ
WcFsaT8bkS+rvxIOZhNrlj604OYZhe4VU86R9TXsv/wiJCld6a1xIYIepE6RosA1
Fucq+US4ts1Ih60xj+0GbhgfoUett5jQyQLboDqQfRYOTHaeNx/msctNh0puw3NR
g8uZRMJu5MbL0hQr1rgzR7fvGjv5TAlPTFtfGiaggczQnd6s13J3GbiN41yyja4H
YN9NROWt7Fp36SiclMa5XvrMGBW1D0lctDnrn47eWRbREjR6dQYgXDyP5u5HUR7A
i9SeUMCOKypLOj/FCg+/8+iuPrPDJQJxL87HU5FVfr2INTwnQkq1NL2fBXIDXgU/
NAZafXUfQ+k3X6kjLWbdyt9Kf5Xp2hgeMAU2CmQT2nZhG2Ix0L7BznenzYXt9txG
q7IOzMC9xsspn7lqwtRidCH86VudvyFbGO+SYVxmasO/KCk+9TkaQsJsGx7J96vz
khD+4AUHaB5tmZ6pB1g+ZME0X1rGD3T8NXgRQSUqRdLRI6G0zAbmZRzcs2EwN4zG
/y7J5aoikN0PXKtVEaFJ03rKq9llli38GDg7AJZ9EzgratLIaECsfVVYLRJ/knVu
tm13bAW4FFP4x/DDGjSCjOMX+9P3YhrNOVFV2+9pYeWze8q7lW+6r0DK0gr4Af8t
2Ewk03d8QFeOFpKzT0HZDXk4++jcoJWF6SB7bLpzIfR2NECJnsC9EZnhYJ92i//V
GspUzUdFMiowAK5wE8/fmw9YbW/gGiB0rLDuNtIwLdk7i3gZazgAOEachIg/JVMs
mcayP5aqIQOvGlKx75KypEtivLUlpCnVHFSLUDlgUTpxuVVHDyescNFHEvHR4PKk
Kny/OwmwcsYqsADXS2RiPu88YoCfPQOv6GeWyKpqLHZnqHrug8TfUtJucnqJol74
8khzjoUEjhmPA0adELtHh1Sog5LmawkHQF8tkExjXaKprh15UEEf4F6IkiIuYSqT
bWr7TczfRXRR0HNc0R+XfrLbH0UypdIXTI7ijrP5xvVTi19+cNKaB0WU831AHBNO
42FYWvTHSZZZAJYaZTScUzz1PIURns/BbC0pTc6vj++xCpMQ+lTvRfiqjTzLPuuV
dVV+zPpln+/qY73ehtVNFDJ4GDJyqFGdHnWJew8KEtZXTh2j2uPKbwEIfepn8eEJ
Bbb+Nmp80CjSN100P+V+RIxEJh8bCvA8eJss91KGmGg596hvVWm28iI0PHswHKQS
dRLz/1vZ7Ix1FAdWATtI+9mLd7UKUK2nqxHcjBHrOCOwMixcMJbIYqBcc+XbvMfS
cT48FM+S/kSSXEOJGC9Blcgz1Y3UaJqusIkBEzkc2BVXoP1bpez9W65FC8uj+/+b
zK1JAafhc43104tO90Wq35nV4oFMnK9VgGQPtNDUJr5bufn2svMAacgo1LwDztbW
c+3dksbjwh5Z0MhxNyX9B5BRCSjRZaEouQ8cNnFB3As87X1XZ3maQNh09qzl/Lup
RGzdSKpaaqi25LpuaeXyyA2kfEInKp50cgohdBiJuT2VL3spqR3IIb1N8cArEmZk
8mND5aWbjGsxhUNCX4zRMV/lkC0TBFT1dd7/yOMjx/u8iqypF0pzbRbxeNKGgnvb
ASXgLtAI/dpyzimVwhlBe9fACCBNaKb5s6FXXzz1IbhLRFSPXkC0RJ7/EhJx4LzL
qfye52JZn8/QboG8bi5h30QgVm/6zKSVyKgm32s8/IYow02QPYc8d7BWtprmSFfo
ur7p0+RfedLuZRaTTpJCRJvyJiBenLyjdhLr8xLO2tFnwiYLuz9cdBjp7TR+HzP4
NJdlA6ntQ6pi4HGr9e5NO6Kl9YCu8qSzC6YGdcs5Njacx3pK/pAvwiqEkON8c2/7
oILaOjRWPm1YKgwbLLG81cTeHJ9cJT5Xv+4oK73aNeXetmlq87ByGyBVUbFWLwGG
KyAR8hEvfkdZXWJLJy/2WIojM8BwN9xG4/4ZBP/r9htFZM3G6X4LcRUegFjPvUK3
ZHua24uJNorF0z+XWqN3GtQc/ou9sZHUy3vqSlcce4A7UytT+BI/Kn8goMhanCb0
RevQqj+2G02tIKYUH5UXud14lUdOlmTWNDcMHz8n5UjSZhCqwlorNkGZ+t+tQzqy
3OAYeiBk7VBM95xwyHGRnrVoAW7WkaL9IGvjTo/5wDwt2bPsbbfHU61z56luK7fm
pCwZrjbI69Gkgm1Qfldtr4W/BpXUpyiTH1gE3fmS2SzX1Gsoxsoyz20mgrtiMtGe
W97ZkSMCGx5odEK3UurIAK9LEiSvYR0+9LJ/h22LpKGlaXMGr5L1uC8P7pwXd3lJ
ReKRzDD93IJB5PhK5Pw5jZl+l0NRoBKazIVeg6l9GIe503/GKBdS9JsaC59AVP1S
yW9e08mWpRJSukS476HtZbP1s4hHKZvSN+ioVR88GvD6HORZQx6Ho6hSk1q8I3E3
8COnUP0BhVugT/BjSHhp6zcOB+TkGXPJFaU0hkc4/VSiS6NY2eSJFzdxX8a0nT5n
XM3NbiXdCF9njVLtIzqAWitMVROMYqgvohwKYhrNkWKXG3p+NELEB4OV9/w7Aci5
UhLpUG+83GMBIMN8iWY4WMPn+k8V+7GSFIJYLF4bEkd1Hs2i3//hrbazYcP6IydW
H49FUMiyTC2Kmk+5JVvwzG4Y9QSDqLUHqXo3ACQindf7xlk8bC+doBrlUJpIP1eG
suwLG7+3AU0WWjKH6bknabB6iFuuiGyzybNZNvzCW3k4jUXAtvaBA5SHuG1rj1uY
RAp8UrXfWf8IvfkiSguOeB2XUX0Y3CV2VNRIDBo6x9rZ/w5clKDEzxhHFz9WxBmg
DSh0Fcc337Qerpxy7fEamPv+QE6/a9WWyCbrLFdUy4c5u+kXq/9xhUo917SEIij/
yzV38nDEksbF6D71jccBYwePzNHY8VNPy9FhDpJKt5eHZxtG2xv3krJubqpHbWnT
fjK6HbdXDUuQl9jJLhmd90eYPKps8tmQK0jpxZ6Owd0HyNEL88H0U/bgGZRr/J8f
II+mXLVRkpFt0YkNOWIuqG3wPucBQM5pVbjlypxYLHAXCE1zKBXQP2qyLP90nUtS
SYGWUdgk6ehxSniEPznCNMEhGI8spqug7D+Oixalfu+uv5SQkXgmtrhlMkx1FpUS
GslJXjAqGQEWxTs4ZRV3upcJs5vz9GpmanGvkQ71RuSGLA1/SJ7vix0X9KyCKxar
zv/+9RF10eZhx1aFKl01fA0iWCrJfKOj2vfQ1JaqGWlwSJnTeahGbXkb1gKJfhNb
5pSehXYmWPDMOqZxpnfXeT7gseHnJgVzTra0WAHiL794qPdjw86Mixa/Jq2BmT4U
2xDD3A27i+mUT2gDuj5MvF0LbjtNAel4S7Lo3IOxxvVTw+taJ+ixZvUzQVaq5TYr
v0phyKp0SlpTvbV1g2G1FoEz/CKyYhDzFhI5ofCR5HvPqvQlX+pMI3qAr4EATJ4p
3GAOY04XuSDvQBt8KZVo64rYhZlXmqtk8T605+nvsvoGctzDHkouWs6hv3m3X+c1
vGMfUpEbfJUXDj0FIvMBjAZPR6DR0WIM9cl1tmhMAIgudo2nrZFQzIyZ+gqnZN4o
8kofBHZR3Mz9oPa6x2cWk03WrJ8k41yFNV60x0vrroOgyGPUMOOSBg4CUCF58StJ
jS6oKFpcwnZkPAamMmSjlmeXIAfLdD0f90G6D2odJSuCIOdTqNp3peWB+iVRTwBa
kQ9NiuTPTM5R/xf8HdTzD6UsRxofC704BwEVvDSbGiNjbxhRXDIHS/D/4F1/MBDv
BXvGTG/WKFop133hXBPnQrFZIMIpju5BrUlY5iEyu3seovWGF/TRPdyGCYYi3tPG
eBACYf02N2riU/P1SmP+v1rYvAO1paexRX9++PHhMhGJsfYyEXPN1tXP1ky1Duiv
mBA1xoLCwxFQ87wrNxb9438otyAgPdnjyR0P2C3S70b9/UgLLvcYKFOxt+TLaBbZ
VOcKj4sIrfiN/RMDmIMvTe/NDpNZctcXqEbdGU8bcddS8dr+jq9jjcTEwhZtLZ5M
tAaCinF56ztkTPIB6EzTz8c77tEkuGFnQMOrKxJJBakbArzU6ochr7qrpwgXqYCY
mGDEs958UFwEiMcTdHYFC7HmTjNcamQHabmK9qWkoLoWVM0Vsx6jW1QyJKlpUund
EUQuvsTqMhx01Z/k6n9x6El1tYdcaPV3tdouftst+R+d3vAOL+Iux6MqTGgUBset
laov/nbYxiXiJos6TOQapnNq+9BbxUVaWh6gX1zqS+OcWXMZG5SqwjH8OAdArij1
mW49YeX3NwEpf1HDLsiP3YjRBSEIyt7MC45t6lKi0JCsjjOKEDw8/9dVaFXQdHqO
yRs75kbzKvyggjHrvNEC3Sv3XpxNaCSXbxpPucxEBZR94CcvhtkHHla2nfRQjL3i
r0Zanp9+Q/3lSwGVsk3RvPBb0HxZqDXnyjiRITpPVw1GvQpIcDGtubMX9Yi2goD5
BDKJyv9kNmKhBGiOhuRyG+2HPeuFHr05kmBVA6iebvjQu2A124GwxGl9Wq9pWQ3K
UZU4P/MgelASrLmIgE7mZl200LqeYUDpAJNo+i1ArtvzOUyyFhCYTb1AR5AQAz3s
bkzEEH+2ih1k845Wkskq6esLKxZ4UCIHLKjCpu1FqFHnYMgoZa9yXGBIfbEzgLIB
SB1Xo0ZkV2FZptEBJsPHg4MHsF6Pum8LdkKiHPNsXD8Bpv/49chlsZBVK/vhOX+y
FGUPiKbirKv6iDVox1T8ImsrcTfq67kuHWz1uaRRTFSxRdH3QPFEfbDs1ys1wPqy
xFE8IpfXrpTRpBdw276ZCv9tWrudxNU+1W6NABmbCQ1kTRqljYRj26Z87FDen/NH
g12vrhKBSe9A/XigvpqMnuiq8Yy5g4FlXlkjujr4Ym0UaBLntMGtjXrXWIo3Rbd5
Bm2YoEjgHp3iI8+IQtVXB7zLekbpNAivZ/BtI2AsNjri9G5OIXwHMoYOnqny0nY8
aIFcPLnnIRUvbEeVCKKkWWsIi/HIIFrtNn8XzlVkT2s9QJdY9P7L3fJYaxQKa43P
GY2FtxjnCSpRk9nwXiQU3cUzpiPMFH+rptlkWWq/19IdHCfF2upJGkabLFoiDAPF
0L9XIuJB0d/2vPEwoXqgJni1XLWHRwo1dfInY9gfu7eI/Pb9z8Cv5Mr/g84qkCq8
oGcNXO82bPfNst5aFMpisQlS2nUhLCVbuyO9ggiJAcJ6E/37PL2xU/UQ9TtqpT13
qe0UxPOo4rQFrzWm8KAWWQQt4Kv0B+2J+ivYs2yggbS5EYIRvF2IqHaVDbXNmmVx
QSQo4aCj8niDnQWcdg+YM5RBEWWBM+CiEw3McYzK0qlD0j9Up5wgaJaROYcM2zJG
MCkKYiE9Y9tE/9VzPRJAePBDtxWeuaLRYxy6U51d4oE45YJmYlcFRQ35snLZ5/Xo
kxOmKUxaKVBNfHOb+N0frHRfvb3dzOW8Z62/XiPNlpf36prwNasoeq0G/zurRqCZ
xz5ZEFAjbKK3xaYdmnXKVs0QpJ3lixKzFpcj1Ji1usLgBP5zoyLa6w9h/wXD0OGW
8ZpPXFcXDrscEEp9Q9Pyi008gULyxQXpn+WzM+S/bBqgfQyq57+TJzIcdMZb3q0Z
E+Y/GgIDOBXRitGDFMhHSN5GUzUa7rNupwlmJm+W8SIc/wd1SGESiccbjTmMqy+c
AqCFyY9Q6WXvjzfDcs0kMxTkI6fB5tf0gPpJoETUWWA8lWWITHrCmuV9O6KQ/P1e
5qPmF0xt3ithZadjHjhSKlW5viATKSmAAjDFGoBCT8+pRhH1e3Ky3uNsPvDYN3H0
sIc+XA1nyystHGWVMMZSPlbHvAnWcBqXFtTM0GwzSczH5dKdP1Q1kbQn/pdp3TXg
v5WD+MHG8PTEXlK8I9h8qYqaMH2Tob5mKI6DpEdICR8cxqf8j2IQBMuJFjQek4I2
YWOKzduMjDUxzDn7lEk9Fbuhmvobs/Fk1DEOzJjqRcsuRUoWu4Jrvl6BlyyOEy/4
eFOz7bvHoJTxXEB3zq+axhyQvhtR7pNmXcYWj73bYlRS5vy6efwznCIBjQEru6EE
4/Qhc2wcipsVhfkLbhR0Se6ctayfYAQ4xOdaQdPrh94WSE6hcgx50c3kYpd8gbWn
61oEq+OWvH2eQZLGOTmV8HCx4F6VLeo3M9IZH7R1M/CdkQ9Za5WVGLrFOxqfWRdx
NjgLINRmzD5JpgKtTytR5+/sZ0hL4Duf6OST0k8W3QLG1WfOOlEnQZ0X0kUla6it
WZLcWHf4/V7nj+cZXwuRqE53IffxZCFY6JqBWwEmM7h0b8uwZvbRfN/f9iXNgKM9
jBK1xTLRaMES8AW70S/S0OdmdQ2NgGtnz7qFu8hWLv6kCqozpWmeSds9DRV5PyON
VoPtCkbgicbunhDQk+Jbwkj/Z+Xo/UnhB5Or7cFt61RVD7uGIKlCZ/KzhMOKJOkr
BpNOG26yl8MI7xahGuXPL+1Nprq4FKq32MHq/cHfVWPnDWeEQ6FYgj8rH3U0r/PM
7aqV5QU3K5RshIySGMgf/w0QLcW8i+pOBMrR0TQOoRhblfva4oHBqTD5Ynnfz+FY
lGQGb0mYJyhrLNBWjtu5m55mJH+Q0FZ8LrEyyJ6phcv8CyFxq3ypuNSQwf9lyPv6
GtpRK8A2WElabSQbfw8v6M8QmtksrBrTruHeGyxwEgiAwUwTnNjqKGWJN4qk9UL2
QyaSvmGA7kHEmYFaEZ5OWAmKM/b8fkmjVthn7yZ7qhbAu9sMSkSW0a8MnzubCCbo
96FAJyG+9xwZQuHNhVFX9Neh9VQEhh70C8pP9a1+oBZPkbYwfck9fJJ6EFhxJti2
297c1xKae+kHxwrzvtAOX3I6jeXTJTaZa0k76+CUDOAuye2nRuiYW264qFhsq+VZ
wv3vhb04z42XIeJxbMqbhvVo8ZWtqKGewWC1+HvmQPbPAsDNV29fLEMxEkfmy/Km
YaCA+o7NIDmAAhxKSwhupSc2wVd29NPjTvbGGPv3Yei1in1CZRaQWa8/NucZgWjf
ly1LrtIQRi+nDlnOx7hU7CzkklhWMj9gOn6ACFQM3H/fjCKMshNtnEEK/MIKsicA
Vql15fjZVfhqTvtgl+hv4gnoihXhBi0rFImUb+eVn73QzU70WwZYaL7Zs/kPziHf
50Iylsp636F9zXl3pvzBTNAgyl1vwKAh7/v+Y0WOgVp4Rb8b3vds5bcO7RFPk4yn
4uxfHRxYJhHkwnbJlmdgx05R1pPcMLM1H5QhbICmi9wnBiCRmHYMScR6HBm1zzv7
HG+QYyOH1/laoYgyZjbH9f6qC8ynhs+gcYM5D1jxlTd3JbBQ//XeHCTHg01Grzrz
h0gIYIKmhNVN1NFIFOo/5JUq/r71JeYDX2TkYMbqkf9Yg9/vcCTVcpNsoWWYrmOY
t7omtdf4OovOKWesdqnaova/8g3OlqwO4ZZmD8TCxsYOlp0erKSj8lUBmkAO+h1K
SbHJPM+LPC8SXRCI7N424LrPaTchy2IFeUhBxy/zUDR/qHlCRdineKI4YaNUHkkH
GDh23KvB7Lpdirtr/gXhRAgHszF04GlkSVSutved+2siVH0JHX/ef3eOS4lJtOqZ
s0RSJltS5yPigY+8SzTbUKHR1IKRs3c9dv+CtQ/YIAj6FKD51CGG3+y5CAPfRg13
t3tUAgJLpObfsO33lVYbpNWxTn1N23uGWUknq916dsfMTa1avAB6jl2ZkiKQCQhb
npFPqCJfKYfmSowJEDoGl8/0FnkasLxx04I3js4xbx7ONjzQ0w/5isYYkC3wkywa
6ZuzsBr1nWafUyWB6gQXz+9cg/EUGLtzX/bK1Q9gVor29oIy8qjQHiCz/dlj5Zwu
q3g4L95B8CZ7u9QyJZkJ/SPlr+nBqRVi25LsTfq+n9uubJeFxD0/XeJxFImUVLm1
vbYQmiQ4CeOJSVSipzhNPnyyIr3gMfJ0XQNYlNatOrVsvoQpHOYJipOEm7Uo/WK1
wWtNDqQc94OZY+s1+Tv+PG/ZxYNRsxOopRy3ML6Uyi+iN+oJnmZovjcMWUnufZdu
Cn23+wRDucc6dxniHMHcfNFsMkoK/Jdq/ITP9b63nb0nAjr62guWU/RvqgLydvmm
hARwlvEAqN27e0B9MwrKXN7qpD3GULR5rwgNxmcbF9IJsCZIcDANBRFBKcrSjt78
iIZuMJSzTrAvxZ8JvYpMhGj0TjYWT7BVrbIQsNIhJBSN82O9schWz9S0hSEREs3t
zS+Yu/mAMcF4szACynSzVS1fVnGN+kC5rhzXQTea6KKmWQbo/rm72E0yGOTa/ZSJ
Ce7NuVNhUDE7Z31g/XSdBiDOOasOUyFZkRQnEhYjmirCHb6YPO90vymYPbhjS7Jt
O+XrfPm5I83SXB7fR+LJhlkG0xOCwOJeTMZiKBK7UiPZxT5ve7fbM6yFon5rhVQD
+I9BkBorHrwJ6n7WF03h45kEqJlGHEpj9URHyAzLqy6OelxX9IDfNV52d0ZKrnDL
zemCtBwXu6KSmPW9RXC1uYezo4Q/+jv9OJ6pTP2RoCl9dayZ+w29plgIHkGifpyK
9cAuPp8msB1X6g/zHclkTz6MMv4UbWrea/WzvWlAUuaKSuDw73Z+Oo2RZam9APpu
jg35IpBNaOFttvPr6wxKKHhPZoHGjfxX/Q4NsOUf4BPHdGkq4EKV5r7vl1YR28Uz
qcHCOxsrh5zDeYx/0pWZJ0xnVRB26NZk+weQxPQuXVgR4Kh6yJtBaqr+ZJcnU+d3
Iuiwmn3a1G5ivbPXnKOuJYRyzWzaHSXHJD7zm8l9yF2R+fn4/p82/Ym9QTTg+aD1
Fy/Rnb0FuQ3Od0WDXgq7IRUz9HMEeqxhwDFI5aRJgNib+4WWbCNhQV4ifKGZYQbc
OL/04j6C/gGMk0HJMSJWchNZsHybhOHrvLZu2KkP7X1PfqhrrzUiUgZHwogW0m5U
sQ7XSUlvLGWj40RmkctaUGMlVQRlaCvGgeAIhcE6NC8L+Yv+R2tWLFcLg31T+Tb7
AQhYujeq2cKhcGGz8gD2a72itmIJRQhXRFlZoFh3MZ33AMerrTolxFZ7+u1+BvZe
n0gkPZhRASp+7KBhtWt8Tl0gBOkNpnjZvjSXhjKIIDC9iRoXc72RPpRs+3c2V+Po
Ar48/9Ldnw7X+HXcRkEA1VHx95b8febNWADpmKBzP2VWY74qDGCGypeJ8fzukEy+
sso5t4nMcMADbG+y1v/l5eJH2KP038cGbXaWAlfzEXJ4a22aULqYirMWo++5PCsy
DK6kn+vdQSvwHh1eq4hIf9pukh61qYirbbGaDduF9H+kA9tVSp28MwwttNYZicTN
Gh22SasYJG6m5qMFQHV1Hf/gbjLeMU/wy+UdbeegJpHerLcaBjyr0mMHMdD4nBJ/
JRXVldUWZUgCSoqLazH2Vr0EQvZsrATyebCNp0wtKiKNfZ9Aoe1Njlgdam0SpxhN
UtvgHj5tDthsI4H8udwTijheQt431FuxwWz8jM48B0RB3UoFcoazYkRC9Mi6WbTM
GyAZlH1DRjq7HC6HvzEt3yfbQ7lAJ0ywlNGDi2h5EuIIhsH3ODyPXUbJ/TChjfGD
hg1+T/SVDXDzvIZ8CzWhV2vMueHJRQKuF85LPHLijszp01r00EZn41Jb/+Monok3
jf68/Zm7QXhXvSq9SPUHil1JWrwSdrUY47Ec4GwVeyzFi3p3Qo5ajLPTTOyVXhbs
t+dPm7Q5LsvoHppFd1tPkwIKw7QZn+Ca1ee4VLAkOnjh+mdylQWkUkSYSJaEGBmj
X87ENN1Avz7X8BzT666IwPyWKwtm4eBIT1J5/HLb3miiXET14xQJZy8Kjs20e5DG
s2rv124Gjg5vBU3FKvPnfCMy3Elc775RMbwpN+iUXLEek+7tLxMEwD8t0idweFAy
Q0z91HJn0IUUD1MMx3lGFTnuszhv2S6zJHhfi/JX+VnmA5Qq0gv+0IHZeKxT0LnW
dW7LL+z/yoaUEQSoG7/WfG3zZtzHy49GSuHi4/sYJpiwZUemjbh4JY1tmfa3AflS
L0X9rPVBEXdo8LBZRQ11xZWih3W+fyhD2dT24tB9Tj1Dj7xfPU7i5bU3+LSrk0en
N0gljVwuFnV9XMeMFaEMGyzIgSP0zs1mE9FUShnLiyC1z/X+9QI91UjFCEvIY/kQ
1lwix9JZ9wSfaYl55hN9T99TppBEM9Gz//roAK3H0NE/KjngYXrQRib6+WDZWbZR
rD7ah0wXNluHHi+FSOeSso5PTuBijIx9zrNjsXPYuwRf+wKFysggmiE5Fi5KW2qc
FiVHy8FCKNXcuu50ly1+DhESbHdtav51FLibkB+YJWMVwNbJR+vtJ5kc27HdYHkt
DXS0b+DQNR9cPiuioSw5vtpU+LjE5Y/uV/57K13wqbTD42OMAEh0RaMVXXU/zay0
YGr96UGePJpmcYBFrm1J/FLryKcPETG2LjhVXZWu7qPGuKsuk/bypgYDrfTvajq3
AO17tAfnmK4RltIba7sSeHUn3YqjC4ImKTu4w1gWhf2WsS62Uto1N9kt/a2hOYpj
CBdcdPGVEtJwRksFs2H8RudHaUjyUnRD9Fqnc0U4620iCJF8mvubOX8SNFSitbYo
IxpFM3Co8Z6k0F4GR61es0iK6vlSBQYgl1BYi05xOaHobcEuPPuCJpKluaZcr+cw
7qdAjhO6yd3ctuU5w5L/GFq6xhCHFBheq1//INTzIprv0xzRko2wvGRBxJuw2Qo4
ZfrOkK6HqiNmhYtFT0hcwQVNYjfC2Ad30sIpqdIYxzn3AgDkq+IiZERSEqE7O0wU
IHpiGyHpNANNFxeYXs0zNvkW2Wh3u9jdFFZo5qdYQG16aNVTk9wpz31eJTAUJYKR
lE0Kqe19zIM8cHD0jwVCgE6oMQTj9+obgY1gaTFbLCr3WfsSlamV8aGG+W2YB0Vv
0ePSSbSEaQpDTyicPN/RUZsQ75BjxxKVXWl+z5cWdwDHD5mNB78Fm49z6rKnZqBB
EsRgzGPr8NtBV7tg6vmdcdywPxI5B4eZ2wqao5IQ38FjF7tOH0MTjAzjynqK4Vxp
Iyc7/rNCOr33RmqNg75cTWVewVKdJI3ljSWc2r7QIrkNl49Fy2uejml0euPMj3T2
tdxzCLhxlfzh5cOAHIuVZGS76bZ13Rik2L8o/b65Nj2qveNbUzhXhBVWnB46x4ur
00KaRZoGHgohD+pWXArXYDihlxRbo4PDNPm2ckwUweV5QtmVKjqcfDfAJQkUQ6Gz
pItzALT0uJEtomAC9Ffawr/uRoII6CXUhWWXXP5e+fwQ5IkS7CUC2QG5MLRNJwsY
fbiqo8iLQzGdZufMpZ/Uu/O1l31fv2ZNP4tWL7JnkSpGOTIEN1l1oXSLZQUM2/hL
Ktg+FVuAIEoJOdhw9/U9XstPFJi6qoCH4xlZnzdzCCwzSiU2Xo9KUv9hPUzallEn
o9dvyGV1bK59ZHaO75C0ksy7id0uJRvR4u5okj/gC+m6JqgRI27xgCKXO8GDgMsA
OGEPV0qxejIPLomIt9ftAdPHS8M67s3n50slpT5K0xlLsN8n1FBJsAu9F+bEZJlu
ViY0dfgxwnU+6GORcCWica+8C5L3UvBPILDDaMjsMuwjiySrcTzz4A2UK4ui6eFt
2uBXanetcK6DSjEXWuo7JZIjlegi1mIYxmYi2gAFrxkuPd2JXicM6g8hmfU8YOVr
ZWM93+fLYmF2mbQMiHXbIhaJ4sm2047goC2Zeyt3YQSNEJatuwjyMxCTr69s5UuW
xjCrGpps5ClXs+sFLOgpU1LkM0otDwBcOHKb2N2DwuUlOmX6DORFineCpWZuVnXo
hvdHsGtXZF0iese+qwmwKvRKx4verE860+1p2Ee4cTTSiyn/pD3ImJTFpSVp7SSm
9NJuOPPgV8oUxLQRC9w2asJWaLML0IhYdPNp2zQr0/wxhFsb08ZxgOUaizmv14Hc
QJfBOrlmVOp2diFnqiw8+XGrvE+bJFo03U1VnvLEhNJ5+n4zNL3NNJS+qnC7jHX5
w+U6VZY2fvug5L3De2L/RHaoForfks7NZq/J/2rMzer7/LNCN5LO+Z6xe3q+nw/J
6bSTD13Z99yFaeGn/idW/pHimI8j0qAJFSYfSNebOlwl7WZH3mV6Bqmh+CPEsbMH
idL2eH7wFbaswBhSqMvjsV5mKVuS/qgt3CPwwBb3Vfqvjt1fVmjwYuU/egJ8Awx0
p3ZmcGHqlqr1p9eEUUi4Mj30abDEeeuleC1iFixDGRVvO7Uu+hT7o0ZWeD80WMP0
u1PnQmKjhs+FwwZUVW0wKz05u4EH2x0t49tUsAWPkH6h300sSIrxntoHn6/JSnXF
rea+gAmr5r8USzYrwPFnqQWJrduaFbggid8nce7ZAhHJWBSdCGNQlhTMtJkKYOsF
ryIRmgtzMTQdHwQHf0J4cDT2xfHh3Baaszs0MHqgvfovIHv4o8WPwm0rN56KKKDW
6gJfp9HB0zM+s5AApOxpHZdVaANc+31n1g6VHaI4Z9Ntr0+6inhRLvU2VcDnlLe0
PGEGzchmkWwX3VTEiKY6OPcHTr94FlCF8WRvCuv57bGY5HqwE1QM0sNqhmTwKh/0
9Ervt/zX0Zo6BH8euXfgMiSpxFEUr3u+KM2X1PSYTKxkjVghNBpUlDdS8jcauOJS
IvZRQz3NbtENfSj5X5ZSuf2GjNgYJBzuaZufC6vHoWjWlWsPVJqA2qu1OYWpX2P5
6TzKb0K2YX0jBb/9P4WKHQag/Dq6/3bMxCScCG99N+9EyGOSuZiNofbNNsa4SxFo
xQHI5ONHp+4/aqump+Cqb43GWtjTLLbhYvwJumE6VwyucV2d1jUXXyNyMV9vT9oX
TtdDegiEzmkWyMboNeBZa63jtQIlyJ5eoR699v9aCO+IrxAIQ95RSiUfX3e7HBXJ
M/M81jH/t+2m44S4lapB52gTNSxnEQpGvzs5qJs4ZryFv4Am6tz7l1YRawAhT04P
GKRV6hR4bwWQbrOG9aq8RpiWilTdVIUuK8R/acjPFByugcfkCgoVo2JOYsF45n/z
27wqJvQljkb0Fn5EzrhhGWth/5XrmkalDvvf6sPvPxLC5uj7YaEEETxO6S+3UqKD
zPa1XNQTT/xscOgWnBii9HrMSqVvYHR8ismPALJUQdmqBt+FK5yMxba0W6TpDZ8y
YJvUcXQLiphMWuPDdYuA64dax84UgBpPezjcqfOkejWQNSIPUSXatfFs6sUy/ayE
PePczlxLyPztdZwLwIrTx6fNggc66KOP1hFU3qLzcPxURPovDhzqE2qvKuBH1MQm
MGAWjCcEqfLdAAbIzhPaxDKruyKThSMrhZqmGz5ejZPmiiXu83lqkWjYyoIKZLU0
JmAjnKzknd6/x6/EH6yEqhpcc13PkSL7dt8U+9wYeC9tjxOOiLcC9XOx+H1kPee3
Y2HpR7iRoivoD305WAF9/U8PhCKdtp1yUJUEXBgP29+RxEbk7zwM8NhlLdCLRVUw
yUZTHmB8fmD9R3ZSyXHMb95Ph0GTGETuQFs2qOtOIdIHGdHD7qhol8LTcqkTywzv
eRSGNeYJ2GwL3jHKxUZRIJZ02W7lWJu6zBefDRs3OGlZnojtAG4V7jhWQQCgPeKe
CpxlwpnTW36wvrxbi4/65aKloU4acokdGCajZ4SNuMMSwgb29fNrCMxHrpbtyFTf
+NeXYofISbV6m+fkTptZ144g7XVoIb72mFUUjSeh+lWKxBze5YpWWJTS3IzQTZel
Z01ofU8m9G7KzrWYMZpzse/fMDdVQsDKIbvPD69Wfhu1ASUTaae3cBuGSYTzHfC1
HE80qQ34fr2eM6gcBX0qWrf4626675F+sUafWWsflQhQvCndMMCLlF6BpbDlHjEt
0IIGcgedt25k5VPAcJ0NgA6ChIWuDh/vDblnuZXG31y0Au55oQQg/qpIT2dpsAVY
a5gSvt33+HaguqcJ7oLyu4b/pE9SFnO/QBw26bD1K/mGuYa2Qg4iDPNqf8iUqB/J
YaoLBP1md8klMl/P8tsEx5S78MGPrp5rAeq48YnC0bty5qfC2HLN6FGUVGQsQOXA
CsnTUujK9HktZv9Vy6JzVSCwEAlBeLAYG/DB2lhNtUf6eJBqFjSNxvy/OwcHEbol
3h0tS6nLoLmUAown83jmMwGArP7Ldnw7inv2S+XeCeJTFIUSCaD05BIPg/Jshfco
ubVoBKS0P409vCTuZgCMdFwag3wILAs/+CG6IrUCUdCG16/uMoI7fWGvcUTMwe5g
ApGOS7PEYFfdtz8MOc4oHMwna0P79cQU9E5LcFQIa7GZlis1eT0CFDD3RVZoztap
1lCAyD2h9isA8CuoJRiKfAHluV12W2jYsa/Bc3rhsx02AhfoD/LbgapfWiTJFMp+
IueCxyqydZpMzT7cLATiBkLco92WGT/9ow4RTLIMWlifNBY3WV1WhtLDZ+QtLxT9
tgGrlL6w1PJMhvJ2GMQim7Vofa1zcQ658FvXOqxSwEOQNTmihlc53JfcJAJLxH7G
Gas5Ab13CPYR9BRw5mM75Au/yyO2RMj8PzZQnW1wwHMyG8TyeEtjBAWM73zSFSmA
QaMGGXj9mBLMyODBgUQNJacmG9PC5PNkDI98BvsMpJ5OocJFXXGMwEkZpAUH/EV9
VbmT49KaBVR4A3TtRPYFIzNUbk5nXsJoTDFkzin1E+ICyxz238m/DL6JbwEyeLwI
fIVpBvtB7ovZxxAHdg724tOZMXfRHRo2Fx2bhC3YrECVQUCzDPFpULSSMfbdeJ5P
Jg65H7NTGbcbP7bngpSnGhcCqkuz8TS/ZLq+5ANlU5iuxUFzPwMV9eYhqp6kJpg4
11V/f5c3KPdvxmRiJcG94EAiDn7R0arZIcJFZD7F8GIcT2T53wOlvGkGao9slMKJ
B2S97kkpiFqzbNMfHvefuLsBpNiaHFJ9DUTdi1XvGNv63EKepMt28upCu5/1Ahln
W9Z/T8IPNLT05sKWugZD5HcPoXTnH8QXvUNdZ/wirLIYpKVAvvEt5k9Af9G+/a4A
1gw61Lw6IuHnxMkxa62LnKlf8uoHHWlYmMeganQaMHA89CBSsj5UlcW+EAZbBRmK
a9js9kA/3GJp6rht6oL+mktQ6RqA6xHWDGWRdgouE4f07GNfdSZg66GF+FJPj9+G
mhCHFhcFSHG/SvS73B415zOLM6cWBXgixW2lv1Y8FmuXJu45RwxjurAcTt6MM8Rn
H0kjk/y2n2l9Ll8sFISK81DkEhHMnwKQ4IIhuN6ytjcyjCl3QvASCgg4woNz0k8R
lcpSoZ6euqLv4GsR6OfD5WeT622Vkg0iimvqAr9b2oaByNvDhqUJlFUNCc08vw0o
nTeEs/ezEUoxt+G2JvefzyxMbhUG6RlgDH7pAm2y2JbsirN5mm9bU/Amb5f039SZ
OElBs73pSuPagjz8xdUXUKUQAGsa15qb6bCS677Rh6JZAjJYUe/HxrE2Th8PiMvU
7+oZZr0Uo5/OrL3nPQfTSGGximh9JpXBJvp6QwrH3QRPWFO5XfgkAU4R1Bx+PtRc
Xu0nnwgsViBv8v9vPtV5Nu7lyK7LMOQa+AIhviThQuAIfdmcdoW7LulVRE2HSiuN
f0kU7aohBWP5x3GjOEZOJbEOhFIe8L5MuGakecZWRDs9LmAdcDSr++qZ/GdFoN3a
9Du50+aQVFcxJrYQksakw1mpr0Q5qbcJ9jTbM27P7ZdKWFAuky4aWu0HdaNS4mJU
Dpt9dZnOZwB2AjBHn10TCLIuhyeJjhrF5GfHo3cvdV6BVV5sRv8uAfCPa9F4DEm0
2YiiMauOfZ4qx84ThBCsf70SNtPpqCSkw1fEahKw/w1zU1xKJ00x4QNXjG6m9cS8
va2cYfex4tgmG3+AQKcp52UEUJye2qvktufhCl1A3oNs/+6+2aNERkEi/UTHpGRT
9Q540c/fqd9zrGzrxNuqMaYdk64nHQTiMf0KiS3iGAK/k51r6e9kfHsQE1M69OBY
a0ElfIs5wW6QFTyFeG73gcufMD7GiSPat1stjzjDb17t+i+WbKjzbKBuexJjvinV
bK7ID3RMjwAn0ikIctXWw1PDqffcEeHlV+6mywEey9YlP2qqxhiRwQUJP0x1M6CF
o2XfnmsoAi4MWvuTM9xUfs4MmqNEWg6IuG4TK7xEZzbxMXBXxDBfwjFJ5IXf2zHD
0hw31BUIzqAq3cG5OtAuelg3b6dGHPCaxkv2GP/FS/asM4KLUpE+Pz95CkimROd7
F/sMidE6zv++6sRv2DQoopq+2x0+7GtXKzJq04woT4h4VyGzhuEtegXIChUfdQz5
W6IYbrysKuogxbQFIkywEUufjjF7M7qu9bXdj7tKYpTBo5BEEupNpDnPZQVIAg/6
SAEgppA8tMhwgkideNNTZvQE+5jn4xDOzeS2cwgJ5EUKS5aa2N5a63HsGBTWB7HQ
mWDgZfF5RpadZw2IIUWEQfg8ThanTU9XFxdVBst+/yA4s4LfiLc7A/bq0Mg4T7tD
yZfdewX3Va4+zUdJNFBonQDGqWv10XbpQpHb0lDhgKlMjG9ZriZaaWZrGztIaWDn
oMGtNuNIF0NDJavTPfm16dNsc6i4ydDq4jmSE577BGTjHy+AgoXfriM22kPMWh4d
BUW7dAibkTiDlmsH4JpCS8+/bB0qldtf23lOPqABKPn+mQ0m2OAIApv206PmSbtC
UbKBPS7dkxdQWqmba4d+D25D7AGO03k4yNFFPtZLZDNqVWatzLoEwAmHlpMDBn3g
P/+sd7rvKli2HX6oN4sB0/UH2j2xycuiHdt/3IvsxO79QF2p3pavojZGMX0LRWln
WDRitz9yP+pRYhefK8e/f+LrwgbBtPP61KvI4dJJV8wfK8grZd0UaZFwcOhJfUrK
XTFGiNRYAY/4ySv6paN3NAE14ZFsNMeeYRB8uBTTK4MaS1iTYXiLoUVjD/EvYgUG
yxK7WPNEG/nQZSBZnqtEbwUb3xId6S/KLlmaCcyL7DVeIq9iQQv8zsa1uhv2nhX0
YTv+2XSwGj4tQT9KPUlGmpZhN4fbKgUiKISOx/GDDEkrghtum8rsvqoncjtyGhtg
nDW5UQDgIwpZ6UYMsB9RueXtjRpuSapex8ist+3P/2sG4dB6Ev8R0fETvIJyCoT7
6AF+WiOZ1J+/XiwNmGm7uadTKe4afRv9PPY6qIQ3LfqYUr0iQ7ERfbca11LhsZkQ
g2djp4OLW7mblDgVRgWFDOvg73rvepSrx3+FMi8vN6ko5RZyFoXH69jcag6fa2I2
EBhJdBBVEqgNvqssY5X00te4Hb+t3+9iamJI3c5mkwVc2A/3nu0o99RuIP1uPGje
Gi7pgyJUe/NqnjvQHOXjhJbGC3RJ0bxhNvSeft0sCZGcyNDB6cX6uMRLhMHJ3OKW
y1w+jjD6yfYJtIRgD5HmD14ZYZ9n5rJCJm1Sxxg//oylesBptdPlPJSv/wZ0hNu5
Mg9dLmYnC4mUPFR5JVNTRbWRkOKOs2i/XRUeQZl2JAPXtDjCCX+ZC9tqHoE6Ws5u
EcimChMUud2B0TRA/OMlnjjQvjKdJhcAZBpyxPRbrUDAOGF4fBlzpL868PqNfj3E
dL6azz/UbNjfQ/8Ad6TVUHploXlo8PPn1I4dI6V4Ziqtd4qUzU8lF9iLRREUz0Vn
qqXDMXb5Oh3RjhiSGnJEO0sft2EC+9VyFWPSV1Kt0/5URABFSmb9xZ2f+V8lUt/j
c0jpkQNux+IxGOWWAJcYF5Tc6/XDrqvM8nol7TTcOmk9jA++dWmc+GUWIxwEOTBb
qJJV4WAYY+3v1swhzZphFGZKL6ywomoe+ntUbQU5mVl0IGVwm0XiY+yVEE3NZ6QX
T24y+21XUnDCkeVVTJTmDfhBa3ldhxsJBEqwUIGCQ8e2g362ntjxy2068mCFwTKm
A3jM1M35kTSrc1lLhMEd+dEbqI8mt4i5+Ip2gkH+RdDDBmUzqXykaUf8beeJH9sT
f76m+I8yFFDCq5dnDacCWTS4zxrfbTCbaK2dp3MICgRN3uk6NvRA5E54/mNtWF7X
yUByHtkfhf4OSpWlmJVyTOLWwYJOu5NaJsW6QBPNIuhxvFq9sb5EfY1StUZ1QUOh
mpHj4OikeFPLQqGRPjAD/eXD5PYRWiws1n5FTZwhjB7s9Bz13EG9ZMREW4YjZafT
be1mQ0sjSoO2VcrlBeqscJbIh2RGWlWCSPDfpfOvnGedeSgtQFewUnfPMRAuZylQ
UXBeOpV9hUIOTasBOLiNxnwgrMYTuXcogrGVMS+YtI9vJV03lZXyDd4H1HNTsK7f
scSkL7f9QjpLXOvwySKPE9KZL+K5FxsstE97RIQJoshNX6Pk1t+Ar0RNg0uKp2tA
CY6R28uk1ONLUn40IFVhNgcLqRwyqHGlAlgiroL05s5aFNJ7NYgZFeQhRkr3GYwh
sUszh3Tf77VxisvByD5HANLE4lBqCLTXfSTv4yq6ypnC5I9R3WjZxIQIoiEiUKTs
ZKNuLIZxblgUKKy4x5/jNydZmZb3/56b/+9p3E+N2wdQj/T+KmclisBNAd6pRJ3n
8bNVPBVZH2yA7tjDLj0mjnGmsy5LDB+BWOowYWGhDzkzJtWpHd2AGXw1GuAtbT+J
c23FXOE68oeGwNUkDoKow5N2ZJeU1pRn81abm34gqLqLTwu64VaIFoD+lUc/50lB
Q9vF95qUx/nhop7VF3MvHQhsINnTqR9/iXDEPgDHrgWbgZzixJqneuybMV1J1sWx
tPBjKYeP1Hj/EpvrqCPHjQ4C3SAEXo3UsSLnyN0RlGzn7mQtz+RExsY4inxeYKtr
NtYldudcY88iYJ5GfZaavyd1CVw9T/nlcVGdNto/nCnPMClUcoJlsX8ofLHGYPTe
H6+pwjrLrMmveikLO8NlwtFTJXS26g46h6yLRq0d8MlAYNDV+dUdXiNAQYeFiUe9
cW8btFYfHijo3xvFE4zzd/Uy6HKxFsaUnSpAwESiwR4q1uWTNeEgzMfA8c8lbeCs
HbRgWtcPaid61dQY8hKYCUGu6Qi4pfTh0DwCc2pPewtbMkvDTiBpGYYRK6aaQFIL
qOJtsBKGmCIgdUYR9M3v5zor2dZDdG94UyFdkILWwXd1isXvT3HUScbLhwB975bA
5OaP1gyGNpW9KJRSQHynZ1jfnPaJrMFmd9AGBZ6ZuYrBO2wF5iI59uzHyVYgOtFj
8/SR6Rh9xRxlSriQZsK29y7Kj0HgcSyM8l6MVkToCDe/ee9849SwuSPCwspnDp4r
ti5BgllAIBwJAL6E9dwJKHe5w9DEb/DooMyghtzJFyHhFDiz6/wTRyGJh9d0fpAM
QZnAcocKK6SD1SjbiCPDMLCPiOBw3/vFKPRyb2SLJJZrbmabDAmJuCA57CLd0FlB
tBUwk9gkm9atS5gF9AJHEOrF8LSN7WKnaYelVLscqc0oInTs4XYtrj49g7nb89Ur
KbF4jZ9ptP3feyKNpGRQdx+IW+Tf4SONSGICu4cJzQ0egPxHo0PgkvvFGHzBKOef
i/2a0VQxP2t8WfC3ndgIxda3KBhjXyLJOM5Qx3fXQ9npVrlRcprZG01mgozC8Ffn
7kLrWaS48KwMG11RxdTxn+e3rFA+0bikuXC2srZnsJj6BND4uW+5lFOvMmMY2C6R
kqGF2BN7u3AKKFMaeI04cP8IeIt9VjpJpTL3/dWrQ191xPD5P6hKhJJ5zbBEoW37
X/rzGFofqRiHolPQGBKdUSjUsh9uL5di4gC5KCLo2wOHQeynjsBBu9iMgfat4dGm
VCqDJ2ITtlDS/vS3lJDCfKCY2hRBZYItsWGAeRo9fcExyt8lsljnIiV2CSwE+uoa
i0kVRIPsxySM0hJvWuF5+7vVo9ri953y7c3SdGiRcH65V7lY8Z02UY/FPBws2SYw
BheZ5WwLMtkee29q4wmNYaN+Py/NjcD5DTEh2Yaq22k5n9ekIdI9RbDXbMpuoeTg
jdHSBolVYcLyvnMdgfvjqE6eiURwvAkbyuENR9TIwvMm/g5ieenl1wjsMURuGJIl
3Py8/04sjOUBOIBEsmOUVPZvM1zVZA5arpF3A1Nb7va2VUfFnDxQvPcF3fJ1uAlv
KMi/8sDnJpPr2whG6/ujiCJZGnopBR9xtO+MH6Xg+YBgqPsg+/17JZ1741WICyUz
EI3a7owubzhkyW4iN+vohzPbwxRo3x/BvBI9ndpdvHJR4IChJ9zWu0sHZonzcJzT
vm8kA5NzgVmwzXoIZmpA60CcNSOxvsO04hWnBXsH+GpAAw7QYJsmQEsn/gtGZ9Av
R8Xad/4ml9QlF2UndgCrs8XEjbVEABIHfiijA+imgLF/la2ax/u18JEchX9OQN81
Lx2uLKi22MPsy9R5C/HP/gzju15EwAQT5vgV/zfKA3oW0k4lu0IG6Ns2DbAXg9eL
p6qMwxoOrpG0vuT2kMfaev3A8/oKC3pfIjwbbliVp4eetTD/APvMVnPGN5VbF9FP
dBwJWbMavAPIYBOQ02dDl1KLgki3bLQJNMieBMsbq1a8wMQAaNM5CAI3qyx+m50E
YKcMXrIkINUvX4yYbkUaFWBob8b1c2VnQLImsIHLuiv6lBcdbChyXVWdNnfNIDcX
wmujJH0VheBq4/i5UeRr8qt/zI97oX+mu1NMRLS2J45gYmeO27fPHUEHWUZMpWTA
y60u5LUIjn9hO3N78w6ycVjabXeiarc9DZXllcvsXZIlQ6UHNAWe1Gy2369PRqbU
buCs+i7DqL7J5FPDEka2UGyVcsK/I1F9dJXkLWCbZx3zuGCJP7T7QyF+VWb6au9s
dgN2Sx6lOxDgcnslJhCNTtAHQloF1IOXCAUOkeJYHrEApwcl8E9Q6tIeGxG956rC
4iYRNEdtw3KilMvHvO9r1Fw2Z5XGpGOyRjltcvyZfTjG4HuvV/8JnK7/3s2r/toE
3kNDK8Kjt7k/crwMTLYm2RB7FaJT2jfz+mFGOT4mITsw+p+/oqudUQQ/Qjy+/hr1
C0G3Y+6cOiYHtkAUMa9uXc3i5p0XsUZBz2PmJSdajHUnb9c9A8EOFeC5InSezUZs
T76mUqD0ubkOSUscVjUzNzxW+oDMhvACoQPfd/izIlPXO6XXgGqKVluc2RGs/yeZ
LXUfufTENaP1mstw2gu0vVOmVPddk1nPo069yVakpeol1i0qCXK0k+t5ONkT/7zl
ZQ+rlIMvz9JumqN249Ibq4UJkLaNleQnbmavbgp4doEPm0Yk35913TP7WPOwgG9P
mJVfbBGeTAEg6Rb/cUtgRxcWzGHxyzREb31fbHmV5gzMLG3LXxfhtOI1PZ91gtc/
ZTNzMnVuPnjww9k3Z7ynbunsqJ0+WgC9D5H8qmUXv4dIneeuvt5O9ko8PBqF3dDN
Vcx+2lIOWup35fM59/SQCrMZRr3Bu2jCt9wbujktO70hmjjCtOeAoN88DmKa+qAp
xhA/gbtogh3abuFFHWMoSX+jF0RGwVJACCtE+SjHs3jq1FcgcG+O/Omw21lOt4y0
C5wX3tILaUq1xAUyYqP5sTE8HX7sM3NHFrBe8r+Qs/0XqCZSreveHEm3jJV6FKEb
Z+YH53VLfkPqrNk2+qSmkC/Si74BaMWjSc32KLZr5QyAhoGOURO4TWhAE+fVvciH
qX+neqkOqfjVvs10vu72Hi+tPVQcIE9tgtxAy3qs1DgNmr5wGX8Eti+iIkfKVjd9
rzr+rIc0YPC57ZNRCOfeiSdnhVJqQMSlwljzBut00h4l4A72txMbWBsIIKR/0XGa
fygxBpoytIkpitB7VR20NyQz0Yf1oyQJJzin1uumSRjycNv1oGKe35XFTjTPwSOO
eYUg7KbQU11/8f9o9o7YFAPBlUnNxPUOcldwjHwLvBbqYPAFtiJ7ylENBghcQQuC
Zihws4Orq+eWeCW8rG6fnIWEeWnQ4Uca/A33ho+CtNTuG35A+ekFqaeK6H+H8Gdz
S3K2trV10Z8L+Org2CkhMjriwrq9f1m6UH7HzvOkEGuclvF/hZiSoOCRzBhQtbXX
2ituW/2Q8hg6XZyWK/tzApG2P1YAdSuDmonxDUCAH/pGhaSJvRroHI/1e0rk4koS
h5bj9pihrXrusNy/UvJ8Tvd0vSJnh5qFwb819ghbJbHqH51/iqE2cm3eKjMirOdi
l2Ib4zKwDzPnIkaRX9lPKzvNxyNnPApiJ4Z8gFweKHa/QyFAv91JkrMm2klNCje8
EBj0dGc/Wbp535iRaLxUb5IhWYOyyH4Wbr+g4FOsHsw5SyHr06vGeCWT/co6JMqK
Wjtm4dxR9Z1GdoWsb2i26c5fXBO4T4/4lYZKNwVu1ESl/gNdPFFb777g0gjjaxHR
XOv0Rtg21hasNtd6ZxqKLLHqbDxPPzpOeQbq6ExjrGTakQKLtZl7eEqS8MNBllSC
noUjXNVhSbOvmPtNTS+JFU+KqI5/HoEWkmkioPwCOQwvMmMjhCJh0t8mvzvLpMc0
N/1XX6rM8fEDj53hr5R1dIbpIiCFTy9O7+3Mb3rHlpH2BrfCxIF47cvbX30u6dRF
sPAirWhEnMq0ITvK/EBNXbQFLOWwd09xtcshx1kInsetRrS7jVEUcsHS6ABNgdBk
mPvGbF9n3VUF9xtt3Bhe8Q+Ui2bSBmKVnxYiDBX3J/yzi26BpfaVODQvjDW1yI4l
9dvhsa/mB4zAdxavgYMoDduVL8C6XtHw5HAFyNRWEKPiKsm/gOTY8xQxlja8bmU9
3DKoCluTaQ8acU+nmeyIyOufDg9XgHaUP5bcyBll6vHM7Ne6dVJAbWEXYihjTfSD
/DkKQxusQKEjGWdSGKjNIP0sKRir6zmvf8ZweHrr823ZT1rXckxs4KxV5JElJCww
NSdBIbz2aaigbo0pM1y0jYY3SGCH06idU4Tmij1R8ozE4r2gouAoe1IakrupMi9+
RJZp5tVlHLzPhtLLVkyLGAVneQasZeGMhpxTd+ObpOsTpgmfLl8bFKaB+bxJfy2L
PqFf9kHSspXeD9K4lqAY9e4Y7oqRJtWTjS02iacuXdYi8fFbf2vgmtHi9oeapMyh
oTjy1ZXhD4igKWhfMDUQq0wT0oHenSjUoFvN85Bb7CAgEZlFGkO19WEv538+ysly
tW+OFGdEaTuDIs1WX7s6k1ErgDU5lNfgMSr9fnYCdhfv1jUJZH1WWziTAE6B0btM
SkD7EpznBAsPWqJq768Q52gTiQyI6PfmKfH35VbuXy8PsAX0cJpoU9+KfKhbWyWo
m6Bzr5D+o/tUOBcElq1eO8UFMVsFx0Jb9G/S8GfoVgw+dChsr0UBrbsXcoRmVyvm
2k/JWx3jN5CrUJHPBbp96lm5KyEbn+4Ge0XD9fDS9mWDDzGjnltp2wkZ1jJWxhDg
KVy5b0LG8l6ga1khOagFi3kmOweYEJ5/EIANg3BOGc2dZxaqcNHYBlYKCev3qMz3
c8VVtnmENsoSTSmovNdF7Bbtu0/vLZ1jmuF7yRDqJJY3LWTx59psQ4Vf/ePTSOpw
NjYec0Tyf64fDARNE5zk7NVq0IAWaZIUf75haag9JxAuoZSb9iXCPeuYpjvpBb5j
h+LA4F2t1dzhwrJjlSMAjFmhF11iPfDxkyw5l6Fai2wVpuShcQYf7/JqE6FBMsug
NRdE819A5AxQxNwem0HfqHef0EC2EhyFRSpdtpwnlBiSGJmOYHG1VbseizFzGvU9
UGCrVfnke0R5hgWxhrOJVjMjVuuoKK7f0W6t8xPC3jFfPyql1hNFkyYalE+GXzwh
4xQ4mjvWksCf+I7MhShesseis81c0w/u2VNd1GS/CQVThE3fs0przx62c/JQzwmB
P69Apa3jWNUDgOY2b2SM+s//GogaYLPKwLTdsx2C8XlevXZwl9GBraL8QlYo86r5
JgdPvRjW8LiTu0M/NbVrs0ge2IwVFV7UCQAQBRUJ7isiskBiB4lDITigQ0y+Udfp
rztfRJL1MHp+zR4pvy96r/atUlb4gn6GVpKUbjz3/lBMhsHBdH/iYIquzbmKmGLv
63cqv9gtxCtENDApkjEhh4zOn3aGmRTRfYdFKUQZZ4ci3A+URhSgZD7975PF8BZL
AX5CtwtVGtUJtml4UoAuHub7N44MvjsNubHJSwCcDIuQ6ENHaxFf44CKkP12iIN5
xIcI9PIIv5xLjKKu5BzfRryOMvD+oDQgBc7h3ZpTmIIxOYXLxOSGWoP1yfjO3c9F
Rcphljo1wSXM+54SMpF5nd7hbTA/4b2JPNqiWoESP7HrEe8L6M7HntU/mlA/AcHs
YcxXp7s5NIWBKkjPg34CHMSCvkaCM2ZR1UkdLNqpUFOEVIwyZOxfkr8jEId4lya3
zWBJ+hyaQXPp4lOdIOwYmKx3dVEJAsuwpYoOtS+G8zivgoH6h0QGbTWLwDtap8IU
N8HiyRx+gQCWUSGMTetCXvdU3FKff58nhJnKlbbxZnZL+2tAPm9lEH3MJZnlGrIA
4d49kioelAtv5KklrAv3LgTwcqfy8oZNFSVoNjeRUOwauKtvt+krfwKj2EYnQGGp
aeP9KRuIJ8Dg8/Sg6JqT7cbLhXbmzeZFOEveI8sNNqd2S1eysJ7LbPM7ngj6WUYf
g4KJ8kRfPSxDngmwMwD2zHhyeg/pEWok6rLdB5MNhMU+NGugIZS13CIforVf03Bx
qYeE31dlEdejL4H54Kn11ATTFZbmN/eSlD7z3QCW+iLBjAgf1p6bav/ktsJ913P9
cqRXkChKXlL4U909hF4zsM6KoY+Kea8jlzp15eigN1MfuIJAZmZh6JlwIFghEw0D
kpF9j6Oa/SRKLkleaba9PSMHbMkiL8IgkdWfzqLrjsugATjn0QM6BodiIK/wO7OH
9wQP5Tr2GFbOIOuQCaWN0nDpuLh/I9+A47zU3Rjfzyg4GtCAjZOtHVyQhjj3duK2
It6ChASqyPN4KFceuV3zVZolaWBl1EUG5juRy2h73LaWtQJt35zqNId+J/5pgWSF
g7vZ+58XzvNoSsJAR+DHqFDqFyEUME5Dy7bFcfmpnyd9FI3hQtqWtEmwKe4JGf0D
vG03N8/poSHeThP3xW956UesmmEL83hhl5XG6Uh4IR/u0I1gC4n33TgSjSiJq2TV
kZIzzZ47KPgDqHobSng2/QHGSMMa02ykSr/uDDTrCtYB5308gm7mnSfNSEVGs70D
AIhZETOxqx6kx/AF3a8W/uRRCoeOrvchCDecvjyfb9S7lmfNmGZgUr8ELAoUhX/X
P6niiz9izXJfb0AK2/glgjyxupC9dtJO/wnVNpMD1BRn41t6rG5mnkZO4PJtJCic
b1dnhPVQgDpibFCTRJ3joCUgBaUiS7XG9ZSrdroiQkxHvbkunIxSnYG9EtLm/4my
cGoptSXLJ/KCajACxaZNsnvn83Yk32gy8KGU0gDQS7GoolRCjJqch4N74n/ecgWn
iayE2WAQcy24LLGt76Ib0r7T/VgkgLXic5AfxDTuDx2/D2q+Za1AULud6E3+Gq0U
aV6W2i4T8umHNL0lO12oC1Pqa4OcdlHSgoAAUBFzbJPBEu5w1JFdsacWLIPk+TM9
Nwhmyvz2PiJaf0XzmZj1UPxmq7bZn32oCM7Rrj6VcldivjQzPPYi+qXBFJp7YJEh
gcT21PmadrUFvmfqSDBe+2EkMkTNtMTw0yKqHvvdgCfZsasPwBQZZn7ut0vZzBaB
XKcSdJRL1h8EuRXt272fIIrhe75uZnbQ5E2mxDUhMHnMqaKKT4yUAyZLn+kR2t5N
znTwhs6cIdSZGsYM21PbB4mZAh6PmhJdebQxear2NzdGNAwGmEfk+aD5G6MVacVa
VVMiL9U8MuWFB0BVh/AjB07kf8t0kpteY7GvpN7sCw8iLfRJ5WFsZojo3uC0rCgP
ND8t/pSxB8LohH7YroB1xchMHsA7dt5MgC+2Yngt2ZUBg/ojCix1lAq5NivmS26w
hY6wUZdM83NgpoovFZW92cyckqIAeEMrG8Hgtn0qxTisq+p7p8BTRjz7C5EcFtK5
hw4A7zQaHx1ZeaUpU/MFwf+kDDUWTFC710aZArnq2DBmGN0Kg5N0qdHkIyObFPtY
6T3FiwZDREqxUsP1MogbHqjKVSmRFk7CbabgcTHB4D2QpKSMxPAVUMzY8jx76jiM
/35NIZrWax8ObOYnD9Quh8Mgc5KxdDOOfr/5Gl1Xtzu/VTsi2SR5WZiKEH32HP9/
jIwlY9/8/k/D+kDq7O3XJvDUqyzQPRAE+VbMKr02KIzKT7aaTbNV+Tlz1vRDYRXI
CA5cfNZTeeQ53ZPKzpAdssMZILUMIGBCjo2u10ZDogElNeJywyOmzNfpGRVL+a3l
+azmCc+wqJnJgUDARsf+LrGJf73GAVCgfBPbvvsaWdNUQGydFosk1KiZKRzD3ad1
jjWgX6tkdSk4u27XJzzuSPpAa6v18Fet+Ca8bvntLRpMSUBmkXGxgpitnR2mzu08
0TZdnwMgY6+ZZKWXfxAYwe4y5H94/8DNr7qN2ZON1rQTX7EMXS6B5rNAOGoPUTjT
l8oyOIM/DZOtRDJPmcn+zVCDIJM/pL1mXOHnWd2SuTXy6ieR5oUgoNFyrO9y87yI
XyjPu8/TnwzIcZi4gwOX6s+GN7hkq2MBMoRXS0GL2qbAAIFHHvrZRclv6VVwdUt2
aIwAUSVKTKIAtudWtot4hWPeeC1BJgKdWJLpfMOqM0We2c72Wbz5f5X2APKrwUit
VxkVcmVBmieCf2ao2YZyzNQBuLnZ8Yht07q4AGSb/knMtD5BKgfsAvEkV9ieB3yr
KSQUNTWHMNpnjXFj+LR2IPJ6Fhte4k+6bOdkhj6kPc9fgWtaG/I6UDspSBbIBpIA
LNA9lwoM2td07OoijUpsBktLSy/UWUbM4zbts3IQjD8DE9vGtB/gkWOHT0UUkZC9
dUl3gPFrPH8N17ViUoonAlrQV2d5NbhOHgyKGDfBkMcLvN8mkTPKst0YeTo8w2lL
5V4SMbmp32FnuU3FPKkFBM6ZkSbMb/WkljV1ysgMA9tk5h8q4uV+abTYarWu77Po
yiKlYapOmiVyjd52OW5xYjL8ORHBbrXSF8r5U9Qza24fmojyX5ljyseNkYiB5Phx
vi9yjEgxDSS8bprPOcgOmWiI1xTXmtVbvBC3zkjF804yS/9g+PZXiQRygynpqgwf
85+2mgg4h7/F5Kk0hhU/4ykBI24ljyYcAd4MVIUDsDmMWDhah1D02fmOsZfNw6vh
KDJQnuxLV6V4IU2/toZLV7Mhey7Z/b6qZHtv9Vfqrfte2Hs2u7z+AUlrpIx7V2i2
hLQ+p2v0lSjkM6b4rGnEiuGSlQsNDGnsDDG8vnU9b6eXONnNqMETy9NaUaayDCwY
ySGRcg0SH7YTnAISSoTcIMm7OsCl6I/Z67dCia6aRioY430xjp8ZMX5KLINgdVfB
NP6OqXWY5GGUQxSTJ2zVVb5ZvJvDtlp2pXbIfXs9H2KcgkNwrHRwQ1YxIXxKJYNa
1fXK49eyTCEdAJmYWQPWHOIVmhNKEsGzqIgnRNbRTuPSy44QOibKP3I1bZoKT2HN
0fs9Ck3KtNxMj6sAYcjJ0QWMKI6iY7aVCdaTi+fhcPGtlmrd+OM6KH4kUTy+BtqS
v8RjP0hF9ziWUqdaW+bcU/HijUpL25TxxX9TfEngBtmiaSjhF7IBVKYOmoRiDW0Q
auqYOXaykJH1sdlDRGzABVuqlCcZJg2SDkiab1DaS87IkRlrrprRrso7Ow0Pi578
YeNTSPYFESDAFa0xjzbTO3nbGQ9yzSZ3bpKpdl9kEw+VQALe+JsrnO68jVNbxuGs
PxbgEwS1SRXuiTKsjLaBM+3KF6mVD8InVqp5AIoRtBL/BHBECHeSWi5KEr9p3yJZ
Bq7QY8VdIxi4UbdFUkDiZ+P5oOgAw6zMyWon16AVbwtDlbYEacVBp5o5PioD8NOm
MTNDHs7Uw3icOZQy9MYqo2hCo56W/PChf5M4iOFRW0/7661Xpv8L2jM5TVZsAQQc
Mv/NUisQu6qFZsceo0CGrp4bpd6peK8tS2nC66m/njjZowmDAsAUUbmGUUOuFS4H
MM9xFjUGDPQv9BELEZMug2qVkDS5c1Q9TSoOffo5bQyePbbEvwCZgG7oU6MStt+R
YTtDkks41h4Ykl5LW57Wjj2ejO9zRD6VFWbwVOJIjuef2D+CHJrFs0+MlquRr7Av
KDkWq0N7xZiX+sxnli6o5GgB0Qtb+C5+WuQQ3+RZq7m0zKhr8YNIycF6QoWw6Cr3
9iWocYVt41s8o2LqULEG37BkYQwhIxJcHK29lsJ/NQiqU7fmpCYZJ/IvZlCyBuUq
0gIHum+eiygh4a+sWYQ9sLfpt/mCg4oHkmNQDr4F7NDcAuW0kRiBCyUpw4V/Ja47
u6/HPvpiVcLZJ2EURbg3PnAZnfGUCsR+y4G3dkv6Vn2YCV5dE1KQV2VCCIxszbJT
6RDRC7gqWhGRTp9Iuema3bvPMvQbjmdOJwVOHzE1gEBOaRugMOgGusSeniZ9wZ/z
qRuGHV3zHJqrdLN1mSWVQdhNHiFkhDqjcS6f6Y9Sl6CAMZVmicWnEAnKVurWW/8H
Z6FsRkC9oRJV6zw7CKA4zXqmCpSQP+CUjTCoduPVxN9UeqszyvLGcNLTawI6wdwq
lb+uRjkaSCM4RJ0SoxSlzlZjeZsTAJZyoYdjRSTir6UMqcVoA2vys2yqb6q8A8WO
yNIwiq4GIcgeN2o2hhM5QnnLguoVjkO47nKqgXPDF2PKLxwvhZJuL/18MW564MlK
l5+g/OsLo01g2igK2gTJW9gAJkUoIi8vHJkhienSxxexv+les4IxHamXGks6ADfr
SuwRye5XqrldoLuM8adJ9wZnXPfGt9G3NQrn5aZC3uez1sDMEzchmY7S8HIxM42A
uUaTfxl/LnhsF9aOBmmRScu8cm25MHW8cu06A2Fk0XX6puow/MnN3HpiJpx6/iKU
8TTLAemxTYvTmsc5IXBd8yxMHs0AMUoh02QeAf1Z9AddaOkxoRG3WlMOylWga3iV
J4dKb8u5UYVNsibhuOziY8EwZNPp0DtZzIbIf2LG121YcrSyT63IXc0fO4tyW8Xh
rZW7JJxoq/2ld8MNeXR6bGUMPxBwzQc5mz18vxRwdQk+O8awZJKg3xJH5Ji9QtcN
pT2jx+2j3TvhfHiaFIu11yxLnBtTGu1DGgqYsRKE+xNUNbK/3/ajWJkY1XMirUwj
d45PU8+Xy+ecWJ8JTkm1U3Bj+Tclkg+eehk0Zv3rQJjYVTcszLX2zv0IGiAE1elZ
HHj9v88wlQydjTOZjphZZKdP6BCa7ippnsYL1acAGvhhl1j+09yeIK9im6hA8P5T
YVzkFBgITeYolaUhuX+I7cbWJpwIxUNZl7bN03nPRkPYWT15ZefhpgX2QmcYRekC
jegcHw3lV9roBjFTTbC/aLs1L9DOXcrjmSxDb36Pm3PV1rK/fMmPIbz9xqqL++Jp
1oDZG88gsX4Y4lsYDCx7JD/6zScLcZqgArq16avZ+gvZRkA+22wCtBZ0L//Xilmh
Rtms+RXm89LuecZR8N+GkuhMTk/DzLHpohJeWmRGUNBhHH2F3Y/vp0flXj0LGaNZ
tBJgvD7DkHJ/4jQVQGp6kpUv9paI3SJRAdJFyGS1BRa0nG4nuPrQZt9wE1zUD20N
WgkqF8GFTRTGrPqidUf3VtfyExC4+bH7LK/eOK5aLwrRGh/rlm8AsbRnZDV7ZoAF
7edu2Nppz+OFA0OfXuby1dvEm09yvsBARRwDs98pcMadwvP7bspHX4So6tr/0QJE
RjGh5ApeKmB4va6Qoih6teK3G5wgK6nM7ZCxsCtKULvVwEeixDNWnLMiC/eC2fuW
Os6+8pv2DpKErhf3wSFDXaBemwFKE8ZUoxOc+5XMAaG2JiWvrJEuHv35T44Vjqsr
nxAbtFFxo36ZUoT5diQxWta8qMXpjntQOE1cNXYyYi1XLbe8REc3h11pfvWJNBJP
3E+UCzHFjS3G2B79qLFAUzWLntbYkrXbjzVpubZ9AFxXhVw8ikeSkziBikJL0VLM
Vi6K/Pt//cKUlRooKr3SWvzBMTSKJ9Nibs7qfBWZl1DD4djCadvg/uHP445itnQX
qW06ndvsc/VF1wpW25dUOL1PZ6o9bTs7tW6PmweHK8g4J9yvBbHuZQ+GBHK3TN6G
sLRn+6mVTRObsuRON4YmUb6sVlH5Hy6YNkI9R0ffVK8iArPg6oU6q9ldh7u+MBOs
35zmCw7LbdxgZgs6EwWGch87r7DftgO5vX+2DmJhqR31UnFxjA+KzWD+zO/nVd8t
ObRrLYsqTUFToI30JQ73+g8kdkwPljADMZhzMANyWwT6pxBx1b0Tx+oIO0LvGH+W
sIqnOsYocDoVf4ljoY3DvpsqfXY+5acMG5v1lj5e+Ev9HU+uoS2yR7tG5ygpjkgT
M83q/4NMEXi4XRa0OS8+qYRJ7RDCp0AVVbpZvbTA8DnnAaUMbIQZ5nycH9eDZyR+
zjrT7vljpehRBbYV+3C+BPpUCFzxlD1zpdHKxPvuAbAdrEYvI4A4P79XiGoQJSVo
aPO4Z6jE5+kV9Wj/P3DWDnbOMNFavFRwSjn98cvD9Xchi46GR629QmCLfxiYomg7
bo6/7TC5fNn96h755H2qxTGoRONaQ6MSnkUoeAsvyG1MWwF0LKEGAEIVtogG8qU0
ujv1FMiGCZdRpzqjVDVSy5g7BYXzXxDK+xjcxod4/duQjBNVvXPrsUaJ1+1dAjyG
bgDCjKXO/mL7o5tc6leXvb5/T/yW3h0NRiy6ByZzD7AyIEs/i2cShW89TrDgZe7k
whjyEukHAEfedgnB0JgKmPgdclkBO5oNZsFB9EdiBJiisw+ak7EbgIDUNrBpuevc
HSs7+x4Ec0xMAVjJ7DEsGOzdTzfgkN/EYnA4dV7sHe/nBqS6GbPWhDYRykZ4l5UZ
gn5hnlCbiq57eZWOaUYVP/0W7wpf3TD7x8gmvk/D+Nz3a2/B+80F5YLOBw2nfLFi
CCjMPR6KKpPQ0fGW5CMnBrPnUR5cv76SKN4Hopz+8aNP9SWXqlAvhZHYwUCWB3LI
VJ5kQvNxErcj5NZNzYwwtk3XTREO5KO//sa0WZk9hNzpv4QvayWvtCneyo2T5g4l
pw+baV0XkC43DqHm2CHzxYHODnuvPP4iohuGDHHzn+CzegNHub3i0ynEuUdnKkyT
Ky2X+0GS3nZ3ttfBE21AFWIZzXY+SoWVgRHvBfsj/KKjtNpW39UG3ALedwe5jftE
GoyzVsb3MUvACT8uyFZEO+9X9torYkuITpfMhse0bAkLNojhmx2JxtVDRJ87MNjp
HFj+V+GPHTadYiHR4bpLhlaiLHU+ksHwsyS/v4FyVi68f2ELZVg7VTwrKOAgjVJN
mOOMpdWyYAL3ltSz22cV+tYL+YfcR/A9Z9IHYt6YP2qf/Ld+sARlu/bxBt9Wj9zy
5BUEB03AVXAZdaugLjCHq2YZ3Sk1D/HkIdJTE2qlfykwZ+QCy3Ash2aaiIfKZ3Kq
Ou3H2Y4tPCvoXRQDRsGVLjl3TsK8elhG4DY6zbr9waejtVW0ZDmpVg4hZjq3m6sx
8kSbUifT30+9t2Cv8fcgBEZ6HLDJ1RShRMet5sWVSkwYWHAzKc3TU1xZX25gnQEy
q1B2/FT+bmmVTrdhmwo8U9n4yeAJxmXXoSkU5Fuc4Ygxa1TCaCInxNn3uXx5b2uW
TqtRRpYdVslnK57kaBYjJ6Je7fHFBdRpT15n4NuKNAIVdSkWWu8/doMS1DuPQzPE
912baXfQh5TLPkDI3PWTakmZK7pR0gT9tNLR72PJI/ieKwColew15DZQ0VOdFmfu
IRdwxeSh2fEKOvp+PJMM+k7aBUuB2mreafIEa+AqsygiHyJVzBbpe6Z1D+tNiiUH
rvWzWfOHWNuD4uOhnlGZqZniIGWrBP9BrB8UQoK5VGHawdT9DhQjJCsNGxViyxbk
ztkLsvJ+b6vXr8SIuBuC5Z7nKDr2GUycu8hCCqkHhLQQf60ygZs/WBeG2rPcFCKv
q1W5XzeQqcHvzB1IcgcfWa77fmfepEESv6CPcmi1hxaBezbVGxuTspss9L5aMtOV
nNkEFZA0IcQfOXMbmNaul+FAaHdRqbCuCoQjWEChAQXoT4acs3ZrD6gXDdFfEtWz
AePEQo4jBihLhR5U5mHCyx9Z2/p+r5D9weWeOyWn0gcN4LhgPFAcBa9Lfm4C33ys
vTg0OmN2btHzhTJg87RTv15zpd4oq+c/oTgmf8z0011DN59Im+AU9rni6fVQ+Hqh
mMkk4ik/1rPWNFdZEIfw621UUo9GjccFSh8XpkuJZ1VCgvUU8gNNQTTGz/Xldu4S
O2fXdsxn38CtPGVNVWDWJCx7/HDZnOxFhCkOSXTIIk6fclFZQVhALss2E3Xl7nPW
TjVHS+uOhoKaNmLAmKr+iPyIfvLNmfQCppF2tTCn+HOh2mWgmaipRoSQ3+g2blD2
YR4SY4R+xatfQfqF3ZnHqqa8AlLtbTuPyM2wqBCOJm6zyBRziXaNn8Wc+3saD8u6
GiEgBxMXnxjpOTnTSSCkUStzWOwfHAQdtI9ZdfMHZxkkTH7uW7tHs3Anz+c58kia
O5beke3+60PUkhT3YXo7l5oiJxWDbdu2eBC4TmRbh4PrZIw4XK89xD2jy2yBdcmU
ZXI8B0PBwjhPkZ2Fzx2KaI0nxS3Lp6/6GZb8vAa3trB4c6WTJHoP0ppWUi8/ThlV
zhFHr2M6eWfa1OH1SpLpne2zAuAm1sYMLblyc4TsgvH/vD50KMnpKR2dMaWjYcPn
zYlWfJha0ivBn3ZPor4A8YIYbanpCJYnwmoXeclAU6hK/ayfvl6pQ7nlahG0uPB1
tK/gYVq+hCjVjLaim48eWlp38G6P/6w3IvZTOLtID/dr83DczOuu/CwuG0Q/5AsU
ky8S5OcRcgvvnbEEv2JbSqsUZAfjhGwqlCKxkG8utAFw3LVbYPj/s8n73JC2Rybj
IF18pon9l3CmPN7BlvDCu89S2rc+eYx+17NtbByuCu06NPs69r0w10zRNXyK92hd
m5bfNxnq1lhxRvWVzo1q/rMKboRorufhO8sQlSNBchCC+4KK71YclGOkCqKL7eIX
r7xPrRdWVSWdgDhn0tideP+w8Eatc3syzfwe3AtakQas2iuvK1W9rGkTUrkPp6c7
bDsDVZa+hVXmin5VW3Z35oDF6rA2j2MvoQ8NYXXCgJO7iw+Za0tHwtfE6RmBFwlR
1SYrjZJM3GfC2ovfBz97IW8SN3/SoJisLGbyDlmfDBdaUhduxuGNbsx4j+5QOgOu
Ve/g17PQrx8DkU5bREmHIASXqjc82H8YcY8LaZqH9lxELSrYyy/G5XZStTH77sty
9f+v5i6AfjfK9bQUULx80BXuFbj+uBl2zc4CndsqdF214g+biGeiXulYt9S82aGl
wng+NZJnSqk0ho/g9ly54JBxW+KQ7pZmstJHAC/P/J/Z6m0l02xugIjGcadRXQTo
cUBmag8h7zj16XGSQNI7MVZ4oMbw9UKdhf5OWgFS5S3YwTbUeSvE/0OGMcaH0wOC
Id8tTMLFtNBpUVNUq1ve1H+kv9+HiU2lpmVzhw65M7dKrshgwHg2dO47NTB5D3CO
iuLNhHi7X3Af9U7SHZYhV+8KLwQv0UIGDy1QLfdIBqcX970otMTAuOgHYXN0srhY
uEDs+XpUnCjkcVfOUcw3c/OCJmUuXxBfwujZBoOIAHzC5Pxn3jjRnlF9e16sObjo
LMqyFYwDsBldsCWYiLxTG7egcojIj5gHy8rfRSWo31LdlFGk6JGOEJK5QuypogmN
TEIei8YhTXPa1lQRTfhL/HdMN0z43zw790ikuQhtJ3OBuHhScv4g34kjMCE+r7/Z
aLLMQjEpOB31NjURqqzsNmGGa9Emr+6/O+bAO3sZkldPnT77lvv1vBTeS8Uj/X47
ryqe+ZnF7cva7Ja+7Tlg+/llZdQfI7m+NKqo/gWqEdPk64dtO66VC/rYKPr1gDwH
rj8QhrN2j6OvwSNnccPN665QtQFstZ9r1HPGO73PWNN4uYXCHHQ1GE4DfKTlQW5O
Unptl8P72BBCqZLfJwOfNGJcj0lM2rEThCneNv5nSVNbMo1Bh5JAsnQxzs8GnAH0
oxmOd7dNTRqouyx7ybBGHAKD36aLkzmDEYormZOfYRgZVfeOKrUPH9JMCpdv+CGC
+Bv0CQz1+yZDhNfEaRRFCeznkhfi1LtKksbELBN9r77kSi7ZxT5k4AFgay7anskI
gIbsrrENjLpj3te7hTSNX9uyeO6+nej/qL/jDJleIrWjFE54MwAmKLOwOnehP2KN
74Xw90vDyy3+MZ8f8xBCUGdBc6YfJY4fo/PirBpAx6ikd34Ffe2ghq6b2zW5Ztn7
1ZtD/3UFssmjjIWkSke+oUSixc1kqa/U7+O3NaXdL7uiwCix+KfNHHgRvO2bj/je
MQ+tUstXHwmDvlx2rmiYXmP8jNFV3pAOcdVrmEi6Gs6UdCzPtkbjESbeaxLJHc5L
Gkq43oZ2K6dRh5DtKDm02ZLdRJd/u3Edn7TyCo5gjVbsLNVumAkOZu5zZmptkZwr
UjAVDrytTiqw2DYz+gQqaEFL+vDm3x7SFgE0dEm6G2bdtGt7/qy5fiB/iLwijeWZ
3ZMCwPqhGt//7E/Jr0c+ebZF2OnvwTtiom8Q5fKg3jUzHYhd2SgPMqWAA/mca6yR
iMrtPiM2CBQHgLdBj/6O87CeOzpSN97Y0lXzJYw6X0xcsZeXD2AlyFgFUjqPvc8W
ANjPAlHNs3hjoWEvI9D796fuLPfpc9j+1qQNVbEsLrUyUKOP9z5qIHH1wWKULNHB
pUnGf98D+c9miK/Snb7ctfubx76UJjDC8uD7MXheNHXBBZX8eYKOJBqQkXAq3NpQ
9ec7j2Lptn+cEqdJxUhlsC3zrJKl7TkUurBJ0q3moAqu+NhsLjUcOuhlzl9BB9Dc
qrrhNNhwQTC0lK8reS8smUvscdfNOd/jeIMw8MbBLyZVU6qrxw+Be9LNThtUo7Vx
qY/sM804TDPgQW6xo4EDeqI6DdGA+r5rUv63zLvac/arlZ+Ozx/EG1cOG97vvLlD
IxMe3RtNSbr/GS360fK90CW+UL8bpz+uaAItmoTXpC/ALUWX6lu2+HDECHwnjMzG
u6SMZO/SewoznBHzgiQSOJpa+45N9ihsdwq0B2shAJwHxDDkHgTerSG6Wk5npex4
gcM/dORZ3/ghgJDVOUB5ScMeKSB4m0JhWVXodCcIPlQquuUCj9HibOotRJajJV6e
FhC23P3fpuDTT2JjV29VqkV1J00UhIWKQ4erwy+N2NRd4QvoV9inZvv0KqRewoaY
2RQOWld1a6FrAxpGNSUvSCIbNm2GyUeCoEbZohDsBAJzyFPPpG1GaMnYp8ypZsWM
GKC/mpncb5Qy1YGRxS+avYOAb3IPIM+eIGWCmxmrnloszE1qGOep6o2rAFsuoyZa
qH09+nBPDD4Ll5xe5uA28RbmXRMsMVyU3mhv+mGFLxFZyaNqdo98ZtHiLN4S3EQY
f3XFN5jLuEU3Wr8nopIS2s7AHItzjlmrlB1ElP5hyJ8Pn5UU+JOBkYe6Q8s9sAjX
2qQ0mPXSKxnFB4Mf/upFq6oD+FlTuVbiwSnKSMvmDNST6pG5Xiu8n1xoOxfqj3S3
Gt4HQtM9qjU7KmvOeElCHGZekoygK6jqrDyozcsyH+LZylLct181yilCLLNI/qsO
CJt8T3SGxLXfKUXwZKgxB3yeS0DkodfZUOwXkCzTemHkCKvWxyTpbTmzt8pIzeke
pBiG4L0P420KGhXIzxhi/ynWr/HFZ1J+xdGJPdh79xOH/wK+mMOD7OBxcc2UBGqs
L22JUpmc4FjJMYdOw9wZvQrzRHFcuQccE6yb5m7+WOJkNx4w0AnoIA2jDUUZlshG
N5icB0KV6kSVp33XZtjb7HgwPjVlNhlx9dXXT4To4K6/vms09sY5XDEPQkxwsNYB
Yqwe7+H9mCZy32GxAwkZxaesZFBMaSgRiGMVs2Z7/m37h4HMt6Pfnxl+sbvHLDge
awyghzg0B6/44Ujrfe60cV1S822TqK/nn/S5S9tQ684X3mJQL13k1Yy8ct1UdAQd
eAdPaQjGDk408oIA0yplfIzTxCUHbbd+syXcRo7m7j52F/Yoq/Zey4QGJkgfM+Qb
MYfX5YQasMmh7R+DVGwJkrU7e6MafsSBnMJWVYwjiaEzXXrVCNnbb5dg1W2awmGT
g4vcxxi/vKjSax9Ahv57dZZBUolXjZM40DEghMxbGxwU49cEGBnuJ9CPHOAtCn1O
ETgrKkBdlbDCcf5Lsne1bNwcwcs78lTcErU2l60HMC6mp32SBF8ouLQeWRdj2/6v
Um9pQQumC1FtFzM5a6iiV2yODGgR4Qv/oXZWw6PTp3MdwzDY3U5+3NjpNmWDmXcv
Aqvu9YM/SWH+0Nd18YDL/dSIdB+TEt0E/3cwwx3BR1I0d3XqHlDnN5Zjel2/lsrA
wkM5fBSua1IMEFAEYwaQa3aPwH9c+VoJu6xQgqgvGXM9/CKYqjX4joouKa4Z0M7C
jYVQrNQ9K8tmKrJcnLKO9UBBKpcDrMeqoVhuFStJcRLjsqCu6scSfdXc/NR3JopK
TKAcncbI+ExrGv2TSstJp/1yebBEth13t91ClHiauakSQTaMVUnrjsrAIUVljeGJ
YCHdga+LpWYspimbn0Ny4PrWVtXf8xUo8UDqwgpxaYXnLf3ZO/nMXsG9/dX70cQF
EDcUejaVHQvrCC+V7iv5Bpa30RfFv0yhIUSX9L/MXpQQtADY+Wv59TOO5jtsfQh7
a+P4lTVlsyuEmrsY2vhGrqBmSDMKmW7q7ov8CQW4urtB8FM7tj8kdiqFMONN+Mj9
+lfGqAscptLDZ8ZywMGHZPQw7XZv5NkrLMtueyi6k8b0v8BYz0QDRdxsVPMRY1UO
u14tj4nmoT2odwOAhedZ0lWeRmb8E4DUp+aTt+cDHmK1m6m/RaYePJJbb7BzgKQd
lWzbeIKxh9zncQ4qj6/RXGjdnAIApfTsKd2lGDICXX8ABae1UeL7dZIxfLtUXv0q
n0XqKGpWxGuLUT0QNYN1UBYRUSGCf8XKFRFE6anEGbPWJ3Q20mmF7Bv9IIEjeTdo
ioPS7s/lqurNdzXSJvDKNXbEATMZG2sY50Ez8TsMWgMHE4mwkaEhYZkvw2kX2YSb
HciQdN5BnGpIRnBxYZ8bkUeeucECXJLoJAXkCwPJOi1Qb20FxGMn0jfU1YUMZsg4
AIG/i5AJzwUge6oc4cueumC4mNGachlkWnKWxKO58Qqd9/FT3ICkbx3jSke0xVzQ
imoy2Vfddt8tfFatolaF6c8l8+fo6J4Emdur3AanZ/Kkxz+ZGk29QWHvhtug85Uk
NdPTofqFFGwq84kBNh2CP+uqVq8rP5BzetjeS8WmC0Eazj36U8blvyaoYVUrfiZR
7hxnyv3NPbAFQMCOC4K3tBlOe4ENoqOqHtnNN5b/Ah5rbxQdGYUFe7HdUOaHjwJB
hZx235dwAIlAuCeUqaPklJ4OI12wH8p2gH8JOmyvAa8IL8c6cPCxhWtEuR3HSSXW
MB2gGARdxSxF3QCeNcnXWS3ctxeMVLva2wNMSbxe0NFuGXUy2kN3nFV359OGn+Kv
e8mG0ZGXjVLT9YOvlyIUKLkV0aqGzcOQWAtWdi2r911uM58OipauzHWQEelul1o1
Pq0N189BoCS8cljTunCfZR5stweQ1ismJPD7mICwCZvIOLkP1h+8gCAAOhEZMmWb
Q7G3g8HKRBCihSB9sng8VvZlcGb/TtASgh6hhs0HLPBj4ZDyJzO4nVP2zt2/ecMv
u6EzdOLjQP5BjCNGb5oJK55zss0oO8X4DzJGIRNgxD51fOBI+apBmiB05TmrH9Zr
DRwU1B1aTaAISpDn478MP9s8/a0+N9bo3ECYG796Ul0mSjrLsz/NFnwSD2IUaNNo
sSRkDSBLKB9hRxTGewK1fjL+BneTk3++ZWz/3vez8Pb5jWOeAHAqtSVBZws+7YAu
bYBMaTnEFf1Dh1EAo3yXY19wP16AMw5GJ1Gj5+2OHXwyL0WCIXHp44rxw2zmA8eg
26Zs8qWetSUbdgExaJjFvbc8LkkIcdUGiLDBVi1IVm9wgF6+ZBcKT0xAyC+IxMNz
ovwuL0N7e6iLT+m6o/r0QdR1cGMm/P4+/YoZsgu6Ye1pgsnuew0RFvMxbGKsXyp6
Iajcqy5N1PREC/O8lr8CXv0LgfNeTvROZnIJS3lKmSUROdhhtbwGjfyj8UtB3a1B
/0gTRk2OHz+O72ePgDRH9r9SmRPnMNMD43xkw6ONR/WntjvIbkMgOphdtXFNKsoW
3FmJQiMOXyaBM1zaGuiglD18DXJqjCi5nWD8jIQFoZt0ooavmPpVVXnnvR1yO8tf
eq1WlLra3vO1yPM7FTecy91XC3QOtriAIj4L7hoVuggbVNZdHrFUdU1tGC85G9b5
xEj0LKwbyHG4gy0XJ72EBpAJybHQH1YU7aGgsXE0Em83glqnlWuKb3/AlKc5hB7t
bfbeKPCwFTYekR5/STPRDdgUtQH2xN143uO2e9Slpyd9ceDczmTgb/cpxtZWpDv/
269GOMQhqOn9by9Xn2P0yLQavxMh4q/zc5VoOuIz1+LGt4G6NYoFJB3MUBndvRvj
g/gPT4/Wu+qefs2Fk5OFn/gQNJkFY5ENFKky+XLbgRcDKnmSq+txIX68QqnzzYOK
uYPJWMk7A9S9hZRpGOMkCQc5tgR7sQlG/yYNjKd0yg0gXP66EwUQJ40gGObr1Abs
1HJTjIuRBwvuKz2DjxqTDnbwbVOEqAa+z9GA6If3QIVadVfcSDDo38eRKloGD/7i
1Yh81BpMB/xgBdYH80AT8xngByY0RIK1/9wpGSF7DqrasSM+4s60RiuSWiQnoGI8
I6eVavNGXOj9OUgxgwBhKCiwpcdxuxx8VWwbJ9QL+d0T1SmwyxYHfuL+A4KHwA4T
hgfusbNoqeci0QUsStESmg970LYcUcBU2WK8Aqp5ztGldboemkMATmMaicdJrmqc
B7UbraOw55UKacnash4u+sB6GfYrmCeaEOGfmsHxUfMWLL36WckHriU32b85sSRg
JU4VpXWEuUPCxTsxjcmjbS4gMt97H07JH3/RYsRZwnL7PinDNKXc80uaeaUnyRYJ
w9nyd6pkc4IKIsxDQHjOvuwMpaluoohlYbIcJQ+XPSzVJr0ztIcSfrYlcwYQqauN
cGwbdayKdZ05+xzEGFBcaRIepQ7BtQCnIZhC9psbwZMugzTjQe5gH7cf0lvisLj3
eIKmk9BPWHg15kqHf2wQNY5PemUHnHFaZIAOno6swE0ZxcMHaV2OBghP/f7ceDMd
IZSNExCmMjqeiBXnk/RgUK9uDukKX5KrdAHZXcOQVKggL+rWjY+YxggEFVfH9ygn
PxqBFm2R4dmsj1Qthb7DmAqrRbFOAZ7R1X2iFlh8rw7uO2Y36n3iFWQC2xaiBLGm
0srOCLFS6D1q8qniUKk1MTsMa6wzzRWZuZgUASB/y0GO/JQJVyxea6sdfMQuPkvx
Diq+LwetnaHn4Ys6Qa3/auyYCYDsOmp//oRohMT4xuaM/PynCJm29bpAnIuPr1q+
b+YxAJds6Iug+0wRd3hWURjxlQP4ACrNRYiAlZVFBuxKebTJvidrP55vOgfCJ/X3
4CwIKVV2bgu51+Ox5HnSLAKp0HE+G26bmkbx6t45xn3Ner5/c6XC6VqpnMxEl7NB
HBw79HDL1a+YG4Kb4ccflJ3VeempRJ+UPLAJbkRryVmXKWhuWOswHf8fw26KFUwO
QqtdaiEo+EUD86wTfVcItstNdBOQCW0oYHpigFKazulxmGuOyTK3lE8nvCyqTdAV
zJcWIMvjXe30CV9K+ej1pdqQwP4WrNNVd9gtFd52B4UjJAgSt3Kov5S55QaZQOie
j+q//rC2EOqdKNBHhu9FCiyVPc3lKU8nqNZdaDxpBFqFAHt9gLVzbYK4+Jx8zVwl
qyyIxtAREaOX3kSfTFBCcR/igYNeEDk6GwjMbDflE68G+KU7AL4m6tR3sFeDtwRM
t+sx1ltAiwl0MFrS8dB9ASZZQnL356Q1UQbxhTXmigyQg0cE1K4rPWmvMtS45ztD
QjIfMvra2RISG+iyh4J0vktzwoDB065Pcox6cPR1mg64LspWky9wkd6gwdFCLKmc
rexYjAxGKcytjcpk3WDbxn7RiEqOUGDkYMrZaHQJThzBBG7J0dLhka6ZK8E8J5Rq
QFdQ6m+oe7vjbn/HQir6iwF9L/iEpyUHUg8lBIja/41XfN4AgbI0z/nf2DJnYG6W
gyDK7b0O80iqQ8irkwiC7seRaC7T/L1g3ykAEApETirq9Aglv+Nxq7sBsGXDOHYB
muAW7n3s3nogvHeMWQiOqJsSscb44WyszirfNsbLNH2v9oYXFkqyeabONk2p4Qo2
brfDhdkHjEShOg8hhWfrAScmpfYT02RhR/UuXheexzfaLiDNCtDuGFz55cldgRpB
D287VIjLBPifxXA2+KBhhmXNolBIPBwi1HNgmdgSn3jtZxFCVU6C3Miy9VISDLHl
1+WOjQUD88YodTot8rOvTeS4TNwOqZ5hISZOZwI6r2HAfdHrLeHK3EUX3+h6tJMv
6qzUC7MfuRRwV8kv9jT9cqDeRQazk2IS84oJYJ+WfgS27+H2SZVWS/4AEGRbtpQ9
L+teqHPefRe9rrjjxsb8qk97MH4eoeYyKBCG+gGsq1dEkp5u29uCoqwvGw9N/Fs4
+t5TyQGwXT9Q3E67ge+hH/XBEcECIZ2Xmq3Gn2KFn5hg66Ar/KQUlMlHcWRdjMI7
/Lx9xk+GJUeBydtBjQA42JKctcDiYKeUm/8fImYMNaB9s5PR+/EQgZBqZPM0q/AG
byx97H1l9pdouHaBCKiTnXO2TpIFExp24PBuI0BgbQoxLQitViY8KjwVHrauYsu3
GUDJVSI2A3EAwhZYK+e5DUpe1vRcUj2/lk2/VQvj5ctmyLh971Kzv7srLr2XFaQk
3UzylOOzd3whn5hGbonXquM/cH/+B5QVtXa0QDxjxS0kk4UBUpAZUgCDhJXsHpQv
uJmSvfwh+RqTSdXDXVaLxNWx5B7kdWm1YhzQ50SVAOniv6hhfNqepjDev8phbFvC
cdXgzgQ76AfKgr32kQNNAfxr6uBx5wTtd+ZAqHqLNHbsmL5b5T02weWauG8DgNTy
aidyN/P+W7Cd8vxXymAx1KDW6/0p8hFkM+oZ+yPSNISbP5Yi2V1QImviAulnOszt
Ud2VS0xNqQIK0ahD0/R11VlHoRo0krciHlVIee27GPsd21AHtumUqtlBf4MkRy8L
bwAN1NWBF3pdyT4zwZduoT+gbxvzGMAOgHdXK7sunzT4tj2+oBH8mhzpO6jVMonf
GcuOWg5XSn1R89OvsIW1W33PXqtZ0kNT9QvZt4KyesSL2PUNlcaROVALnobiiVvq
6JaOWavLkbG6pYL+QjRP8KmHiqtLzaypi2HmRAaMg2CLOJ2JykGrjx5/hEkNHLvO
qLrDRmZ/stcMJhr6l0DCztIBrogr9P0KJlBlIBqZGPNzQpdg3DFMSnm8/AfDSUZi
o7jBrxkIlsA7h/UKC7sDIjvd+J+XEzR+x4sf64vZShvwlthp4Od73XCRCkSLQpEx
r0cBietUM15A+SPNIToXcGPIvXmKIyLvf9/ROhybIe+rlv5WDFerq3krRbbCMyfM
Gj5VstBv9S4vavGft9qVocDSXRkGnlDI/ymeAUf6Vn79fgkvFj83YC8KIEAR2+AE
P1SgR/VMIwV1h2b86KHjGlkHZePPxWcHJcqNm46vZKiNEKewizqmCJ/bQ4tUyUVw
GDA92OzvZ6o4RLNlkStyYaufxiAAUgSiW6a5xm0PS2w9yk2r7ydT7CZVTfM0tteO
bFbyZdyn5IHOuBmu9MRiLhLKcboNWoTZfUiKQiPEdvw1h+ZvxRoeYOkrhc+PsTvH
7vDIXhJgnW9/hQ2f2jCsCRHa0waUNKrUhW6851HMGS/xs1YHaDZjgll1WPhtO21K
JbxeQeDdQ26Z5UcDiyit/BwFSBXI8uYFfZGtq3BFKc72ohmZNsxhHJGStbDxT9CN
O8uSiENDQD8M9UXTUwD2bRBtSoVVYuqADikxVekVrHJf24d5hUj04EqA/y4sdGHa
KzO17oe9nUZ7PBRFR9m699RQ9wu6dK1LEt2gPXCkC7fBXR/VKcOl4DOoRWSHGVfF
hdKh8O3wk9zTOVpp+oHQPLJRP16BCvurJgoMWvWHcmKemte5Z9ANN5pNBvI+qNVp
mB7h+RZVEuazLkQXbmP9JJhj1DH2+icWYT6zhOvqiNqmEFbGqK8EKegdgw9mu+dV
y9UmhLhkIRJe8E3blGBzGp0EO6GIQkvkH++symJMAgrpMErbmui2ilFC85OtpFY9
eatUvFjH/j2sp924FMNWw9POROSGyagV6lujTBEUVCHJfi3cJrDEcMFQ/cHiEcD4
f+8HwPqlclaY8cwl6M5Vhkp4VUxPLHOYX5XQjWnuKMB4C2BUBSAsFMv3jMgkEgJD
/PVtdLhibAdxwr3BbhA1r41n8FAY9Wk/tNZECmpOUbrtCK7vB0wvTmLKQkOR9WIv
m4gqmewZ3xYsCRWWYMkjsnTQ33Nc9OtoaWXkMR4DNf1alO3XSwNRD33pg4yfwU1B
iJnyhp69FQtfuRtEXKHF7f6Rizfw9PAjc5t/HYpDiXOwodSJmuI/VRejEeqPJ96O
qI99/uCRNy+EY3AVI+lsjGl/xi1vlzbYUg12UlBKU58MVd8+2lOyrx2GBDVHctQ3
Wq0ncD7MuNH8lcgLrszznf3fTaIG3hTgQVSDTwJ4jJF7NP9dKdsnnK1JZ1MIixkK
Zi/8dG9ehc7HrxtzVIdzDSXMxe+f3E5dPwCG0W5Roc8wjMAgFXtHnuDvmJ/oF+tt
AJgY0HuA1ogCOzeWqSIDTEMP0jric1EJGXF05P8pKf+QdDGo4lunXYJM0R4F04DQ
U5UD8dKB+Syn4BHP3aw4AlYL6Tmtm/JsXpI3fS5P6h60khOxufzSAqsJqiaXu8k+
X3uzhua5u0l31uGzE8YIOmUvI3te8x0KvPwJ129SHDrwUF9AeoHgsLMsbnhNGcdZ
jB1fvsez4VFh9bNeiQXBuMji620lUaJ5UZ947nHBPGVAa4K0CzOqC5+KWGYJ46s5
F0+xUSyt2H5jF208e5/aFBP70bpBYxYluuuusEkeI6wa/a60ew5KJ9ZgPBZJRv+v
BaFTHxVPmwC5fR3KRSM+SwcprhhCIs6JFLxjNnqHhWqIhHpai2A8wcc7pBdpBVVs
mz9K0bIjlh+xVWeFLy9HcPZ63On99ocD1++Fi4zPtmC54kZI62R4rG13ze+Ucgd1
35wuq0uMViBfEgqcLLjzl34OEfiHTuCbWMqCZwcD9NiYuh65DTWyWLE9HezFosaX
maJk6mr01Rs4i3zsjEkkWWDe++j4L7bxmHBLV6laD64M+FYjDTfmR9Zy1UECBI6m
qnspPOmlLpEm9WL1+7rkFVKf39eVhICRU2ON3NHtThAgd42EaENMjllOcC3lLAQu
1mHn3Wnc9OlyErPpxezsqX5cYFPoTXIhLIYk7eo5BZ7bCDihRzQviST7K7dEKv8g
NTP1pYxfoBRtHRBHdbt3WznonrONi8NKJ8exnUs5IvMFglEgcsOfw93wkayMnGSy
mHlm2sHpynwAryo+qpQtlkbi0i1tLS4Y/BJcc71sq3YC7p5dhQ3nFbh/ecgVl44y
lJpHogtzDi9oUe+bnpYHJZAn8xy3MlLKfeoWdbJh1wDFNeV/9lZNybaRG4F4nSiH
YQQvqAb08pnKhaW7xEo0RIoHmS2CylYxBuyS9X4BtKZEz6wfVNUyUDZVrWw0ijg5
18/vq2ezkMKtRB6eNHDK1s80qIOnCE5RlOgerHhBQnaFif1MoZY3yoEaryFcHI9x
o0Sz03SL77pGENVR3zfyMFYfR+5wi3rU61xKBb8VOAdvKlUpLs9pa075Mhv69kdM
uKnT5PzWF6kgXCRZHkfChW/63u90htI4PBkYq+0phSEyzDlfIycM91OrXdHOEIUZ
Rx1KUkWqX+4XPvPUqHnsp1xh77+bVDia1YQgBEzw1Wsc6099RbGtSNJ7QFhbpg22
HJ/lYOrbTmrthKJv3QmiAVdanGxmUgt3MF4c9/W0jHGjHJllpXZRdZAi/Gz4kmMQ
nwOksA+7KxtYo3wHoKQU7PX1E/y2/tItHDLu833c2IdGl6kLTYN+CmaDMYs41wAX
vjlMrcXl+WdfPqyzSK2P+rPAsEFpkXPMzUApMVq81bZBDrAFwlMjFg8o0oHmxQ9K
psMKJd/PBqTfYPV86TPh6N9CuaSXOxOjiEdJW/VlC+m8eD4wyKs00Piz3KdFKVlO
Z5s31AK6bbropdloZ9sz3RjBuSiZgFCVcDejyOKywPsPvwgQhCwhE/zg6KxiT8Yz
zkmP/0BzAksrPBpBhV0nsA6XFsvvAJQ1OSRKBiL+Ek+DO4Q8qhSbmEYwwS6R8skI
ggEYJ/qWvmWITNtR39r4shaTGDv/17EwYC9yXALMEBr/1nhjXG7p38KZotY2qriz
FnB1Ax57BAo544HrhxnoBqmBkRzoqU1WZIrVRc64hX6CpSDevtWjmiLfqFSsb5oC
4o7Im3YtdpFxNWHq3dCu1CAl8AsrLpOVNaEu7L8h+qxP7oPldm2FM57BpGWQ3vLW
5PQa039H5DJFmMSic1RF10mDulfqFgoLNB4gOqA15r/CtmJ02F3Xwj9yafbXG1oT
JSsWpBdwtFGbK86btm4q3hsYE8PAxPcmAaS9QUlKtdC3oqGqmbbCsx8BVxtzMpXv
8Q9mnM5GXmB4hZYToNtCK0kOM1MssxMojlwRVwcrnHW1btvzkZYvHpGiTnkeJSVp
Jz01LDPHP1mcxlFor6pFq4L5yG/Le04EbM19jivj3kP9hBq9pKR9fKd9tUNL+PXI
8sKC002z2YE4wotg6M2OuRTVpSEwXTrjAn56Qn8xWqu0Xpg6JYVvXipmE/VbOgdW
tNvLLm93fYf9rfngKlOpIbEIK/AhqV2prx0Az4PK1YjuRgbLVZ7Pa4/YdfQ/ZEEm
m2bflCvwQbaR/YjgaIAGmTz6HHxRf9cE6SrkiOVwwxVtcHCTBmmIsbyy3Rl96Fsp
0NEjveDUH5ITPhIMsvmtNjj4LAdKMu+ovFjnXEmeIByTjIuStivV5l+RDq//7X6L
v/Cr5KcwuuIVvI2GvR0wrlPjSdVldvoArmd6lsj6tXnMjtKejt1FBzP5wbuzpE6C
Tq6JUH/fB3ac/CEN3O6Bp2F8ZtPs7ee2Kt60bc+HvUDOVMwX9PRLDBtbEZMd1uIM
tKWTMe9jBF4Rtep1+sH/nm7hKyduAXtIZIswQC13vtFHPixiOP2DCygzkKWMcG3S
JeEfmh/AgAijYW+wopVIQSLNyernkUFWkPsjnf7tveFpFW1zuE2sMqT3v15Y8CK/
UXqI5JIhqVsYw1SIFh4lc8k04mcPrTB3Hbf2SP6QEbiuA2wjcVHFA/BRXyKp0W4S
8F9hFv4jNah2LAtkccOU16t+5iT8m6dzPLpSjMuYS+CNiCqmnQ1SVXbg1SLAZp/s
HayyGeer36DnqIKNRajSQJLPds4411+VXxiTu8BsaapjgbYB1dTFjm1D4azCrF15
6WLoA4eDIQU9S54OtKLHrWbucP7I/KI49surCBTRJJGOCrh0UgiiobAdSylEPBmH
8YB82MjpIE5eh9u+9PIcFyLhNwQAVY2gzecSvf95lC0OCN546WrUJ6SzQPwXEt3W
KyzhXTgt6D3rTsjFBfgG1T+xsgrt7b/aWwsWG+Rrx46k7Ku1Qiv/XFoOykJFah1S
S8mPgJuhC37T+nVGeoJckjD9rDl2fQDgIZybzyLON3hNYQAV4PH1QV6+IDAzWrFH
i38qnv4qh4xnHzjwec45Pbm7bc2Kz0O9P8n/OwtSUh3N2rR4iztmCvwJts9vpUOq
EFC+HIXqa/yYtOdeVoAHwHAilKmtKwigQiKs7iFXcAPQRtfe1Qttogy8unjPtxCC
3/T+Uy8XptNqfBM2B482yaMNhZsSy+co5HaogfXDDE1lxD0svoKSW56BrB+NhWIg
3wcwZaLCXR1jIJV0/MHo8FglfTht3q7OnnZS9t+LxpHtEDBYP/lyRh6T1RA/1Rgj
1dS8cY8J/ngTP0vXxk6ZJCVRXYsiERXbRMBWwX/T9kR9UZyxiBs0QNN/33iJfJXs
+iuKhPA6N0xMq8LNl0Ql/JC2CrSOaqPYPYJLpwXygSylI9QXZU+102CnqIlETXgC
5USEaSzLsZtSxj38ZqbgChsxK4/fkcQViRYOXSNNJwW3pcJQK+/YHld9GVOUgUuG
PP3mT6VDHBdgdH95L0oNAA7SNxoxV2NBdbOxG3OYwO0gXPLHOII2GsBjuy4uXLvE
gB91CNvQdqCpmRokMBrL5WanDxd2O8apCgBV9Snh5aLSW1moG4BXT4AFtFprk/DL
jkOgnVnOxLhX+fdYVRHJn7BETgp8YimFZSh16d597YMhsku3w4dp59/MDE3p3pa1
Gta9r99cun75LlI/uIiAOvuYvpMJabJq06mEkrmh4ewuNJfJ39b+yXYjW8vY/ADc
AeiXYuZvDQmUS08fVzsXIex7xEgLzgsxpvwt5Di2rIqM0Pwk42/GJ6DZqMNzpOI1
zvsghX5lxcUtizil2fycPYd/ba0H97BFVEem/B57znZjBwv6ByQV+iOPB0R71BnW
ibLOWcZALUIvbdo1OYd/gSVyhTwGJvOWmLsOfVVEAy8FjGeQx9/gKWy3+6bpbGN+
vlP5YXk9s3U83BJY8nw/FBc8FE2OT6YV5iav1IgPxEZR8uR2Dd0/ACSU+t/g6ZWe
0KjaDDgnaD6a079CmlSUhyqSdV3YEMaz5mOZVZey3BxEufWrZFtv+X9a0uXWSAYv
oCi7Y99iOkLwYP9Nkue2/FKN+Xjk+N2jfeRSuK/iW3ULnIb7cqWQZoNTnDMHYhvY
5MteB4vCHL9ybL5ks44eH0MEghSGgVJlYNNf+kmcDwzQs7wYT6GnDKd6cNKwAKWY
4EBFKqXpN+xJ9uKMGl49uDwiyUh0xzr87NYB3D0cgtdMJl1//WumF2tJKcO1i4ev
72bGhsXADP6PaCoHJA1ryLyNlOkA2RF+dclaXbQxQlhnbgIRo1ssc0cAD9Pt8Q5t
69+haoGCO1MkZIaI2M+GuR/LfcZCHTKIMXPIcWXL6E964McA0iJqdTY28ToAbb3L
+Q2tRX/gULW19tjBwQ0EU0T3GKiK6BkvatUQYk/zNMKi9xHISEcj/nZS4GJiZakq
OaKjDjq89EL7W0qY7VuUJGgCXaLbqyk3vOiwPYUFV4c9+VIvC9Av2aQ+OtIlfhbP
IZKYZnTag9muC7eLBnZTGhQcRSsOmJGdarc0jyntGnWbCAxt84ZvaGi/XXMh/LdS
TeIY8vqovCrNo5YX1nkPAdBI7LxV/PFuEfGiv9i7KyDXrGKZibg1mHAF3UyVctKn
fGXEiuOTxh3gpeCCBq0YUeRGvSkCqaQ7EvqsvDVrQR6FESgp62y+paqcmz/nF3/j
F3lgCxuAmzXofa5SuaNGP9dfqb8wCit8N72zfXLAUL7r3LVfJS/vn9iPPwK2zK7d
/CQVCdgtjtYmKIG6kbqyfEPStXR+33WHJFhpOZLNyLzACEVrrjP9z+rn9hrpUHFL
OnkUW8FBmIWhrSTr00ujXQexOHFx5XLmlr2CdK0QWf7Hqs9Zv57x5DYxwH+UaLCP
GvhlGpHImz97n0BXsittOWUnnYaGwgBfdduql/YHH65H6nQaPIlBZABlC09xL5DP
UsuLWU/6fCmR/2IhXRvdVxbg2/fVeLg6TPpgjb9uaUhhBXAbevxOpuPaEY8JG8qq
HFZbOSc23iTJJuoZjEnTG1ZaX3NfxiyHa1PBGz+kTK+vcFWC3GOAlEEB9iwCDuij
4wv+3nZOZuuC4TTLrkh/SkQ4gIr/fsWTMD5FlUOTHW7PAaLiU3K4oMmN8KjmTvXt
l7hyoGg5N95yqunm6D8IlxjtvdlZhwbj0wUcvvg/LE91iltatnpFgXYib9vhvFy4
uT6Lp6Kh+DYyAoqk+yTXAq6Clk6pn/hlGmTPpAUxi5W0cQX8X996mtGsQbNXkSnm
XEInYjZIe+XIEdh2qTlXT1XqdVqBggRfJBkZQiGSB8rjnB2zbjPO6fkWcnnx2xkJ
V4a3ILKm79oQKDIiKv+rWwk3/1jaULWHGVKXXl+EmTMqDJBf7aNwpCeBNRUkhHJ2
W/rWaHrAEzhvrfppUoppBuBVNY4bWvvW0N5ZyaFckYTGqjuUbvV5ovB2fyyCDZh9
4Z1yuXpMorJJR6NODwspwTMZKAxMqVG58ZLdCr7QiChg6WpL0w1c6D2m0rxmcEV0
dGiWIEpuQ8Blgpa0wv8WB16tO1S4cVHKaZKBCjLvLzYuHlzbglO6DOKIk947nGey
q1AHwOL0C6Na8IgoNn1ZSsZaKxwHP3OOvrGI6DMWZWq09vOO3il9ChPlVRZzzFyC
R67pqzigPCY0F6PO86Kblrt09fLwV4zhgOOwfutX74x9CQ3I2Q73yMIjOwU6F1Gt
uDjTLVXD14A+X1zDXVv7ZW5dd9i6C6Avh0ZpoRzQoqSjl2w0Xs2ABgBLRQBQCgir
H5G3+xshDs7UWGxv6EC4z48QlVYM5lL5Bq+NVH8TscemDwn5oo0EnAiIUtW3TB45
A7ms5qBu6DqcS9Dwx9j8Mcx+7fQDfGC94LSyTjz3YWsdEn56X4ZQvGEoUPnqY3OO
sl3Z1Uqu9mosNwcjjeSZDLQhZybrpYvbmrNR738AxdDmH0GgT5vetI2OQl9vAkcU
d+w9yLOMF2vUIuylrq/rEwjB5cilxdiATiPLC68es6LBNS97KWPsBBkGB6zQ9T0z
7ig2I760ts3evDA9h+Ba6LCGEEURuoaILdRlCw7lbcj4LgjbOlZl4/0QwVcW09+7
JsPJYWcwCn7WNAqt6fV2UPoUYn8e/AzutHunbHntl5rCWNsIMpYIuAKwxhtCNUg6
bsyhq0pOjczMmwbW8HIKULHB/62RHmFi6v06kzZPs3FUpSMG7fEcOmbSjVwSj/B4
+yuS3jwvnsYou5McvSVZL/A6YwGmG+WWDbYQTWZ3x4MhMCvPl0PrG7x+CsJ38CMA
2d/qGZ+/X3BBOReZ5kx86L74qzmuWU4+225iUIJdW7i6C96CUVfgNu/lhmwgDioj
8GV7TGrUi3YrOB2dqjuSYuwBjoIbDP1cP3Tjwa8ke4Y2u+Jk21lgISW98jgy9/rC
13lKsyQzayXV1b9PYQfSdtubXyASk6aGNiLrjkIB/oBTrxm/XISq1tDwO6RyvoPD
v2u7wcG/A7/D+zVQwF/41rHnOfgVN+htRVfXEfdJalx5pLyGqj2iUIkkU1EPyJg4
0ipYS7lsduJfSbye+QeQm4C9qa92cQOJgccaw6vn1LkGGyxOE2ASS0DOQUTOT78q
FH8zHfQhnZPeLGPz+FK02m7nzdLDKj4WpOQD4dl8v02eOJFd05yM40MBxllcy+hD
gBqJXMtTHTF78D55f+i9v5Ccvl8QT1qv+Q6YFSoUjBewnAkZAMFmPGg7ZM0+XM0w
B1G4j4im6OR8upj0jowTRzhiBIY0AI7/gIGq7EqZMFMDcJgebKnTNnXxO34vsrE/
g615kYzpqaLMKNiZQzSyAAXXqKBxnwU1p+NcSVBbjkWH1K0yovjhnw0kwCMoglv4
MYlBVYgjdpm7P2pacrTBBxrtl6HWP375LgGEOJdeTRdA1KH5JvTCm4VZdB2IAr+s
T3yBHLoACyD0ROA2tg1k0c9euMbXL2l6+pFsQ77D62PTc7IQLoSYqQaoOiTGL5xd
cQRQErzc77KH0CDTk5GtrmRywhAf+/78284gGjbVrgWNDH4NulbNnvRlxRO0WFwi
Wo2dDq2fmpY9LtYHW3plHShgBTE9ieY8zmFsTK/zJaT1dO7hB7S71OkE7HWKkcOE
R2/ohjFyGGDXMH6NMCOfwEFafx2mzLwSKh0cUUKQeEA3OWsMDOg7fqQ/dx4q1sv0
VqSglxtWyDZJTJd9E5fidgoNGPOp6YrO0NOe1EWjTxad6axAjXuZpyhG06ZcINR9
g7bCEtxQXnAO6W0Zy+tqqr0Ignj1zvjQzMqExwHpgm2HiF+QvBx8jwHRg5FSmGux
0XWdv2mg8y09JYQ1HwlB4AlXhRoUeQhPznL41Kyed525LxAZlalGYj1LlVTcvPYO
mErZSiZhl0ZgI3igt87lRfAyGYhZicQm8hShtotupNaOUGW+e3K1T0uLDm7Kz/9p
2vbmg618RIXIvC9uES5/NoQjY+HhWv0itUXfdaPhSaVYPwnIh8eNDdWbs3W66waj
U+nfoHekhIExko2SyZVX+9Xf1mSLJ5BylxKEmb8iQCaEKzn3a49MrBub4N325wZI
I/QSywMphUR8Mxb9t5151mB+YXGsQPYEoy4SBZH15fr8Hy7ijBLK+SIEyBn2anZn
Q7nWkhIonEOiVYzf7vBacVngRg1Inw88iIiKA9RyiK+LHFLg/B5IStJbbHZ44Yrk
/66fdxWqsU6/lfQHe6Z0/2Y3RNsqZIqhERu8oKzvoawNdGA9GCePWD3kxjTkWOKZ
MRswVoEE/jS3PtO2FkwCfUrTq+XEepWrdvuJHyMyMWVQakt08n2RF4oDm2RS0WF6
3SDOTbXFG6+jBYw8S0N7JexF8dMbSJjQdw9tNphUPi0kPNTsBNqesAa1/0+iVUOW
4bU2RBzJo/dDxTm1CtQkBKq0uTEvTVD4cvn3c9BgVWNN/X7r8Vwv+YnCGaJabT9b
NrxpC7GxZdAPcFg9PCmEPAp4O0UWO8wG+TC9WnKOrYNHZIvWVXAoHXqCwNBkbmWF
querUHEo8UO1sJSdF7sXdhX0ZlmifO55B1VUoW7mRGTb1C53Lpp+QmYQp825Qf/e
GpdeF/YChXSNcfy8BgpadWuomT8Ui72O6u24t+Xc6riqmHevmRJ9w+xNOFWuuwb2
wVQuYVHMF9D5hLP8X1aU9Yz8HwPy7nIz6QBqqUBDwtp6vOyymQl7kNxmUXyMtMmb
vLQQYv9t9HtpecHfyQVWtpdHiBiTStNkCZOJ35qZ4mkfM4y9CwYzBGlf+TkXauoH
NnyzX1J8oOPzGA81tEqxdVj1q2HUtzKhj6WwnfwgT7OEWOR3qYCs1y0x5kZdipgh
3QiFm4Ao1hK/J0NszHqVq7hcqG89kpw6x9oDH33Y5xNjIpCMr3SZyrrDFSqag/pU
lkq1xp7mD8XB2Q4x9WHqMmS0s4/J2ZWeiVXX8N5HK5cURRT0yfRhGC0dhs1OMilF
l5sBQY62tvTetdLojqdohT42UETk2WRvuLVu9kejDKgvqo54VOE6P2k8IwtwzE9r
mUkmLBnZWyLQ/EpMyQJgINMYZ1qaabOifz0umIpd7868MEyA9OfGbrhJ9YsDRb83
/Js6MuQXiiq/kiexnFgMwBUBqjtCtZ7PPc1SS8nhzHXRRP/uAoNYwMntUGycy8QI
P5rq6ZoX3V4y8dK8mYnmxTSfwGqVv0ht30gQnz3MCpRJRmAq0qAD7yYwJLZP8nxP
S5gt+nHzhFjfiQdTsJphWFcy7LCFUfHnI2kq3XPLUU+HBvVMnyLizbFHV/OVaQ2/
tvOw4mWVfOsC3aFupXth+bGuHs0ONBlt2J4g3nju1h5+Zi3DEy9TZB/D+9VfcyQv
ZfB9BRfmqPkbEGpXIRB2JU8uZPlrkjMpO4TCUOUjWRGV+N/911YeNQZq1At5y00P
BL0RTnlcs4dF3L00LKugs6tC0/UstgiO1EN2N28+cWSURC68glWvYKZBt54XRrdJ
xoLj05uTeeRqfS42n2fNikBq+xqZ6SE5GwWQULqSAxbzbMgc3eDeEcTenRPCUJKX
8oG0gBRlj3KRoBZWUKWZ2RUEjcNCpB+hxkqSbee2uusbhy0uD+0TFqKd7Dc9nxPQ
BB54MNtiVNltg1KlpJQ1OMEB/BrsP6Uw5Q/C2a74e9vN3T+6bpxLcsO8orZ/egyh
PiFXC0mZzFk/W/aMBxLTJnqKr5dYAwqvB20R88bMDAMCKxf+1IZbfX/gmZNYvvv7
hEitsUMg0fH56xSjMCUNv/72qBg59a2t3JmW+6aF4O7HQkL0AOiGDSayd0qucFlv
5dLrHE2NPcflMPssUuRnUzaV4GoRZv7rcFtW9JkpDgn4vAUi7vJV44Iw6BznIjBg
WFwwojPoCcoyZcPiw7ejEN7IOp9ocRJEyadpW9UYLWyAm/0elfaZvOboOtnWFAmG
LaD3y/+8Hfy7WT9+LwT/HxwPlOpce6+BizoV6SWvj0bbkxI7akJfQnup4yHRqlSa
55Dx5mP+R4P0on4Ph9vUuEnVVZtxvxM2I5nrfGd2RQd8bsWkvxRJXYAzjuCk8Gwz
Er4J9WpBGFu5dsRlDoqv6tDlBWRgE96JszO7Fk8it1eCOrizcTX7pIZszci3rvN5
nFgPFOsP25je4x/m8r10t1jR4YR84OHPzzEBCyDqpdLrsBHcs+43IRgXk+ST7n/J
2l9OJGpS6dMfzGm4Tbhc3nACVEjXA4+0jLMN7G6WND43f8YS5jXGgePpZHlP3wSG
6DtmhvQPQG2GsbMICEzugY+Pn6JOETikOxmE7d9/EtvD+DL9A0KvsBPeWpHvbly2
2Ws03yYIhgzEvGdFUiHe9HLvG6PKOmvlsIGEXwyQ8gkrTfXNru7EaBo4FLnQWaGL
ZASod1RQRhzFAx7k3KrY29tm4O4JJ901iIYO2Ls+dvYj8vn2dkxAwMUmsflHnfxc
2OmsTc6T3dA7eYeH/XZiz1gqKFiyIV7qB4Y1czM410Fi7E+c2fra0hVtYDATJ8Ki
DYmjM6CNWx2EfVBcZga+b+J8VkJ5Gh19rMf0FbBYTAHkJ0b/Bcw/npDvcPUbAtx8
2LNCWWis0nLKhb8/IGEQ4W9MFzqGvCyk1tKtZLEZ88hgCuAitYVVZolmGBEMUz7D
VG4uLriak6p2U2uq/B7ENKUEZYbeQts4CXDZL7q42qZTYlUuqjdAJiFqQc6pnE9H
tt3hVNSjSliGfJVq30eP0sMRKWS440OSrak5JhjIcp7nn8DibD8RK1LrKT/ol7Zd
3++ubS/5pXOZVR4AxiC5SWI/DnWUfs6tlpW99HR4SyLBdyEiLRyrORodam2gDGTU
NG9T6KXj7RVH7qZuFZUuWVSbWB6QQTP3p5Qedf3ZjWW+3RRPmTgOaaa0f29MxKXC
jTRlr+e9nH8/i8qY+RBAdk3uWSZZbmxeA8acSceAERimZ3J6SML57/1M5MuvcYuU
+sAkFXCRAgxNVfTLzWezBwOnwziRJ1QmLcfzqswWrKq+U4nOGa3XSx4ciM5KZ1Zl
m0fMPi5c/VrqXO81RAziaahZw8+Wj86C7TfbtMZ6Y61NLhyRupFFpcvJHBSUWDhw
Gu51MNrxf1oaTMEf7OBMRGNdMwUqjs7AbseELqQ6lOLxMid2srbm8qVIGfb1k8bR
+5aPOzLJUqWIK9lUkGtdGieVdI5nqMUJ4XgCEt7OlN/AF3a9vuI/6/QpR3oNvVWL
NhWSpYQFDOh96/kz+RAXXEaFd65N312/miIpCGn6coh+J3vM10/8ALBcSX8KecsN
QqrlaafuACxIyDl84W5XYe3w1p0w0YANm+TmsWY7botrodKQtoacQjUBMB+9vQ4O
2wzxnRWX6bB6EBNn3ptgy8YVDQ2kRBSV1HCgVo/alGh5mB26PocHHzD0iXPufRXp
yMAPMqazLbGZ5hWkt5QvWf0aouZyIwzVQPh4Npsoede8LOdrb11XwKjvFZe31Kyh
g38ZopobJWc0/PWFnV9jIBL/mz45ksSZRovGEe+Z6yx+FBO7ARFxes5MQ7852DsS
fa4CG3xl5SHG67ZRFFpYHaGYeYlUDFJ3vjo0O4BpCETvnW/eLNGl8yDW4bnIc5Yv
7b7l+X+m06nUXs3hb39QbW9iTFckJHQXnL0KGHPUXVGqrMilAbGegHXSxEOvjg5I
v203b3yZfT8fFniNUD4y+upyXOaXjPqzxTsvamubDx1WgfwBn0vH2ZGpcHB/jfo6
1hsNkeMi60RrOW6dCTRnkkcur02Ii/+eyI5MHnoIC3MEX4uG38BT60Vn4zZ0+UsE
r6I2/3zJNOEMJIJbfJ1nl4rXpVJOzJKsf69yfQAT52r+dDo/3IuOwVuANSWII/+U
xClUJrDtO0e2pNQwt//nvOfB8cRiPUMOT9eOpjNvZnXFE5egBvrb/Cj8JhA94IOL
oN/oc4kbk3T6NT+znGieqXqCp2vTphVm5l9AB7/w5hjHF8wp3K1bGHX3tcS0ruRP
o68DPRFp9umDkKm3ac4B9HZZ7iFqqfSWjakHuvl5W9erUrhHElSL0RLQT2xz4Cyw
UGPdiwgB2wU3RFbu8goK/qwlyh3DcYfG7AYKw9gtpFwqj/KenHkwdlWdSeBaehVh
lCWqsPysy+BhYMwleSSYENlAEpBDlac77DT2HX3oPnDTJdjzIoxfQtizvOWg2AtQ
pZ4JjhKUbNytg6z6xwWRF2W2bs0cInoj1O6LCbjdWqXi6kMiZKCs/WfkAhDr1j6q
6tKM7cak0FHPjgeKWbdaWiqYQEx9iKvxsCmx6p51eRHx+F+4379vaX7M85C2vzfZ
BlDXxz8UHnavpzl0IDyksGDk01j4R5KhCfdFWl/2Q8uhWZ5ujkD8z0/HxfuMfhMo
IjmxqKSX4ffIFrKh6M7WVgT8z2zM6AL584uqOXmVMboMeXzSZI4182FueC5EG/di
enu5S7ztm5EGwE+4DFp3nEgJnTTTS+i8Z0kY+oea5F6yDoSUzi+kU2b/anbtbt0Q
51WLYszYQWAMWx5jLkuLbkuxWt2dKTpZP2qHXb7Ba+VzMQqf2s6GZcO6vfXVSpRC
mtOiRkDKmAhX/YevvhP8Q4nVywZrsSWiyU5XGgMrln087IjuXsdTXN2mUnQ6gpAw
Zo4vujZ8IoU2nD2BasAMmkqXXOFxtmRtt8CzaVKWWyDAth+DcREUTq3M+BAneClG
ko1PmeL4nqexgGL1FrqG03tqa07wxYXUGEvuNw6GdtAbW0hCcDpI50SYntXtIdDr
q10kvJMDtDk+iU42NZytHCHTqFHHs+WHQVLG3HHGJzO8T0v/1rH2oZB8usPAp3SX
PELBOkMNw1fklFMb7l/+tJ66Q2agaZTZDtJSBeFl8r6/RPw4+aZQIrtiP4JL+hqL
NIPtUj9jcI0HbndWSpn8rlymByHJs/x6/nnCM3dgxwlUjvI1ZE7ehaA6EHRlg9kf
Kd12k7CnLxC0VhzAff4VU9zIt356KmAkiRDvmaU55nlqjm4OQRwYx9xIyg5nzYwH
si5zMtSXKh5h3U9X8Re8puQPXoQUkJ50CGK1G0tHQnk80SaCoQ6KaJ8AnOAOiSEd
vkng3rvqaN8TYg9w0TSzBywsFq7K7iYp5q1ypuREr52tyM00HoJezorm63fdScTM
F76Mqs3Na6ea4vXURrGZiK59/PBYwTfh5nVotRg3tk9E4H0vdYWKHJRoOPt8dYPF
kVA0EphzSxdqrsX0IUDXMuRH8pRGx2v4Z/1riFYMw++g34EfYz/blJFbMSMy+7AF
YK24xuFgH5TBybKYNaksb20uMsWIDPuI2Ij/Qr9OimZuTGrRlieBnU8xAFILTRAr
BEqtTa87Ht4oaXEVv9xJSptkPOiJU+E+WwwoA5yXxj8eeWiBg0b1CDhLyn7AQ+VI
I3MjtoBE78P6mOs4FPn32EaP+NIMfh09KU7vkEiudbaVNcnHWv9xLB8GkyrYqV2a
8n3c7ypIHU6MVtCQbBnBHfkjuHaZ1UgTCW1i+RzapXBRoGOuxoyDiS86K9a6SlIQ
iRao/ZQh40bOoeXXviK/OKgNtpdAsByEwYpF5utNBhxMXC+roPxprpVq/YexfP+w
xhfjN5qIk/k1+62xs+WIiiZfOZktiHUtDXru9zgVcj67PQ7llC34GiFEKg+ngQvU
19zzxQ0XLhpFC1vtimFhDD9w483mJL50iez3RYbwkBSxlHObKOhe12OoLXen4/f8
IQA8bA+t8EtLXyhJSY5Vh7KsypNghf8H84e8OgARddQhuLupbH5YPTAL1ciZdpa9
l5Or3rkIxF0rbIhzIBU/PuCn4C89QglS+hy2ouWXs425+cLtLtBZcdOtv9CeNzeG
VBQI/yLBVaexheMDmDxE7dGKVpooiXHGkaajcMqg5ObmTqDSh0fvIcg5qYhY7jK/
EGjhiP7VKna/G558Ptl005FiakAI76zqbq5o+/SdTbql8cDeXazJ8WKRTkX9ZVR5
goQqJiiyb9TZXi7lgu+wstI10pRCMzg4gVzJxlIMHyARtjAIndoUrcEU7FuWBfvA
qmC3qie0jb3iS/2wzBMS2MpxZ6n4L6fW06c+nHGeYUJXH6npf0s2+mzl6svmnw/g
JUDtKLjrwVTtdrL8AOj9GqYtOsbYiKQpv6VIiJ68KM2Xpqs+fHzoqhDTais2R0Hx
7vwlH2biP4iQSY+QT2ksUQ7r9Lin0nHnO9047LyDKcbGXL81P0B+0lZdt5oqJi6P
SKaIUqOlkAKhLVtv5X9JsTIb0mVQPpjHdmgIJn2quLU+EpThfixjfGG3JAAGVy41
a8/BCbQ5dfP5scZR4M9/aLWObf6D3EU+gkrhAjIeR7xOpZBQtVN7hcuDljWTDysx
ITk/L/mVuezXUHwpQ0AgnHy6uzTjeoa4xwELfShl1G8VxLZ3Xo6BhhxHu8GKrf4+
aNlndL64yO1GEXe77DjQcMINfRShTs5chQ++cGsEBosr1N8wlRcr5yL2PrnO3oCy
nPUiA03P4iyjS/R7+QFwZ7lCdFTPOz9w/oTx0IJ9n6sJbPL/HmM2EnIEyXfm+VAV
RywyjxdxLZQ7I9zMIpOnGPv64g9CbAY56AccdFnBPJU+anDvvygN/hY5XKIaa2ne
zTrMu2epakp+/dZli3TA9OPn9XRVG+2dbmPFE+wzSupv9ZsegKD0juyantaIF34A
ws0QJbeGyzn+xX09DoEP5mrjre22xwwIHEdbQ5Woy3vTVc3s4UtzijUOlOVq1jHk
YTYezejVnNoEB07mGyRVk7WLTMXGQ1uMZyt9aovpxBedr/ydr6weco8hsf6ebmBl
QqSODCnYwbz7kcRog++B5voKYW1XKwVQcYMotWt6B+/u5sGFafwGR3gu4ZZsA6jk
mbGXeSvPfHAMZ+OO6hDOY0g+0ITvtGySmZkid1y0o2n8S6Ihi/8EZlsW+Ra/9+Jd
svR7R2PHNYvhugb3CksQz8W5aCzmrSpyM+DTnxhhj6Qu8GGMD6uXtEvgJtkJ86j9
RgozUo4dYYditjCmotUEDWVqjz9ll+MaV2lyWMkQV/ZQpRlmbEmoj8nHl3F5e+pk
KcZcu2XVOKeqldAWLL3wUWzTcAiv3WbkM973gAgZMgeDPMPNjRzsidika++Z5VoU
uOt4GntjrVD129Ona699PLCGS6YoxnLNhUfRS2CqJdd+9sLY+FpwPXebMAOmcWfc
14pYZKEUR2qJCAJnvJMugT0w1cJ2ejT07CgdE3IZtfYhBNTEKOa7QGrrt/AS2r+N
XfD8xxSI2uD4IxtFPbFgHTr+6MxDh3aumRH6fQU6rC8ssJabs+gg7Q4+y9ivYh9j
somwHbZieHozFBkwtaCBfJ6VA/ki2HikQ2/GWWIugR57lPaiFBJmotCA+QVxuOm7
1vAKbPKNZgQBUgiuhwuhNdaz5IYDmbAKeuhRxk9ftqG6WQ6jopEk9DG1Oh/6BTnY
/QIKtvH6vs3yi3fzCLid1nSy7E2CF5Epey2Ip6gUfCw57iE7jqEXlisuXSZY6WAy
dQ7Jpic2Me2UYAoqktQfvEWgub+dJZsgFYJJMes1jSKTEwCBG9P4NaSzA0WOnjmI
o0TyKr6dL9Vwo1EDJ8QM5bgTRX1OEzzvFaaYHoEvsG1F22Zy8TVwNloihwXkIwr+
c8Z7mebhqc/QlBpXTc1ka2eXfLTqqlg1cy86wUQsdrGLXuCkgcA9xe7f1COcY4DC
ez6RAsIifqTCtggTau88XBQzM2r8vHrh8BDN1ZTvvM6OYO/mmjH5RjR1JOUU+N7j
Qgefa6yGAcP2XvGkolPLqXAtXOT0wcNe23iqdgsiaZqjPup4uKskheXiJ3qOgzNI
43syN4loYLQwqJTxuEX3wcY2ikynhJvVhSsUPq3dDGOtdz8vbNreB1kAwlr7UBTM
HZX1PzZpH5SFPAjZFKfUuoSbPn772KpAbQhwyl31OjxSzxeNQmkwRX4mIDI/BU4V
/x9KsExYX+bbc4oi/0PzqLfyBGQGNhCjIn1SgR1OClJofQ0c4cXENTvcmOdIMkPS
SzbR9gMk9D4W2uX8APVObQB4svadaRTYrjsXHlFn9ucELhVE7bLyQdmf4TkGADSc
52uVTvwqlshH3NfbWx5pUtQh7sg3pRzlOZ07Yj2qmaDrDJifFNDYviBGZQcK5XO4
UW1qCcxPqL40WovwZZR/Cp4glisCV/m6kzKaMbgAwS/GBZi6Apxd4x64cvdi0CpC
e6WjwWz/D8y0E7hFa+U3O+4g6UyncGLdGJQWDI6X9ytCcL05QTQhDvb75zqGvQSh
Mw79X8ut6ER/Xi7suiNMDoLm36Kq4L/GltfuCUo2OCdCBZoxGHioWUrrfeqxybih
4PNzDd3yB80AP/7u8KuFQg9lp4TYEsVgyiHhz4KB0wAOT3MYvSRnhMxcX/D1Xskz
PYoUeVlD0nZuIOuMQVwuc5C5dLqrW1doGQouaUhuI2X7SVImpxOG/MiNYg0Aqj2K
gnDlTu1ipcilXdO4jl8Nv3Vw6LpXc2CgoMdVjilFnIbfFIoTCm6IvCzE/oE+aEa9
JJO96H+oWMSUalhEGTeiZVNodl6tu761Q97FCzw0wL+a2+dDk3FJBbNv6zi3s8Vj
/qPs1bQbxRFv1fUbDEXbhJBcJ1ARQgMvtj2y3f0VchBs/U+YhLqHvY2ryIGP8buw
J20YdVSf5/1xWdEAMs+G8FsRmSciBNaVpuavbruUTvbNZAXj3oU+R6oakRx11b7Y
2YHA3nV9pOj4nEmJtXM8cxtCfE6khe0YHDWnztqQrbwkUvLVgxyTKrK45rqiPdeb
NCeuvXSoUKzNs16pOra2D9m9tPgpBQCTW0v3+ynKQH67hgDi8s2oKIjpZIzrsTkM
QQe3pt5441+/HI4v2q+EMuRpk7N+fyDhogfWT2rg9zqfndKPyZR2GLErTbm+DOyt
Tsg4/uXI37taiORgUvk/vegoEpDR/7W1EmtffX2MnvrSGE24xCKkbca12vnEoeMR
HYZlfsG3qYOF7YvB5yBT5JHhYx9GpE3VvNd9xgOnlf2Z9UU7SRinZ/B1AcpYUKSc
yjrC093eU0APqTU+CMewrG3GpXy6YdjPcRc1eL+kws9eg5USPkJG1szg7mKkGUli
SWG3yZPCLg/ik6Iz/U5AQsTUof1mpFNmTQ5Bdyd4BbPByWvtrD9cEmsTOJyqXppS
B12MI69Z5HNqYp86iFevKpEubbt7+aEFmnwiF5Q1budKVJvXspl4KDhHcSHfb+Xs
T/wCanAeMTnZ5ifDERXa67qAYelK7FTCTHwo5LzWe8bI42M+P+NlUhk9SB4XTU70
oUmTcInWonDwtLRlirTr2LmSmde1sC2IsGPikbvT6PB96Ul9aMOJhpv+nnGSJHU6
DQiKpFlLHtIT1DZCIr6M4qOTd9EXIMgGJ4hrZNjX/mRa56Vxb7desReVAiP9NNok
tAnwKD89AJqvp4GKHsZcKaduANNg93o/3fi1tQ7pBy0BQ5Ja9pQ26DvSio1eG98x
RvPPHbpOyAAHWn03X29HL8ARBXBZ1jP3w0a3OC12pwbLwKARJdkz78RG3y2jc0LA
czLmrOXRuL7MnNwDW1/i8DHc8IRMstorBae5JfCkFj9EafAXNVmYlZThCIjmUo3T
ywXUe2HpUSwr2GAa+O/vix9egMb0bKrgVkBJDt0bStibJ7GmqzBTAkopexqneo3J
3lBReFnQ7lSqUWVvX3QZlaxnhtwJaglCU7DI6Aj0+gfWlhp+8BKtaLqwt2nWXAa5
uhriYElIdPBIWsUtYgK1Uq4nYK6t3fDV1oG9oq5RjWkc6iZGbdnbhN8rd48Nizz+
W4hm+8057akg5gE/6N8dtfN2I+sC3OMFDd125N2MNu9MzrC/Q37fLe5AI2vBqojA
ImIWiuCfjc8XUYy/bmlvL+zFAJhZuIGfcRk5r5Yasudjgja7g7FR8472nxlbqqKJ
WZchjGXSpwYx6FzEKWbDqKF++cTFf+tYVqDWa0hzXPAdr2kZFcmy2DpSxPVijrsD
Yoak/dKNbbPW13f4W0WF7k5x4rzM1Zv7rdXi67fXJMHffxLBRlljyc17xd+n15ys
I9Gq02aO6bTzxeG7V5x2mE9s6SK2/D/x8CkYBx3UYKCdBscBXqrRAq64ePlhm8f2
58B5JowDPK5SAAm1D9hu4/MvVoKGBPRALCr/UB9k0PCjdheZiwYD+A9RdrP/e1nr
HWuMn2pnh3eYQP6g5+xd8OHfxPXzPalsyX0xq1dPOV+UocQH8SLouRKihqkYGZbD
FbbHgn4BiLhbTMkQ51/FuBJGEPKdH8XOBnwuQE2dmM2Vz+wGqEuLOjQAxLs2b+fq
SR1xzWq7tPBRCMF5LOYSjkALdfqjF/EO4RjAJshCc3Nt8V3yLqb72Vh9pAcXOn8p
qDiHPzQ/0wnsVblAP1kLOmFGRHGE/I+AtIxM9zjdJfS3FEQKBiABTfmBh9EDq6dZ
4dEygkIFVYie9jAVxxDI0lmbARqNgtvoWsBAq3Aj/BRCXybAtQ+R1wEn93dAndNa
q6xWXPYvxZhoiIMfZN1DBy8G/WLSR/lZGp7ikfIiyQ76LljZuQso9kqXLq/1+mN6
LqT27BwprIoyoFkaD/hXFVrGAiSMypOQJwAhuHIW8DMNwTA+C5FYdwWqzIyUmiFi
A0b3hR+HWPkS3+qyOs602Inoe0+4zyogKXRvhheJe29pBxjV/Fr/U6wUefGP6tka
zAcaZGf6SI9CCTNn+QkKUOvsGFH1sksh7Qc84C58k87pbWyLh8eqKWVVKnEjy78N
gRF3mmbKa8vtAI0FHDy6tyl0CVtOkbDtPbkvcFrBtChPRwkZ8QhoYPk4k5pMA1je
P5lyiaNXJr2DN+0jw7xZORWJ8hOXTdsixt+5fDDLYm6Td89jXp7NdYdCK9tUEefu
PaQBZi+Eu/ZfVTC1eMOst79WfC0Kq9c0x7yHFTFN3lzeG5af1bQmB4lvWuTPzQyq
Vm0CWCQQzaKpmb/Bl1Tn2usITgxjwul81DCknpOvsFur1nhysj5nJfVxXeaVvOwg
PpJhrkZVKd6fxOKYVqR528EVGpo+cFf1dmxY4fEYgz+LTEtriiwyhuXRI0LMEAbZ
9gKZrUqpU1LNF6ocXC41+FR8taItgNLHg5B+8Uhk2MNwl/g9Nud61rQ5wNz/TrQn
j3JSzl8p3GFzq/eRyvD2jnLiJ79LleKHhIxhZb+Zbr+u+GVpRJKVPCA4JEJ3I95r
rP6EyIXJXvP8+j1GHNty2rVONBR4dMEX8Th7ND116LoP8MSF9LsvbdC6HioOIdkS
voIXUEe9n2ly+XePWky/sHpyskd/DcT/EVs9/NrY/zW/9+ioUhHaLnZiz6IB4ivA
+06KF+Ocn/bLLJAmjZsglTuJYwAuhOjtYsdfWaWQodDcnCAjwEyMumLkfJDDTQ0f
vf1fBmvTkNK/dtT4r8uE0cI2iwMz5fHleRGLNmOkdWM7DeTdzkbADMwIe/wMadpC
XiNNpkBPLOLRwKVaKOdQ6+VjR1GrLwVjEQeCUQWiJPXsio/MAV8lIzSiLgcXv269
9+pwjaGLdZCqHnn6xZ+Pzs51R2w5BNFle+wK/vfCA8UAKr3ZkVLejywGI+Onw0iL
2mMhtnmagVjx5x9PDNnD2L8ZkbPhpY5Y+aF7AP3fLK0qLayiq2GfobO66zuJJuBp
TUQCTJqTi19WmSTQpcUv6gwvPtoMISpFIaeXdRWK9QrS/5FFmF8oobd/JPjNiwDu
mP6F7BtnOLHH23tT6MTFmyAL7CTyAzb3W8WgqXvW04C8+Rb20d68KvuCAp85Rzhy
Y6v4bmPzbeXLwgrEzL+nLtQt/gjCpBBMRIoOs7Z91rQB1PQTzGE56OqXcgGYEAcc
rH5V2BB2C9nlowS/HbK379UskDFTO+7BovgHC5tHdPbUjqPeWhh992bJIIIkL5eB
OZfSeZRpSHZTh5BqlCKKPdNw5SnvxNsW9IsaNxtkX2vAyLts8dMPYCeAAEq/oXml
wgxTKUHrw2JGvwLRtjrKD6sMJq7JgLSA19qRtu+p0CRb2SuVRVbaPCX9CpaHdQK4
NRoE7kTLbXJn6pHS338bUCmpOOJcqr3eT+E6JwAA/1mr/CsIHKONXgatTeMuk5Kv
gzlAD0OyF/I9GQvUq3FxLTMDi4NejSHdLU5UGWHhOlufXESh+VkG6vDiA20afnFi
ehMrRYqxAmqRtGplqEd1yv9e8L/U6TMg/YM133EcrVjf7cFgNnqVbd+Cg/OXcb6r
lnZcN4DYSeSziCpUlhO6bOCcOxp+laiOHB1VcQQsghycD4D5yWrvrNF5/fiK0iUg
ESaA9eh7NFoLZRxn2MRY9z1YvWOT/fIEI7QxEVAGg/lN/20/Uyny+XvC4CFvTkPf
OnlJojA5PoYOCj4gzKGTbZI1T4NvljE6vgbVBWqrJ3JMCUY58PMToCFEfxhEBtoF
0lKSU0QRX36MFhi7+CNVZgNrqu+kAPX2h8rCtI91UZKNh1ahGoji/bDoS6ckMt8m
OcurXHMQwS+uPpIRu7gPwfrlQ3QqWwEkSo7cCtRYy4k7IRXvYDfgiALo9ybfV7AH
qIYPJzx/QwRvEG1On5oX51ZmNRRRTm4e2Y66paTblEpq920DA44UsWnmnvimurYd
dP5dJYtbZOVvYBxduSZRr+p3iXQPq4b/kUw3cj00sP/NXmusUKjAUYWWeO2n7woe
l5bxrTi+t+D1r5v/jX41lLs6lSbIK2bi28aUxmiM6nC/0Jxy6rPCT8F6EbMlkPmJ
Ro2FVTfsJ1fhXmJ3jFLsCe/zBc4tp2PzVDYtYaXfq8/89cp3q/siYKVfat95dOZy
Cz9hcTxk/9QBl3DFxFc2ZCltuEFJLuh5Vdeq9b8W7defM8JswTJA5nugxDvHDkWz
FqOL+RgelgRIKOplHzQ90kx077dYrsd0ERCEAnUqxq3KYuqBS+OcrwK3dG8l0MCV
DOAkGtabpgYCXzsXOcQ+dtv4yhKq0FLI840WrXlQRGOvhXrhzFICpkolhTITBH1Y
VIGxG/XCwyhaztf+K/Mr+EbXcxN244jLl6orTpycROLL5FFiFjRAziI+Vm+zYiFP
9V4RXrtuWFR2DrpZoxvS4atdp0mj3+r/gjri36OLB3eRoRFkxVppMgrIRFB6KT3U
kjFkabj3xbVSJ8i2Vr3k7NjaW6KzQeLCK0Z5Nb/GtQZuTT2wbzf1ukbrN/Vm8fYA
caN26WspqNtnt0JxUgUf3z60siiYdaxvIsUX8mzQM+ZRRh5RwHuEZuaPoxKda8uw
W5iM9zX5eoXOlyBJ1eKZPbNRMq/D9dxmizB2NAWAzJmG3+bORVv+RHjpm8nY9cXJ
eugSFm8H0mfZBT+J1URecSoK7KCqpFbrsJRHe+2h0ntlV0/hmhq+LXdriahaHYNw
C1N69oCfpWj6L7baAQ39jcwViCsCFClEB/+I7HJ1gneGVr3WJe39yrkyJBas0aj8
cr6aUiqabZ8vrFutyizwZ4tjBKo/Yg1f2uVqYFj8PGiptoWZ+Fzm6bGVzYu06EEI
LhW4DqALjeJYJ8mKKlyIefuWT0JYGf1EBT3Z21JetXIiUuXuzUBuJBYgJuICrMEL
EBavQ1xzseAdHg00uRYNz7sMu1ciXwGVGF3309x/7p0P+5yhvCylwFX03RY6CioE
NTPvJWH/i+lvuRGBw502erZ1GYU+6szU9FZTxXY3g9ENMBGszJtkMJ1Rf1znKPRA
/tMMs4L1wiwptGvSPRv8/Km1g/g8VJ3gQmirJmKGYpm2vmTtENtJ4vWbdfdE4qc7
qNaEBR/RXFtljZNMgkormOnqHUz4MEJ3I/OB2Ig8D4g+nkMlGwHgTtTYBsEYviwB
v+a5/6pNHMpMYaKtnW9c+2lrC/ah95d799J0xyhHCU8UBVl0+YJLXMOFJYmM7gVF
DRucopK4vGlccqAGEhdYFSrepN8yZRCFq6Eh6BS3UbxLK9qCw1S1NNI+gnC2US5V
Q4ar+6wTjOK9j9BENt6pZKeEGYd7USNLDAFP2vq0OtuDw5ew/iN2C3lGnpUPTYFl
0GEJ8byvWmzbxMiO7RI986jcv8+FGoYM1WQkbNHHYxs2+XgDLjw/pGCD0405OJ2S
UkaPA6NT/cBRtb3XzBHD2valKtGIkcvTEMu0Gq+I8wO+4dBSXXwCQPPDHwf4jIse
hje7yljEmr8fTbB/xsBMpYktjs3/NGkGupdvfXd0amULH0pQTwu8ctePWfuejvHE
8kPp34GQHChen1M6R2ML6JTLpVEvw4ALbj/ihaoZsGEioKoGn6YCAW3ZiWkyUW5A
eOI+UMmVNvSpOiJUebmkP4WkBHR/iWVEFSfNLYJL9qNXXgaTHeaV7Y8OKu8d4/LP
dp4YmWHqhVEcF0Dp2ck3qgHVV2rcIqxioJm5gyK5/XljoABWVYera556fvFa9WVQ
8bNUdZ7uJOQqLVnYoOrKEb7wMPtmacK6/Ue4bFeoHRr+VU5JKZGN/0GiHhqYP3SG
/l65umSxBEKqY8hSRaZ7cHgcnjfAp6qgEprFhjvkMwfx0F5epvZqLJFMB94hsb37
PGSAYscEiminW1Cob94FLLJM/y7yYmn7dTDwlwY7E95KkWtEyic30zuxYfOBXLCU
a94bK8E4HTtO4xYpAbuUZ7vRlP/oZybWu3o4ORH2n8BE9zg1jRwu0xWSFETYEkKn
RaxP0Jfj0Gns3G7Qx+TkxEiRFvkV2k9PfW4Lp1orw92P8lRZmw2qy0owUtVOf7h2
+Zbjt/LddmKJTSzGTguRkP0jRxr1mjZOCmopg1iqB8qJBm48EUT94BlW0V+BnQMV
4nAT8I+jHBPHByg55lbyapHW2fGIlSjtTjTVHdis/nV8yyokG5K85qj4raYOhIad
0hJgsRdC5kFJ4HRIMuD1uDmxr5jwIcxdpY6hWAsxhyiBg/DDWnmmBLD8GF7WegLa
spkD/bkVydkF5tHFKkuvRhJDNGsJTFEqDurZv8ycD0+Td7/uVucgJ1KRamPouciv
tdVM/U6P6Vvu1sBWYTCiA5QQGdJNHmYYk6/ttqGZLKMfBmfcWD58XfDq3FYq8Fih
8fQYJSF8K9fv7HRV4ac2ijNvfVxAU87GwcZpy3B1Z5NdkC+PZH5WKo7MyIwymkAq
u9oq3Xy/OyAQwnKrNFsvC93xTH4kbFPZnIimneLavAARnBxk9DwVlUO5kdH1Tz8q
p6j3nw8jBWi8ige1FxBl9rxu8wg83q06K+Ev77l+Qdw+Q03ngvZVqRL88cQerRqV
1C80G1uM97zUBmxhE2GrfOsD3rvPknmkAy3otviOIuLGfVBEs0GwyE4Lc4IJaNRq
+Dp9J+ovj2loVBR3KIhbjwMDjjv4AzdDxXLiR5uobBsWMTy63S4e7sGkMyF3QQCs
nI8Y9Mg9sf9KrnsyXidOzZY84IPZxwP4trJp2Q1WNeE2nVwVskfheCUkek0+W7oa
yosqMUGg/bquOlV3XtTie5rWger4TfjeQHGTQf3YUjz9ZMvrvpNLKIZDNNiP78ow
QLo6DpWEjHYV1nKIDDoEMB15W8f2Mwp1CkkjXilhtZt75QFquVDMzzsuib41F4ET
r9qFpfycB7Rod6ERkCiJx190aTHmSr7dRk4MIeJOqOR33xUkhzuEXJh2IAdhgYG9
JdnXJLrXETfptMwZ0bzNHK0kRWaokNB3Dkt6IFByhwvR7SN9wSC+Edi8davxTkAt
9IBM6ACGdryxyHUh7KbpuBfOifxlQJYE0CON++Zh4vm0CUoBzcnL7ZcZL4YjY1EC
QWi2cbIuaqY9x88xIG9Ky6uYVskndEYKr2j6Z2ex+ZOAljS+6w5N4AGvO/u7FJBV
bq4WHA3OVgJGcOC1NGXK4Jr8PHh6apPiSPFGd5Pb9SzJQKF80ixlS0zFYz5Ddlyo
TIfQy9JUnoiTC950DWiiXvXL9CGO7NeASkh7torUsfsk9HnvgT2/RJoXqUTAWm3B
dN9n/QMiCEt9mhJMpmIbseU1vvBNT19CJBI23rICTOqj3aQMe7Oiq+9kU7Qkj7Jz
CWtLsWkoJZmmspxlJEYJL7RIGeDSuzRbvxJMqB6g1yiL/j02FG0OMQpcZui8aTs/
i/GWBkkhVL3kBQt5tmESK3i97J12ah6Jx70360XegmMmru+aYz3n0nQlIZqcEtOk
qYHhi43IkfoZWUocgw+R1wq2ZoyN9MamGthxN6UTlgkFQqx2BI+nOGxd66aOFEdv
YrhC9N71yARGGeHCkZOTQsF3ou6hm0Fso57ODSd5l0B2NlFuJqJ5+XVaAHEFNw4E
a6aQM0/aZnu3tqUQR5kT1KrhHN056zIbtRT3m5HBmUiiMbwPvidrzAN10HiHumVe
e6RNMIddKrBdbl4uNn8+ZpiUjBYcPlHx0KWkLa7QNcR/1zcUFUe6lKTX+lxA4s95
XEiLsegH9szcNC0XoZ1pdj5D3LDGfeT0HYzvgAolkj35tR9mC10GEmuotiblfVDA
v7wSeVbX5yejXoOwIjQ16LV30b2X3Yt+t++7PoJOwAr60Gfz+CnM0XSUxNn7ju0W
InAZgDPOHP54TI01izwRM1CShYw2yfhlJz6qNdhIt0dcntdtyxMM+iT0uD7Ej842
qSMxnCfMN7UNyYxLkasRW9wfkJWQvQmMMZUTkNmbCm1VHABeUwI9kmlybKofUhS3
XGYi8lhgJRvN6K6LFG/Mp3EOhXDOQJK6KxJCG/6F/EO+/HflnOaoemXG3lITu9ZN
TxzvBkmIEgIZPLIagW8LNA6+wI8iCrho5kNdwFvpQez/9rF3GeGXY9gBmeD/C7M7
kRpmKO4FdrCN8iGTqq1BRO/WEEtWf/DbMl6uelfbVbLD5W+ekf1ptm93uqnfgKbH
f/3rtrCfih1vVATZ/RBMIMDTSzdjE1AXAeAk92jKOfOed1npagkdQmhVxV1Wlu/E
SM8KiB2GJtvYIPmkwxfpyWRabRfZ66jVkK5sD1R4pd3Dmo1IW+vlrRv6XBaNu0NC
lohtLbHaMeW4mC48XtTdPvRl6273WtleIhRVKhkrPvDdWSilKFbEP5s0bVFpIfO7
eArn/pqjmPCa6pacpUxpEBxCR/t86SmeuZPDppq/1EbDuXVss6Y//KyEdp+kjQ/F
dS7K1MFwIJwPe1VBlWzupnPWvd4TVJhHy/j9jGYQYS1lAtcMASLY49RHKf5kGgDh
Go/Y35P1AcvVZxNTmCOy5IQsmCv1ojHVXNOfV4H4P1vpK8McwqMrnHiaC9o5G8x6
xctVT5mqL0gLB2z2bvU3tiwaEKIFnO6i9bQkGsSUGlDnxHDY8E/Qy8dXSOUP2vqe
00ytyFtJAn7lwtPf2/fAW3Ezk/q4YP4h/eu+V1q8SIL401AlYGkT0jE420v+0SU3
j/w74saHlfngk22qXvOTJ9WOLWTZrjbCgjZnhtxrwr4JQnxkQGgfDIBUypwpbOUG
oCqz+gJ7eEf15iiYNpEeY+Z/FwM/BfybYKKhMU7VXTEAJHNYv+wodT4ItN11i2B7
Yvv0hkSJ9AFJKIYjGzoAYGbQDB8nmebjvCgay4JuK8ccJcip9311xufHk8WDKzUF
7FBGJLa6ZABvL5PZGIpEpU5fBKfbr/e0VBEAUP+rH8F3VLMJHsIS18tfvG1WPOun
OMdDz6RkRbQOULpns1cDGypUv7jJPA3ZKesA13Z1z66XGYqfuleZtexbLE8Xbp1F
ywCb5yy61FdTmGb/x0cGhB01Ffu9xOKTyyHoZhijTxFBaLHjG+hRBWLHDKOWRVu3
4JhN/dQrd0a5qswHr9EVV4zhMdjrXVZU4hCmr0V8h7X1Q4NbhiKao2nJnL9qzkSH
PZl4G4Hs27/hajILo5R7qm7nR9w1mN+OlZUxB0SEXv/h4cjQjdnxzR0IDhhviykQ
4vvNWHKuA853J2gbkK1ssiDnzFYQO/M2JU/VGUUFNACwp0fZziKPsnTp5guOXNYn
I++sOyoVmkkhox30IYlCrlbAgpBoLFy3fXcM3W+7BYlFVGNuevm6G3zOzLHNG/TP
IHqK75GbgEIJ3BUViwUpGDG6Im+SzBEk6n0LMGLFoA/ANdMzVCHQqsZ2X9lhtgNB
R4XmGOETuQ9A2PHyY5zT5VNAac2mL0CHpl5xZ4Nj3IlI1CgY7BEjGl92wBFKrXc1
lgvTnHFcqygppK/ajnMrzaxLpz53+mV7srfR9wp1dalN0g+CaSEP59fJ99YuJxj1
s5/43SuiaenCjRWQQrbPJ5VOnMMJAtbrK4DP9ln7qfm7EJZxJ69JlogN0DPx235e
wJwy7mjAdjhpXe+GlLMoa/IDLvNH50tK2miotvA1Ddholc2kqH0G6lfmj3J5dHHt
Unu32AKSI71zWVnCIo501JDM7iCu4GrWXX0bWS+07TXDQd9ryq7RTTfxinqY1kR2
HCSt+Jzf1ywXpD3VJaYK2rcUrf/d880ZP3Mck0AC2LuPtwy3/BzLcuZR2lwXq/gT
+TRhw45lLTDg5aLCk2V4N9sVRIzl6DbTVHLIrzfMigCXEO5RZjsN209vD6V986tQ
nH8jkOeErLD3zzfQVpAM8j1he8KfnVE3XMjMuFZGTZkTUsaFOx71x8Yoqd1o9J2L
u9XSqeV8TUTj0eSL1sQsNwfLU5Umxe+46GgCBjUGCpqhknrDflAZE625WbcNrzYc
YXLWfTtC7PUxVcKpOdua4sQYkvvC7lYBDyOxpiTQJExATV21MmcBVzbaiF+JgQcX
9ogNXeLGzotkiQex5fURvlEyh4KTb7RdXaWFGXrSfN8+2nTEkbkOog+nYBTj4EZU
kU7hjIFwPaU9vklsqOKeahhoerVhX9PRCJxVCM5G1MznbV1R8Sa0YDT55HmOSIDN
LMTrEo5GdHeFMS54/4DCFd2Mls0JSennjZGbKEkfrKyr/hVQeaAbGGF+FYc+qgHf
lJFfx8oZ9akdCAdulxdzPwdvquaFqRw04KHTgTAFiIuL24eUXTr/QkzHIkyCVYiT
u0IsAMg2F/wdn0MzuQR5whvKGISrwFQBcd+v7zuWXoH73YZYSSeRDenSvO8/AvM6
d98pBp4d4gAX4qXGz0AoX28YWyWc6BrdBjGlh1DCClW2uqlQWq+YNPIWYf5ZiKIi
mFicjOQ9O7OWmgY6Cq5dh8ZARLwsQz+DjEz4TVas2GzJdh90/WyF2S1ruu9bkuH2
uygq+2Bi2GoN1EX3TIIOmRRm3/dmBUTrOGL87v13pDx0Nw1L9ijXK0XkO/fcJm+i
7aNDwTG4ucXv2X0aoabQ9fJIbIgnrXbrv3ynZQy9aF7LPN0XgUwy6OmnNMvRL/03
NGa0XEweszxNLfIvYknH2973oSbYNSzs1HeBaN4NtDEx18pk3PmLnJc+Ln5Fg7uo
mQZ8cJFyQuetIhLvs3rVY8WBpqpFrT6RVqvyUySUjNxm3K8E7j6QR0bTGsJFihV8
sJnDy2+GTpwhrc+6wqpeCLFs7Yl9COV85RBoJ4p9+gmAd+MGRPQNwb6CjQ3kxYJp
1CouYfUwiEXIEUeeXoDkD6G3hIqDcZmyCO0+2J098SpKtk79ub1Vl1qOADjYt0Yq
nK0rL8YMcpje/6STi45B3z6FCOjOc27jehmf7aL08tDz5UP6bPRzDBdxRS0LiHRn
1W86yibwLeUod6KlHwMXSByt+aiNXmAiV/i55AWH+8CbIqAp6ka6k/rgo481RJlF
Li9BMLX7ReuVnidAPEt0vv8Fe5iKDBBVghJYPhToTFEadvJ2bQo/fjn5zJ4AarDd
a4cdjxfUQ2rGLZs6Q/kPd2iMzYyF7LMUVFNEdDrXyfkkLizEiUE+CLsILIEA71iS
VQIzFUKv+GE44K0GNiK+m4wxRx/hLHFymydMMzKoRLQ8PfURDJPXPML/V8TavpFJ
ZVxZnqUmMOi9CCagHZfv+FfyE9ZzBKEgbG1kYoOi6dGJ3BeTyMIxYQHaIsywcJCk
7vsOyGM4FnNcE2FlFN66Ok4U+8+0IkWqx7L/fR3P6alfX48UfNoOXJztrj1JcXwZ
KZsCQc7QI03jJ2NUwxwUU4mxRNhqZz3UPvKVrFSW0oooE5KhIfAISD35mEZl7vs+
VUaBbBUOt2Y68Xw8ZIHBh+KNia8kYVWXsKvy3RBXEg+ZVqbuqVMk9sSgwnWmspn9
b1oLuNK/Q5ItcOuHIVHXJ4ny6WbwYczjeFd/g/0UvnHYtcMx2ZYR0XNVV9OJbTFe
eqIEG+HHOSNr4JoK86OZaFyudKQmfnIrWPqAyTayot3pAHoFDfyzGhxIHUiM/Yh2
59Gf1Yxt4Y6x14wtDkGy+hfF5AAYIpf8+rVDi6ZpiBLAxDoi0nhQwzUQdnuV+q6u
xX9UNC+weDH0sp7d8MhY7gCikz1N2evR05lVknfpKeWZaHJMbqk5EywNpRgt8NJx
khLjDPnYAC0nHZVSkEoVXPEvpGWPUfElMYHuPNI/tepSwy/5P4S+lkQDdbDhhg8r
/9pMlDdUMCqI8mJr/Lg4jD9gq6ft6+EM4ONuYgt/mb+UVTbouKUbIlh0cPAqFmim
EGWbyrI+MZZIYqcp/MPhs+UtGay3JBXyro5zxFShSFlSIc6hdCDFSTfPOxA9OYHW
/LA9kNuuIGiKZxqOTU3sDfVSQ3fvEwWcF/s5Kz+CLK/6WjNlNn2PE1GLBXyZABgm
+PfVTC6gITnNnbrNjIbnIy6saHQgTnypDwSpFYCHYl42QrtKfdrsnE5U2Wa4lJEu
QAkq9TllIsPKbdxWadnntB2p54bcG7A6HY/65YCfpNwMan4+BfAonS+CqslnxCsS
SD5cOHpVPYVNsN2XjqK/YP57yQlYz7S2S8klrdfIugW2jbgeR1v0PjRe8iFCOqBK
qeX3leahbEuv3gKQFwSTMtX+u8OZHCgTRTtmAOcDy4dbo43Bc6ZiIzNQdO9Ut9te
YMla5TTSn94+UJ5isZeDAlLB79+N2LqNu3TVim95F8j9goRY1bxKd+DaRp06OIm0
pOVTfGt0Xb7N43dthkrcjk/CN+Xsw6i10NCZXYJSsWaDw7MyX/ZnUUwnlG5eaYgB
V3OxV0kMxM8lC3tQn+znv5D3ibLtViCr6HV7dP3GP2iyWDS5+mXulCV3EphflqF/
/VbOvYnTknrWXHcxCZfynU4IOg7RcI2zgNKeiLq/8HgQN2Uu1AVNXuo+vvECq/Ga
V8tY9GH9QYYG3i/BLwSEw9Bi8uv7cijQxh6EIC32Fa0jRk/XY/6H7KMWxfcfUOtx
mi3bp5rgOJKNKUzdZobUl04YWbjNE99erhZ5+GSHpaNEU4ec7+6JZptyeeGYxXxt
AQYbJynkLjyDWlI+mJWPOtMw3DQYdintK7NCDTg81NND8KE49/XkZD5aWtParD5A
TQTIAxoaYSCleifrKyWZzYNpCqSif+Okw8sbpniALLJDSwTZkAM6c/URgtz7GM50
ig4vpiZMg27oT1gnaNXMxptYvLOC4+2xPrRWjjbUkyck/yNs4Rq0VQ/doL1Noi86
FUjmKMdSgC7rPk8AknfN3PgdjowWEzwsv9gTljE2QFR9GaQ70uIRnGR9S/jN64so
qJuRdjEeIaTUl7uy5LfJ/q+mtEVSJDqq5aAjkTJRuIVrqtca68BV1+mrKPCHONb2
703B3oYPTcH51tgw9MIyTMxLUP0ZJDEeEAtH5Ysk7PmweSS3aKcD4Wh64S1h6XjG
KHTDTvqqBlkQ0TIcPubwobk/dl5nhRRr8d35nP7n5wgp/7rCyyP+coZOefCcc4iA
RWFyaC7rRc4Ur4RzruPtc1m/AmZrxdPZ9i6dlnDL9D9fzlvZyCAVfg69lj46SAr4
NBIrAIl8rdBPrFOA+f5hCGoSNzwYtypM3WFEUAK6Nhfu9jGpqdwB/A5to2DEMTQt
2sv8E+DJG9AG12DSmyqJtciCD8ClcfkIevEqYVh2723lf8KFExFDYuKSrEWNPeaA
wAVBsqptGcMgdw53c6bMTJuzUfiIRsRuqoBUoT+QdvmHNwOht5O4FZ6nb5P2zsYg
lTj/K1z6b4JHboQCpAMBFRjz9zGxNPb1I2woqJrO9Ig3jLEtAhUv5k2E2m1oTYug
wErKzDHaenr07xtoYC/kEEVFijHMju5ZqfMvg+OB41KYpbuHlFCA9v3taaxwX7B0
Cyg/ofsB7yWYzA1uhgvrKWhipmrySoahFCRlPdnGzRyKUtgvVW3xWqpi55BVIpS1
v7Eu0e3AmnsR/9Vxoh/QiJh8+neFmsz/DSi1HWUKqGHbcfaHOwE8d8cuUkr4brnR
1RuBbn3jt1JGAZ0glAm8WlbPcbwGErgOtGGVsQnE8WttcwlPBps9LhIfsmheX4vw
czK0XUEnezt+ZqDe3vg4oBv4BYWSjN0PLwNFcjF0+LhnddYxUadVKKpZw9LZ/SuL
Eu1NcbSnInI2BwF9IjbtowUu5CyBHmK2PH7fh9jbnPNThMQOddjV0yrIZ9O8x40n
sKwtOqIrPVd3lkB38Rk83tVpg0Fv9raIYf9YXilrbi2qBMNbfUznyd1uoOkmNKcA
Xk0jm8/huNN/hKmGUk+2h7a+pWsNcX9KarCa/390ZiU67e5vE3Nk89XaDVtsQyn4
NOIuBWWYZNVfPxSCrUgvCNOSLiXtINlKnRSnz+Tlilg36+NOaimZcAd2lb21HD0X
Zwrs2eTXayPxOWUkmosSgNl4ore2csSfLW8/eN3l7eoyJK+roL1JFQad3LJKA25q
xALdsdI/mJI7dg1FfSD7N/xaAfABhIrukVbKQd8RQ9DIwUAfzM9AJg9MfQuPE4fd
1jem/TW086C240858cwd1F+/p4qt3bA7P4rvgb3Z/cXAeW11ry4JirpD7Bd5gYfC
O10/AkL2GCi7361GTzRxgR4XqrPLh21kjlJEAtyDcr1tyVTC5OBGY2Ihe8KyRDp5
cAfzs6IKn+41xy8lC/45+0qe4XZsgJYidVp9RGl2fpqSPdlOe+gxxHKKL65g1RC3
zhVMqyNlHrOZ+KEw8QK6ZdkzaAdmSdwhyYC7ym2V0S0S5DsLTUenptBBOHOpQZCD
XyjLx3r9UlBCSUjG9AbBA+iFZBTi6uhkTJWRcEXtJt9+JWF7+oxW8LkqVzArfEiS
jWOIexFd82Q9yySfzsmLAahKazA3rrWFmHJWdHssWwVOY0zjJX2dbZg5eo8B+cjc
YrTECy/+wM/fIIt0up2x5KHQATSQM4luL4IcrE7UI/AFqx4Z9fSXR+CPAbtBzM9W
OVcmWSVHnptJj5LppUG8T80CAe3IykEmqWagzfrqU8KAy7luCz4T9hVihywepRjz
+LWaTVd4Z1vXo7YrKyLmtZEKQzjfWK45FX99AJS5jEpfRDuXPg9lm5d3CLGuxkv4
D9CsNRmX11d7211rA3Rk6dg4pVJTSkC5l5ewXeseaFEmWyp5OVcYROEV1GkaNcK/
VVSjWx9oGafqmj5mNDXnMuXKScaRJjqLURC4fl2YOOIZqW50snnH0IY0L4h5i8c3
cEurY7axQsbJ3aLLKUyXgCNwWB1pOmx2mQYyNSpv69oFOvCjonpmDicYWc2uW7Jm
YWqwEYSx9tcayD3ddYaToTzmdFU0Qjq7TwxZVdaNBEb+TCII+ZrfhTrXvM1hObuK
KwzZq1g+atK6aBRaLaQYnbDz/ZGrXsTXktcfkxo0kBvP2IjUYPTwrd44vgkoGaga
kmpS8P95JJuPF6rkNQO8VdozTbx6L9h+LRj53HwrZkypYulfTtIfhjfYgvCDz/Aj
zBZe8eZdFb/BTzl7PuCDC/wx6MtHSGV2A7mW7ROkXLKof6S7QNvGCLzbnntGeKAP
564+umlPXArN/Bnqemr8xuXenh94xcN3HuJ6Nro2SXquYn+EnV2rhRuazLpw7bxv
+pT4qB//T/xquSefynQ4qDHLRoHRyxdw04+LNGSYrnXvXpPVOlS1HLnTf8ludYAK
QDBAW/EGZSbuwleqD4MvgK2plh/jDVXgu4zpfssqc/I8GXKPYOt0ZH5+qqCVDPkm
4Yeq8OUMCxVNAe3wXX/IxRL6bkOP/7B718s1zZnHeJ8BE+GPZoA+LEz2HT181E2I
k61hS349uaOdn/dnoGt3q0eay4drNV6OvZHpQUv1dgXmvPROwqRjdsBPpKnA8cSU
oF/awE2bJ4NwQPaI65Va21wYsobgC6I+3K4tUcwu9gOwMzL5KIXfMvGhlsk0IzAc
bjK5I6GdEj/aex0NZl9VvTRBKzvUSM1WOSGtffCB2gRu8zd1Airc3QyNEbHcPIM7
v/H/tizcvmoUhiIWOoF2dUmTqd2P0hBc0dgyDhqjlNaZ9Mn9zFC7Td6J+nYQfRmb
orBQG+a3oVbk9qPckfM80XPU+eybmApFgZzqdipYimp5sMOJuU1VPQbtaqTUbg+l
+dkVTcG1cilXYSfsux94XHX9H8wvr0bImcT31NMUre26fiyTwXvOo5YhZ8w0Q2SR
fO6rNxvxQWNAqlDz3U4o6M9SoluXcLKPDMhByDjuj2MdlF4MwWdz7hZBjvWJ+LXf
SCttjPhUeT4AH0XSfVnHXgYWTQBF3X7Rno3ypePYjZydPjEB976dJgSiK0YLeeyf
hRBGnzvnc3++Gyoif/VjKDqshKrtUYgyfPoRS9eLyFk9rL2NFFb/mztv4aL6UGGZ
YRzO0/wz1JhnFMym+8uWRDXh0lxVvp+G3lCFKobk4ww5bxPFIl398/+tUsW4znYB
WyMItpxh+8D5rDHQcZexflpFM/yM6C1DR8jhcunoy7V7Ushv5cWSLEyw/MmNAtYN
zPNoxq2QuJMcYIvkNs2WNej3vhmoExxqFLdcER8WjMQ66ql0mq1M00PZ2I7IGL0n
4yww6ImX9teUqmU09IOvhHuh22OxUBGXnnkiOQDlj95w8mR7DjKXvBRB2WfMyYWl
F7G2Smx6EmpP39Ls8xMk6IhDMfWW8iQWDf8aFZ8i+U4jfGHCmpFijTWHrLndin+A
ByOH92gGkkp5hoKdCEGKkuxKhkapY62YWYYQhTetsJ+tEsKgJrmvzGhR0qOpv19G
Wq9sTdrkzbobKCIn6PbfFkGoefj9/cqrp6uI+fpsHAc0EnK7BLaM+XJCnrALmcic
ENQxXA3OfxoMBEYVbyj//OtXWn+05/WwQ5b4/57F/OUUAIfMiF8xx05AwDrY90LP
sQFTCx202fJ5ihYkrjGnw9eCLywdPWHuSakRbF1Kftsj7Mn7lZIbx38f1U/oEt3I
NlkB5P78FcnywMUSg9GWOvsc53VinRD7pYR8nSwv8wF7PGil88x2TfvmL0GS8OZr
3jTXqAo3qmETBr72obCITkA4iwMb06ipzYztp8C21pjEEvZ2zJBpPqEejWOyQ7XZ
d9cjm2pKBi616VlS1ydOHKSGe54Z8eqwpNx20rjtrcHrgmRK23kgM2jR7w2Hx+M4
ffkdtOXCiHfcGhdcc44OBtektOzYqR25o/Nf/fVHs2LeHfrXPKJd8PRjvtO2MwGH
X3kMCFwEKJwfGjEJ25gWpeMr2XHA5OPquJSGUywQdUeFfxKn2aY3Cqh/fHhMYTrJ
oOXS/kwCbCk7B/HxU2UPAQliiwHn1OToY1LprZHazkP+5qz1JvdMFTDaijKVBKZX
Ys+S+eC7kFBnUyyGu+78gS0p/qpkCtLQRBehPJI0Y1j2OZ6ZCtMPHyW4idL6jki8
7jfUBTp61FlmuEnFQJkxOtSqls5ajqBT0CujDfDxU1xEMZYiQymfKQzGs6vhEspJ
uMia++b72j2QubgIoalavEtL07cBEBh/9mbqAgUT/bqfaCjRePqO+ohnhhCXCGHP
iVhLv1/7TqOC6pwx7bIr9fQ2BgxWETSreXUIxd6Dy+Br0MTRu7W6XGr+XcEXgkqH
jWcf1p8hhsu7TClNiF7yfIfw99oR2dwqghQVJ7PTRb7pfBnskn4nyXPWIAvEnK+6
jOCTrDYCC71L9Jr4LPdXttzWWUFOd34S02cWNfIXa60wkJoFAK6fsg6//s6h8WPb
Z78hqr6PruwANF5Am6gU8Gh/nbzXfNtgLv7EvnZHIMfo6da4DOjA+kr8DuSQGPR1
GRE8jCXTXpzxnuW3MrC4LqHU/+MAN4js4rn1zw1tMTK9uu8KG/hJm1akVZP68qXO
OyJA4q3TMPhgNaNCOObWOC7d6qQoO8urH50L94kUyhQ9X2EJAvmZ/GBfFT2byZEe
ENyd1rBRV2qgHPPE6z9tEPqWkZEKbS97b6dKU+2PhoO5fibDS5n0CyiiaLIc//ii
jf3f4VUFngT+X+R/fwqXoi2NRIYoO5+fC+D/nxqCSR1NPEkjcm18wq+d6XbXppYH
ucq5P3SLKNqHDwU00smfPwLI2laR5wWo1I9MrdM4UELfipeLPhhGZJ4+u1USNckb
jxCw+LQLRtr90xttGdrCz8hKVLHf705HAdocr0NXebqgeendMrXUTag0hXA44rko
GSynptEddx4D8Jrltcb6R/1bYD9rpEmumJlQRpAmGaqZ+cVVA36FhaIBR9qUGz/m
8m5uBqQ5rstIie4STxb0MWlOVue2JYUCSetKdOL63ccUVeKR7T+c5V6ytXjFviS/
UTsJ8pXuyXvrtD5zvJ8hs41kBFPJHBIzxhUO/SKdL2d5R96hsMrjf+IfWrQP54eu
A3s9NsUd2J5iMtEd4DlK4VCQLp+fb4THEGAWEpwVkEt3gSOPn2vF22dwNlfRPspW
/SulT1XV0/5qCZOe72FFNO9fPxeSF7rldA0qzET1Ao0gewxUDKMyBcGQl616/A2f
JgyUA70xT9VIac9Yfh8+So5ha7XeF/1t89oq+bDr7uLHf5t191CcrPakCOFpcNV/
1lzO4084JdMBRUrYwJyz4+gXVKyDz/Y04qFxf5irpmEF2J+r4pRLqNqBFzIDiGPx
7YhOYJbJ24cDm1jZCjXabN4n0p6PRcJlN7MUffHrtriO+n2vBAzsfVlFAkKCNB3Y
VfTBLAti+5MP9IVpSl1Jmyb0TeDPaOSzh+3jM2WIkpkcL8eHoIoufKZ3IEd6IIgy
IxoZ990mwXNLl7C/X/HZMRngawpgdKEx8vm/Bh30IvLf1W1nNKDU7XRbYSX3PtGr
awWfaOYbYE+vt+3OQZqZ7PXgW7fkv1+GKch+1Wv/2TlPPkJUklaEjv3aSJFquuD2
J1CDv4qyovfF8F1uwAJMxuB/xWEF3jfyRywfs7w0sLtmmwIvQLTk6CRwPYnYgCgL
eDndxyQ4sN4UNuUfYBhx7vCFeDd3bRI9cXyH7B7bG8vdzxDYy5E+0IaW9qf2CVPE
qtURpbgVAlwoY8qXca2xUOu2I0/EgiukBSybflInhYr/dlCIVsgF2u0GyqOnVuLY
JvrkCOajlobztn70APhjedneCUdlOCzZjLL0U4R1Pi9HFfnejcXndDRx3azjVOat
XifSg0mFqACPdhlENHHoyaOoZ+U0ei1ELjnbgC5gmRU+J25fUZCVsAYl1YVFVfTw
gbDax0x230ByvnJm3lFJ6bI0QG999DMaJPik/JcLhMImdKQLSdZ1qnU/3dTRHgJr
dfz2A7Ip9kCe4VCHCk0kjRw0+ROpYAGQad1KZuPGCQGmhQls6dd1d3weuXLLLK2s
UkyWjI5iS1XQrQFqXGPyp749JA/G1Qr9OfQWjaZBYDBsaPgh++ljfQDCTDbjze5c
2lZcBzFltezmxq5VxIJqVyOhQakaulxqV1uwaNCY9cW5XZyN9Dn568f0n5RBX1ec
xduLZyY28V66LOgQ8ejhINVWrGkNmG4QAQ/hQhb+tU00Xdvt0LkRwXcTFxHHJxYm
uPRl+PrlaxobnpOZWml2Fo0Yj3/Rw1mTXeFihOUJtcsU/sRpKcLUa6uTIZJ2fhMs
AfYgVRT7RUUVJOEa1YxeUFRGzuTJx+2IrqqT9VzOTQ2zE28nIx/CRowWrvSRGKwh
QvizRUrqDW/tHJRqgYrC8WTMS7jtpdc67bdkfLopRCAzkOCaSr6ekJQ5AoXHyv8E
fesWFBwTtv8wtdh2QvCAWHkO6dwWDFRh6Rc85VXcUHfAW5NN+zRVRAZO1dkhLjwu
NcpwWfGjiz5sp2/wSkDFT78Ae0RmTYGQW1ajKFsznTVRD6DZ+3RzBYReGMnHHwfk
era0ssj3+63JVdKt3KI43egB5rUDLU99AJq1Rtb1mmWXEsTWNK8iNTK+12GySJ9w
dWXqO7eWTMu//R4oTvOvwR8O1Iml91WBYkXGz2/1goJHuGzmog2+64edvIXqqVk8
AeWNFbdexWXUZruKKL/vOmViauUZBo6oCorvJdBXnfWQufjoUaMS51A0qIASJeSp
EYjVBpNzMEqOISVJd3FASkI8Q0DuUsBZIXTduw3GyylaV9JQCc0XeydhOXbEgXnM
DVVCVaAmEZCPwylVagVIecxKvzFe390yhWFP8Zowq+fqQTA/i+Gf1qgpH1qqcW0+
rtqte6MzD179Ct7hdA7Z+7BiYlq4PXNkvWr9qtKfAdLNZRu4iQx0hWJRGtqn2IqH
ViM5LbnCvjhf96YZLsq/5QP6XY5ySQG/2N4p7LZTwFqlQcqwawOyV/pfrgWUFBBY
KRNhn5NUyGZoyzQCZMveNpIT9H8TsLVQabClApGRaWVFjL3Si4pHKMY+931f3tdC
cbSkD6AroBG1jklQ52c9z0qXHLJiPhs0V5bjtvjE9d2Hr/LtsA0s1SD+hFZavsrY
1pr3lXtEPyE7ey+VWqMe63HG+MovblOhRPTZj/iO3LJ7fwujFbPE9Pyum6Kg7psf
Bn5Wcr19xxRerveJbdgTeKD8AGLyeEvqXhF5cQCJfUPK38S5Wr8Sz+NfLN99mjuT
FGPReqbLS5OTubXGtt+5MDD2f3yubTmjkyhLtxLAz0sOFVAsG9XZBpwkyMwLU88u
zFVfRK4/qTuVGWelraJSdM6tp7wGaux/5+9SrrW7sZ4KTZSqxMotb2mtPqnIg3tD
eKgvzWRLDvfi6bjCpM47w6HAhTuhxL0K946xWGhXW9BTYyQ9Go2d3ywaOz1iYC09
ajSfMnVqWanMWQeZVJMKYtJoctF+YX6CrRnNpgoai1JKMJes6oqQFpRahkJ5RTvo
oCRoXMScllzABukd/Ue6dX4GmwLBj1jREuyVDE0Ik/c/th56SxBeYjsZp/EHusSo
VJtbfWtUR/hyMCwsQ228fETRQqyrAt9lbPzbOspvPxACJnFOfPowizlxEUZOG/IP
3BZcWUkBiXtioUsCgFPow73zFdCCHjkX80yP4sOqpFWzIse9AgPT41e9JyX4rcEj
yQ/JHb6LIhLGSeYZIbtuym2i1Pd9DpLuAJL4r+HsCSoL5ppqmJenPf6lEnaekIBP
kAT3mrcRKrJ4I17285gde8dNcC+dd8mZ+mG1i8mzx5DIK3bWaXxhG61+LK1FnxkE
6SBR8fjioxOXvD57bc8ZyCNmy36XFI6dzWJ4hTeKXYBqxx2IolZ6m0OuftlKJEZ4
3w8G2AgZKABAXW5LUKPyvSlN7GsMqIxoo9HWFayusqbDOMoCu4xsEZrfq8FsN9MK
xreLfFH0b5G9DUtLGfhBuKIrIaEt19AVOUNAlSAu38Ub2Jq01CDsCTqQi1L8HG28
aojWyTP2UNlANMcGCixMPi8P79wmZXKdOkoovX6tYfhiiYfTmVbEjg8ZDYc73o7p
hFC4iP4FP9gAqpN5MZYYDihrhKhLSNPkYPy6wt5zQMYB77+OlN7KXUHxh1lrudMK
rwwnWbhnaW6nQi5nFDUt+YPRaQQyuSEFaD/slBPBpgEO/Wy+F1+ai6OdwhUi/JUd
Y2lyCaeVBVFYaYbJ0WDsqXNO37YE5vot7s6vW6QCrcSwPqYNxSveLjYasHsIVNG3
qY0+TIBveOZuTtpAJHKIPhm0INeLMUmkOCmdR3WYAlgI0cMHXCUpLBg9P/MC0NrO
8TPaRoyGtqnjifwV4EGBzF3ii7gzE07K0GZ1VrrVfAnN51ko9/qJZYvmqcBoyyNb
LI3n+houAE5jouUPnHQElpgg+BThJMDcl6MHU/SvVWef2sejgFbj+q5EK66TgPqN
ICPbo1xE9b3csLTP38i5PylWtMF+Fzn4HD37vCQqkKlnIYFfnjWMFny0iyiR9Cba
KQrFm2wfNDoKMpLQwZy/TkKKgX8bmnHXKqp1gw0biUd8CwpPTiCXtz3p3YTSyKCv
6XBaThIdcycckwo2034e7ygLs9pcYQzhQUtxy0pklUYFlbJ1ktEI6nnCroVIkDXC
wp43wgb+PgR5UeJR+jN1GKlPdRNIsT1nG0d+k44m9XI2W6+RpB0Notd7a1NIiQNq
K34KTpqaFUPRy7vio7cCD8bQ+1Un90XqfzMMpZwOBdSxRQg1yv4mpOjYc7saOjkG
v9buf0p5yOcuQKn1Uv20LQtYeNT90ncixTdThu9hpYHdux5YUgg0SWQFv81CmXAS
e1NneJm9AbuYY9OgIdihmWt7LreMDm3mnw0elb0MWwDnA1gVX20nu8SWtS1J+vZ5
7IrlUGZOI/SGtwJyw8ya1kdvBnCSfOXql5XAn6PDSe6P1vXKCT4q6RA4amCy+d/Q
HUKt0tIJHWqisw+qjD2MeZhEtqd2CsQL73KJIBznkOoRouzEPRfgddCv3c4SDJeF
D0mljmyP52RFiJcipF4Je/GrhTqU3jN4UWi0IUIp4ZKZHDc2aJuYgzPU6k3ciN4v
k+ogUc2hoAtZMX6Cr29kDXCsp8A+b5r2aLS63Y6rAnqnx+nm6YULVifb6jL9dUmk
Vzq1m7ULcR/shL+sbUcieJo8fbLkwO2hZvWHH5DIOEXq1FAzdfzBZo/iBWN0ShZ9
qKZv3RfRFWaO2XexbEXqKu44mJgENfkSiMd5Yy7M6Gf5dgclZpZuCmz2IaQ8Q1Y0
V+j0VRCU0FRU3l98wP+OvgBri4F2oqVun52EMO+zn5D0sAmBJF36F1ueYz00HB6P
7Lq4y+iwuFgn+1LybR+ARZC1D+QWlJSwRFW3ZuEukiHzd4BEWB4rxx9IIERaA9f8
mXGIiE7sY4y5N9l2NYNHZPrziEzjRi91faHo70PG09BTNdYpNIdgiuRFyfjvU8Ne
DauaPfFk4IIsSZD3Ijz6XxK0eN9eQdD20Dj8URDrBK8stxi/cNygIaPs1lyeKj5R
I0HXn4n+6JfV77Z2FpprfV9Eb0O2UksXOIIT/ms4KQCIEICkbLuqeeoH9DXWake2
Qn2hQpuR3+QxZ6+z5KNYq3WH26wxoo+I5FinFq6FKW3gfuK3WFGAgYfo5M/l9j4n
nCfN6g0NpTxw+5SNK5ZNHbo7nt9V0/ceKoXSuZw1IscGa0MxM8ilF3bc9TfLRl0g
OBYR/rRhNcD6aCVBAlYwNX/7jL+szpOhJVdxxOiBc1d+7whizl3jVWd/uTeTzUV7
qsJ8fu9SR0ZMNpAxs0tHQeVwYWuYM4RYCc5avqWiOdETPv9D++uia+ml9l+PsH8V
MskzLXs7goqGCwDegf26extVnitzw4y5yFftN5LgzRQV6Fyyb47fQjBMChreo5zH
oPAro/jcdM2D5fAnfPQKYzlaQTkLWT2cDvPtvrh7cxhF5+GlOcXZ/tLDFIdf53yD
4TF9qVLYpkPLGGeA41VWfkK62UYUGWb4NiQ8AN72MgP49KYHDVuUYsTClJg+xsbk
d8LshiUPIwf2vqOmpzFHVYNa/UCs71FMW3JnQnLT++MgPHCJlSRBtBSROgRAvq7J
FVNRAlDWWdTCJpcMfLJeSfWpyVn5rSMnlcZqwDjl1H9txOBH6teWBA4/9GZsCTCT
N+PiEGhG3ggvSLThdea7/1bBcg5wKJprAUN5DgSgbB/IGXSuCghrkzvOTeSCvc/9
p1zmzPQxAxJUZltwhVS3RjTMTMNkv/JotLmyEkTWJ1CcTTWGSUjDb/oNW1Z6ZD1D
hbtgWWXAfhslIAEfrGTKHZELic9/3MGDqUopIrA/U/+2Hs4qVbgrGzzBxDpoK4S2
rNLf6jDusEJP9sf425aMYgEjuHvPz68tQWPT/yys8+h3GeN9EzFwZqZXXpnBRSkM
aTwstCtrG76a8Tsfns8hbDsc4ZUgUCytooX+6L7wwGSZY9ZIrLZJWPiWcRFRptdM
XaAK0ZRuezKq4l8eSllqQ4UvnjowlNvbtRdY5D6UyifuYlUJw+ys+MFTk+JTcLQi
o4I8Mq4Ba72+0A4JtM8R7DjjHwsnliQs4FowPqaD6TcVpnXSr52LbxvbVwI3nrkW
U2J1IHluOCvJAHp/k2YCe8I/aysJzNXlg6BWTOgurgT21biGfDBfPKQ5nQnZ6XyX
Egh5PRcZ6lPHMDitZjJSdib49r0H+7YDHqEsaf0nhpm3VE7uiD/skSghuXQcoEUh
LXAGYJMGJ1cF64DnZqHLJ4ePVWfEvqMm65/oV42jZbRaqwh6XhO58hcF7+d5NQOC
MUMuVvXzpTEdQvWapcZ1+3496lxdXZdOU7MnYjqJLRtK+PHxbNzCqWyLA7B7KsGG
7AvlTiVt3RX0b5BoGsxX5LWeANiTLW3Yk0nAcq8CQSARpLNl0ZEtmDi7NtWIAy9y
cJK0BBxuWGNA2z4I+B3qWAXcfYCB3lgndr3349Ql98cEY0JubHe7Mu3FVYFdxIj/
fc+7LuyqTqsafMK/pBvfz8mPkVGSstUr5XqRvOMgECnoL6T4bs/nvkvQZCgnOWYm
L29BuJdou5WDMH7vpvb2OkYRkptY+vKMZv0cKMhD2cDlyqPLhQ9L6d9Sf01HnNsD
PufsATXNQcw8qWVD+xI45WJPgQjuWH6KCa/RiuiNlkCBrOMHiA4G3y/cB1GRprO7
6jLlt4mf6hAuakiXn0mQgigfkqmewArBXyomU6eqJ4rNcMWvhTOB3EnPa4Y02mVH
RIb+x3vGIuk660B9DCaiNmq76wZl/0u72repkM3gLy7s/JvPP4FaLfNgJZ1RFcdG
V9J0tNEpzmXSEb3OGzMRiE6OrgX4/7izlyyvdUsgx/xP9yo2k/vndL3bl4UTpCsN
sVjNrmLegFKVu+JuftZiwR5G5IOZPfegwQfhwP+89MWo4BZCLMyO5DRQnnSDx7wL
ycC6Y7CMnBAg84wCHwONIRfqbj7HKgjc+fVDzlNV/V/H6hrkZQuiw4SB0XcOfU3b
7mAP1O9skeNzpP+qZSwQMCenQGx03uepbTm51wG6eCYWXnIixRESbtfsVhli1jl7
vk0oedTB7GQvRffFxovyVN4pYND/6vnDAYlI8A6Mf+0AfQdQ39OnPxvaIlofZ+ol
Wk4bxhZ2EXVObas2P2lQhPRg3PNacDJ22xmgOppLuzf2xNCWczbcAjjGVk3WQ41h
JiVKdTIZG/MQpBlqvIeXoHuP7p8zFZtFzLsVJ0utBRbu1uh6Cq/eCrZSymFjvh+r
3qAgcCwGO07TfjOELi0AsVST5T+Fd9/GXzftagkzRfHieMggJRtqLX+oam9ZvMck
dOL8apcT8aGvR848YpzKOofCjoNlP6QEEw5S28lE6V/e0g8nZ+dse86fVpQ5+ama
RtYp8yV5+lKzrSSQTDjVFq/tWvfiO1UmD4B5HQWKtbNyfli1EjlsvG39ND928LKN
PRLAElhZb+oXLnWjnE5p3EKJrmjm7wfyFV4TejtuEPOJ/cjNuXng4xTqQUKxSYf7
lxXG1btyzUODvCxrMHByGIyLNEbVULNeuY1FXhATtKswAPwNrGTM4su5z7Hj5Nwe
UkljBMqyyfpNzNQDMWIkzjUASgRYeEbfjj/AANmLU7B5N6F/eAOFuhtaZ1UZRXiL
9OFDMZsyW2xHk8MjPQyjm4nKES8kI9ZcFsdmhnbOClDCgvEwPPQ98fKG18Wsc/Yv
LkhOvJd3VB2OnwjkS8fmRjKk5d4lmWUh1NYOtEALfadvjdiQ+o8NAudoJ09H4OXq
YmSCDUXbhatMj8Tym5Cyp6IYah+H20T5N7B7/wk0Zu8QW7l3HRKwtKJZejMulntj
Aer127IiyTn1hpBPQHI4hY+o8tEQbN8kyzC5ir81zNgzYPyUEtciPKBjA5p7KFBu
JeyCWwjoQHy9VcFZpjb7ANE+ryZJzro+UTLa00WKvwaNd+K8RPaMULelbsGp/Bm2
F5aktP9m8JbUyIlZ9IkkP/0XJiQsquIU+FpzmCU2WlPqCQnl7qbXR/nZx51xNfA8
rEF7Iy2AjJORTED/QjTPKNEy9bQVfwgR29caN2LWNfsIAH9tMvtrcSeXIMu6nCIX
Iojinf8xKSXtPUQ5Ozfmd6MEwZWpxfKJaB+ufhjJz3FOtEjnG4UGN9sxISGx1TCZ
06NjHX5sf6oYIuhPJ/mkpMStIvXsBTjxuQbtaPIIkosFUSE3HCh2vNsc/LefMHub
HGHfOhlVEIWbnhGiP9FjIZhQq/zdLk/chv5BRDortzEkkkoj1hDUYN26zMR071Js
JN2csG1cwigAVLfxceB3OAhPMgIusnLU0H+9WyJWmR+4g7QfBfCttRc0aa+UuwY7
fbwQuajh2E0LYmhJ08acaztOjmDkIEy8NhaTE72cl+/nNT6HVk7ZKbejAJdk3bWf
KDvQHcpFUZvsJUWgouzlzEMlvVicrukkUUayiMPY2g+zoMDrGCIMnOodvYW9MRrb
BVX/KEv1Rij/RpxUxz1QwGulj2L4/UKrLY9IxP7gRIj+H1tvfovJtuxe0NYD5OSh
XrKl/pHsCRQ6+lORWvVajzl4ZOeO5J9rn/w2Xi3cMwtx7KJ35eIbyba2tDdn4QX0
Qyzlv0LnpRK1p/KvAY4k2BMuANZ3lobxC3mIwXZuw6KXw2nfTQ7O03oY+jzz/E1v
O2cRtcmQSS+VbfN4oPSRbOaB7/kezds3wgmFDZTM4UJmQoF24XvFzrmk5ZgbVzep
MYKCtS3nfoWR0CSAcQnmA75669GaOhNUM1eeNy/mOvyJKqbRj8NMN8jzR4j2PCmJ
kOt+2SmNqEA2F7TD3HNZl1ymkIcJegrc7jj/VCclR6Kp7F/YpwIglzPGrd9E2eHS
nD/bT9uqcZA3Kn53ZX0u1bPIkA96OSDGLh1YTiMZIoKU9/QCoXfDh9eDKlkayOUj
eglzhqXS6aIFWktyikAEbkiKr7qGJUq7s35YI6KF9fnt+8kbeiLDhoemnn0u/Y1Z
BTvcIl2Te+Hmpe7cPyabsKZWoeaPPiEBDJX9wD3QBEPS8F5S9VCXeCvUfJcDLM86
WPO3aVNcvYznmA8Ulclk9OqIH2MCwZ2s2bNfz1IQCHtwt9qh1HSOQCauY/5HBxpL
xslkInbRr39NFRSvvfVVmmFVFD3Q1PDEi/BSUbuzcd3fPt4jabJgppYrh+rU1FA5
pb66LXo0xHxM2JEAgohNMASQOeyylHU8zwg+Hv0BZqHWoJz/hvp8gppQ/vbx9iDy
YODtoVyiXwFtajRKvMJ7hl0IdVIU789E9CRjmBoofBYrPRwM/LuPcKefLTe/TZQ1
cdxB29FUf1XVHHKY4/sfFckZvfjrq+UD0f7wWSlIakkW2QcWVCD5rbfNoiOtL8H0
Ul7b9mJMyA+Z+ZPP69SYLq9b/pJZXCg1XM/Jmmztb9yYc5YUuSIsgYST3cc1uwUS
mzpuB/OeeCF8z2XIECuhE/Qs89TLza5XCeQEE+SJalI0FdR7m2tBdhjuN/2xyMZh
8RjpU/rlDaK2nF8qh3isBcpUNOMMaLrcOXV25BWVkbAGEjWn73ElkVPxzkQ6/IvN
OSSfpx/AMsMLVidgBTKJHPHfNqn1B95FtLZkQXez4A3MK3Yg50LuNbLBoh+NTR+S
h6xk37kysmwzyV0jKvyurWHZF19ReI8KiRgXIN333cJ/QEVdy5Ztq6Ci1U1QiyqN
W2CY+aodx0oVZv3HjaXueqxU7YLGfXXTMcFtoiDt/8elukhXD4zFezFEuOeiKqeI
t+hO++4jQfWttERBNdakCbe0uiZL9LnvmaLNsTRhOr2rqs8EVqps5NZweWZB2UH9
7ozHt8p9Vl7Z7WemvyEwcug/y7eXRgdpSve+Y+fht7VvHGs+DXchyRQc9wRZQ06r
0avr5pxTS6KCRcZWcoam3s/k8WYF1wGRDIec0LPnv+3d8npQDrrG0ig63VEAOVqe
kiyUMaCh07yfXLD4YHiS5czRv0S5GdxCgkZcSllb5mJjTA7+hsTV6VJPCKvbYvO0
eLZ62ixU1itDkHRahgAjGuzKmtiuxc7uffbjLyiOcVUPS17ZSbF+31T2m1YIS3kV
1goZ4+3pQc1OjMVr++JbLGbd9jxjPsIL1BKFA6PSsTyOCg/8BX4b7ZtXlxaNpiKd
Yf4TsN7A47kW7abcsH1qlV88gnvaE1UWcF3lDxw2e+yZsIpc4ZU0vS1qGzLonTHP
GuTEbA3eavWzH7UYpgTd0r/54eOMDTOTe8HcXDFILVgnBfmrJQoW6JJryuUd3Ec3
9cBysAtwNZr1NNZRDcd/PBKfWuZhyi0CsMoromsFErDsh+s11Z40J6VOj4979GRT
MoyKn128DxWrmgDOA1nKTFqjzJ1jlTVAAszYAVxWPP5tH2VozEBDw12y/Js4+T8Q
k2ypJQr2ODWEeyCGQdFFqckSIX1eNdF3p6fxn9eUwOz4qZwySQ3+CzJ92Igv+acC
I7LqqyAjoei8CcCtcaAh6OLKGp9Q95++ei7oDWtt+KSjv6C8lxh3YmhmP/n0dObB
2JTVqTcgCH46JOpalgczQUDCcmnfEftfFkj7D82C6PbaYsRi6Oi65vHOOGQOtLPJ
N0QnIw5/Hm7YUsx/nRAWFFxU9+pKPrSIBsoMtk20G3XGdzQ946XzUc3n7x3yq9Q0
lRC5cFIx7oma9Go0MKonoTeJKkdRJuxVexRWEBKeBPnG8Ux8H4tVQGSZ65WrIgXK
L4qH98wQL5Nu+agUxxJ4VqGZ5tSvne65isls9SCX/NAl6x5nAvcpS+9aaM/92JbH
HdoqNMvkvSNWyhcGYMGcZ5f4DqgCNhwBslGBzloWfDyvbW3NZega2W04BQ72qhx4
Cx9mfyj1utv7m+yvp1S07AIIjnQdTRv5lMKv+FRRNMAz3QfKoDEdPjetbA5LM1F+
Mj7xhBG9tgdr7l2nbOa8y5Ec2y97M1t8MafyFwFgLMN+omzwTm8MkjVIQg6sqnjz
lh71Wne/nNxJ0jueNGPiylFYts3XLClV0smGtEa+yOQr6PapBH0XiRQpdkD8IOPs
CFCLMtfe6qG+GCNQ5NUDgWaXUoxabxLZEnY494QGZfrOjDqHqXSgdaO39ixGY0+y
1maVtOx03hy6RLGrJx1O3qwtOSX7FXji2qfYV1KFqxrnZJbiWIKob7FYGrGmFQud
F2oO4zrP9wq7ukVmBsk8e6XEqKpK02S+fBkt1b/zxmQ0Xq9RQXh6aQ5Hy6TY8Cf8
+drv8pJhg5ARcA03dXgqT5rZKZ+K8/vPYD8U4r9qWHHbOVgGzS1xxgTjTpfHXnC+
OuMFYjYOTE0CCElEjf0I16MQlwYTF3OW0FCitZaQbwjzyuVRgsY7v7wi4RQYQZ5C
tljPHIy/uvbV5ea+EqfPL+v9z73MtAjk0RKkft60frIupxXj5HfgzFXt1PLmRYD9
auK6N6tJqA7h9+BePLPwzdAEhaS+y5XdA7gGfowlxQtO1LK3NvBjygn/PiRI+fq8
+acfNZ8720XglkHVd82SKyIMWcRtcAVSMsy0VIZFXUnOt5T4iJXT6YLoTCKmaAVJ
cq2jcjX7XickTjVgL6MZfSx2g3DnzThOZdM35hKaxJMKA1d7cY8PtpHCCElYFO0b
36pdiGK9Ql8+Zdk7HEop1miuFH/Aw2lTV54F7Cb88bIU+5iC8owWNWW4KIabI8gA
KNQZy4gj5ZaB0ej3unkXXff0nNy14Ka3/YZqzZE0oAHHy2JztbjQ3Zvi5miX+TEP
+VtO7Yyz2502dYu7nNKLTTzbLpjWmPqavEE55744Rgef2/WY6q8kAcuOTQDQpozX
s5j9QFJD55uLZthyz0J0+XaWCKL4HuXCnKm4vvgefkT+Oi0QXTlSGO5x0Gz0f21B
mGvhUN15vcirYfvuA+zpobxAhe3phP190Jhr6Y3lrq4/BK8xLEoFFFFLHK7TDym/
5bAGsg6U+PVJlHbNmVqroqcf/aWZcc/gqfki3MlL7nqpVbR67pH1QUMXcg98FOzU
2k9DiJwQ4/75uXlaHujCCVN0eLnBHkvgDdaIupb3+/dXyLGb0AiXEHUgTtxz0Nh+
i9cv44SXvHg4QlzY+E7X9+JeABmunvtEb5qbJb7oLrlg6hZII+2J1b/Yt4NuzYKt
Ld6rzc+PcZz+pJvJXXVbpWJo1p/ClpgY2/TW5KXOY11itigVb0kN2MX21sjUyn8/
ZD5b4v9zegynj4Z6vga2Gj2rdWnMFLX2jo0yoioFIkBwWAaE5fq1Plic6pxBEDvj
+0s+rB6lKYUYS4XO1v2ExzISStnBV+lFvrXqRZFf0mTEh0+ymFPnEXJJct3VHOf7
Pwi3dTG9lE0uwALPL/bXhZPjwpp9XESB6jPhQle+ht4uGM6a3E6tlLR+rM2nkWCv
Q9dNljmdtiynFk1RSSOq56vG6KhZUwHnLbU4zg49YTffaVvv7cVA1AeUrXPzkFwl
PrBSerdoshLUUdEw2KdarrCV9wbukpHq9u7X1u3a8tEyYv2dhIxMzzbYuqBLVGDC
IBnO3VwZBS333t8+o4HlCcaC4Lb+oz1vfWphpvNWCNZ+1QqUNDB/IZwWlvHtIP2p
BVnkL6D1GGjfiraaJ02UDM7cLIxf0qGIUuG9nl/inhU08y1DgVSuc1xHo8GwIEUA
L2hS7ND/ImtZpirpZc2V9zMcdnJdPBI4Vn9Etto6loOeyfX9qMy2mPgB4milgCiK
hxf0g3EBQdwskz2lBt4CLg8NTAmACwyMNnHX/fdKg70CS/Ft1TYOxUesXWoKxIKo
oR0/+hp3voeKT/XgZgv4CbMACFqkS8LeOwpugE5lDsyxwjHt7EMolPiUcO0puupV
EN+ZRest3jWEH6fSUls7t5pT5VwkSIibDLImuGINJlSGRQZTscz9fbqdYqgi3bfq
9KUkhVeLroOXarDvg+JG4AkQJTMM8UsmkQ8YaFX8cnD0GoELpA49jBpKi7HbVcMU
g7Eqn9QXgqao0jC6TLMQ/z9BM9pnyfLvoIOesQhEgdNilKjY7QAA/iDp+v7JfbMp
J17HDpJQjDprAToI+2w3V6G9oQft4WV4sgdnjA064YcGtYzR76jdoZzYqlhW3PC3
/XjrEg3HRFtkdQH3Q75Znef5uXSjsv0p4s3SAPY9wJrATi2d1onoL2sqxTu7JYER
dPq9PAuB0ATDQwW0viBbnLqTzxhRarw3/meHRYt4RNP76QCt3C3t40nBS2qg/KYl
DOdS2MJbpXcI1rBlVffbMiBnhWNfndQVyD4xbuBLyT9cx1Om2xM08nPWus8K5rgn
+M3fn4dUc50K5oF3OpZFWu0taQ6XD08LJQMLqx3ufyViOr067M1udhMWta4cBfDJ
Ue4UKtZoWgoe0XrqoVEqPYZbcSpf+68XRjVh7zX/uV8/WggvCa0ysmMnXUe34Ge4
JRPjJTJb1kD96S5VSoIU5eCZY3swH8LyP2Mjs6r5kE2msEoVES56c1kF6WtY/n4Z
NyG2Sb/XMoq42D0Oy1dURihPBMWHz4Q+PB/SCYIl5svOIITTadf0/VsQ8imFCD6C
OzUbrj6OhBnVOc0WLlW+fmQpPWgd5WJcUG1V00eYWwE08Kd/XwXVpmMi7iYNqcGf
EAeNCA6QNPI15ITmw06BbJNF0LiLW4zkfKfWFlsu6NHqIZqBRfKVHsobufENpUSy
Hv4YMTXVhuH4dieBeViXEFtCGO80W6S1wfKFwHmGKqmvxK1CvUVFoR5UX3JQLXwn
Rr13DDRS8rvJBgzJscIbEaNzmoApAbsoY42joG+eQfy/3f1kvQPUDgD57OoZiLao
AXbHyDPckC42BfaRlp+9lE6EepGSZoUai4A6S1hVha2/+4UIMF3P+BflYHkV8Ndc
NICtTNrRdFuOOv6Y9n+SVzGWCgA5mnb8/dVvjBnt8X3XUM/4iFonyjK0Dy1VIh4U
68cD4zJIofeI/ZWsi3q/jYcE7cU5Rm+8gE6enuBtluRks9rQ8OX1A5uFuGVk1gOs
sCxg+RLgjN3oWksugOR6CfSClaNDdCaF0NoSS64mB2RN0E+lhbCQMo+GC9mEamKN
1Pjj+97ZA8bsi9V0ZjFQHpn8iBG3QWVT145IbiZqfu/z8yonJ4eDtzVvHLhbgcGP
7gs/cB/jOSjoMfNFSwuuNqkUWlkfX51aMdMflpUZwXdus7juE6sTmrGr409IMJQV
nagT4bajlJ00sxCAlr05SuIlyG39Ep973wUB5ojOvzx9bnDdg9m6nvxslQo6GXfO
eLs2hB7UOornWuBI0BocBWqRCXZM1f+Dfud5wlj8wqzFH6TpZvDRlshTsSOEPlYd
DswTdBf0aw42LS2eulMv1AaxKOx7u2sC266ns0blSswECHYU9BQm0tYM2JTNKrYm
VPRgIGx5i8btvjLAWUMW+MY4kAZ8DQxVd6lLHmGEkNgyiJTD69Pp7F5GeunE61es
9zeKWWLFOHf/GdvYdY++hOB9IklpRUNh+SK1aXPSkopx9y8sFX/QAl+qbICOGXtf
hYVTwt5NgoaTKZdj2Ar4gP0WkjktIe/EY9kaS+HqMLCrCFFRo7sFUQOlyHTAZE2J
j0rMcgbb11QtQMsQhqhqn7eCkASHUZap5bFMG3P7sCypcHWWmudpHyeaFpTCONoa
71T2x1+80ym5ZGPsu6tPiRpybDmLvmGgsUGNhDa4LO5AtAzWRUquLmR2PJWMpZKS
TPQWCl/S0W56rpr40FHknLr9fyD5qS6Ua57wTbxnGXKlCcZZT9swr0ENK1Nqpubi
DJxXEXWpaiPUbCs+Zb/nExdYYNlLdXafXtUG36uD+d+0G45aRYF8Hhg4Y1qWqW2E
szoaN4i8x05Fi1uNhV7NrDjHwZkqgf9IeRLr3Nj4jsBX28UzLhyz/2/cKMafm5pO
5cQqp2Wfko/J2E3e68f+aNdJdPqir+YXwlreninUi2raWi3mEtIZWLdiT6zlmzWQ
63d04Nci+xkDJzs5rDHD6y2nyFcKiuYFC2ypXdcK2J1sLewBL9+QBWzlXpf97zZM
UsaV+171IGSz6KLpIXbr1p77zhpfyrnLTTeua5Ptfq+TrMvq0BQJH9LEDiZ0/pLk
XdWDp4sNsgaD+8za2oqhLUPjlXZl65GqI1aWPSkV0EGHhiyQbdyxRG5vDCcQJz+0
dtbU4y8ZWVZTqwQVf9wCDqIdOpsYQAS4GJn+dD9Ez+KZJsIA/bgjGBl5vYokPg1u
7acYL7WVBNfBem/UgDHBi4yXckAWQweGSHDLfdTDSVUwmzVml8sdb5UTlgwumqGM
kp/it+zHZEN4q0jh6DQi7DechZov2mrjXaw3gDpjXBCSeLbf3JJMwLsp3f2gLHov
aG9FTWVDfUZ67UUhnUmxdw9FzsCQ+K1oCoHT9p9HAubN++50/w4m/otZp8zBO2Sv
riutppbgPuxS3e5wfPat6+XC0m3vEz5rRvXSO3xeaQkM6pOHyc+xnFJ2MSuPSre/
Ma69mGgaqBLvxhIxi8fiXCmiOhQpoi9Fdi8Ucc0YZ9hIIqReWoZ8dRXg4gtZeJUM
PixgqrYS1uugjNPNzFMhBJ5H++CMxYiGLAevKcbNFHd8L6HEGfQA3WHCQY+CuR4E
bnpN92sDkujkABXHQYQF8HaPIwOmFebLrfXC3ISYSGNZa+C2rvCVBnmjIShRDtJz
fG/xXjEPg12w1GfqVPbpCrSso4+Hb728+YWBOB0h7DHNIjlGkCUt18Dwr2gXSKEi
s/R8gKCVl8Ij7F4cljqTxMUFf85bOIjC1Qgi97Xe2PH9frgMytNto/uHCi0aVzVa
trghYN21W3MZ9aKYLu5msqcuppMI1nXb1VxdKXDcDFycz0nK/4eHPlPhPlQ0kEBY
U81VYte1LU5620EYANZj7VQOX5T2EeG2k5E8pkGeJZ8LopXtShNMsgzGy/jNbfMD
dRZ0IfdXRhjzObhTxJiJEvYSEAd1njADrlmGlSL+52bjJXrqOhowPP5p92nXkFBS
o0iJOblz0a2rtwuI5SE7dkOLLPQAQPeC6hkEpyGEw4qbuwHYVTaFUAoKYgpde/lg
HRySNyMMEAuwoWteG/vh9k9ekJb75QAOQNOqVzpjo1fjIMRcuYgVU42w0OulKbMs
sOemm9arlxOJjT7OYtqaXG1NqmRwZZTpukW+SUdz/elLjGPay4KkXuGZZJGRdN8G
XcbPIG6BBxKexlXGSwRJ7prYYqZJqTU2DAd+NYM5ibRm8dtAjgIze9K/aFYxuShZ
qPHL3KZiRpuDFI3YRNxirzepC/+lZeJkpzGoDH/SiMR2PyPW2Rox5EivsoTQATYY
3kDZYJWF5PPFoBcjvsNwuPVPxbvpBB5g/PzG+JWSL5X4yqDHZgL8oqOthRvUD1u3
14HcYd40TibeyYoXf89lvSpi+yQqrMmdCJNKdP19e1v5KUf/EbmIvJJInXkpb1D6
dzSGpHMvy3bLpuKyNg507h1LmTM4hGTKgvwmnZ4vbd1ZKE/28ds9AAboChxiowuk
Z8vl4gITAafP324eax2x+v6rGJ8qEE0AljWhZrA4p8Hud2l5b9XTuEfrt8Gd9ElL
NN/LMV5Gc+8rPZDahkzad1NxlOgt0CqXPPk4c/SLaklD9qUnfMuKwT4PBJXPzQEB
MY154Siwn58CbwUdVyZZ7/nCMDB6vJwsltIm/doHjeX8ftl8ZToZMQSHE6lGGt8q
GXSgj7pBGIvcBBFN/5/5BsTXgt3/yl09foBJ3vcDRDusZfXswTv3TTi37wi5oN/R
R8Pz5cR9GGVMJcgVV3N1HK2HEM1DTZw6wrX/gYOxU2laztKKTKm4GLR/hPEzEVx/
Tks9/wKnGUttuOd4ow0HFj2ZRQu27+Qmhn9mmganhMq29DGpRAkVRDf6TeujIQeb
OPUYKVHUOH3WgUobgvaPbgquVkP02d5ryFeU6zigtkjDN4dgGistQGiImPd2HZsc
hQKz4oDdYKyqod/0oMPyAAfKBkjzGD9UOKvdPcUZwZOqxqJIg7TL1A7tqQ6K/GdE
W6t+ICqTdOgXXX25zTGffb+ntxxA8PGjunUaKRoL5/09SjUvcMj2GLm4ipZmkQrK
qNjBrMAjMOGdNZWHxM3/Oe2/QhUjz9ehoT26CZ1oPj7DZC8a2HkXmLpQgUY5EfaF
7HJSESUXQol7JmT43ihV7gP2wyuj0M1tJHy7qWMHS5vKHduKtC7T5QM82aBoGJSI
nFzoyyok4xvhGxEZbnH5MqrcZw33N2M1G8wr+Z5lfgZw+SB4u0Os4N3Pa9RFAFoq
VKaQH0lGvlOJvfnHFGT+G3+dnpdWd/2EscuTKN9TTC4X/24EgLfFzR6/HuoxSQcG
AT/8/sVpyBhlevku+Mc6LgWBYsrVRpyglxQR8NyXmkGkL0/OlR6TMoCZ0Ojkt001
F+kjtUQ4Y0LihLWEdeQf4p9DHIWe6jJhHj/ST0QMboYBYRh8HONEzwuPKlycGehJ
feNfiw6r0K8m/rAKWNAh9JKMBjJ5lJAZRhzsHeX9a/uVsodA+Rn8s6HqXM41lJbV
Wnuw6948RA3Y/z80vnA6sighRyjkX3StV+3buSCE3cjxqjJDwPYA1jbAkxiyzw47
E/07lefUuy9Cu+1sgl/ht2anNu7O/oUDeaurqLWTPRodCDEZKhN6zLCfNt+usEBR
F+HEKdqlJj4RsBqTUkJj0tWE+qCKjm+KGq9s8ngoz0tyJZ2a2XerNEdcqZBfoGLm
GVR//RgCK6f3U4BYDLSP2eTzOsaRftgvKe1lr29p5PgrKEJicspCg5HcaJE9TiBp
XTz9DEoi/BHjZhfu7dgRmYyu2pnutHNJcHa4WI5ZVGmMDP62tGtbD+nrUzpZ/fgj
evfPuJCZhR2r8lNzor7ZUZgbeZLFyCAIAzhl/oau9s7cc5pTvHPn240f3XnvXhB5
o1GwrZlKnqvkLq3UnbB2EGXM5lOaQMJqkIguaCtymBGFh26x5Yei3tSk6Hf+z16V
ofsVk7J5d9ZkKciY3Y3JXiklJb/B8kMb4JaBZF1KCiGtVedIbIBHl9DogMupAj3w
YEKL6uUA1fuh00rmZOiaK8KE/wnoOxqWp/TuHtMuuAVlXhMgL8JfHqu6Izto37Qh
+2GCbxcQt2wsYBMVwGgvlohJUROhkDwhWPNATnvOTuo8zCTXNGcLD3EXNngyt2il
qRjj85QXcbeh2MPKgU+Mjbz66rm93np7sgD7aH79utYyJDpRljQ1UOuuMzCdjpjp
cn5L6nV1cv/DvqgiP5+SbVXHsunJSzslL8/TVKNkqxeaBZAMtWxwzksQoSmfi0/l
3uiuvJAXx52tvRjp9i4erc0YSOw6iR0Vs//SLztGwWrm+kWhoEmTEfzPn/evz53t
tVTzgWqKEIPit8OS3M0cxa7LU1GvtWlwF9kaaKfS7FHgCAdXzryyuGZ+GT816G0L
a3UOH0ZHQ5BIHgfyiaiHzzjwVXu+PxjwFM2w0C3WkOkVYsipz+J41rbfC1r+issR
azZSfELtYpgYvLU9jncBgdLLQOz4Gru3Y3Q+fYdDF1GnmHZ0N2KWM5yn8B7lXUE1
w97FROf5Sh5Iz14gPkdWPEUWSEVLEpikO47emPw3MuAaq93Oza4scEjfN/SY7JQi
TmUOnm863O2vCCFu/mEGBHgc1I5FGWtxGvwhwazgxjV/tIY6N1rCKI1MdNBe/XbZ
hka9UMSBli7eXrdQ5SeHd5uWJ9nZCZ5HHS/cTsuXwp0PO8vupzviqkzvvIDDLrTv
+Ma3G3lIPQzTKnW1Qxx4BX7p+V4yx9JfNhJ/Lc1ppqVvJV9mVMFCpGWac9tSSuW7
gGGWN3uhFJiWwYox1PxRSj9VlpuHxNztz80bH2D4w5FcMpdMLNyobxcnY8LQ8IvG
3Cbdn9c4gsucF9AnDJAI8qxG9deIeFDbsOzweNr/5rweT16QMCiEVUvPVm6nvAwx
TQ/WNaGk+bwK8xnNLutsjnVkHgyHUyTGZYxYQJKppshyB3GTSSeiFrZhnllwRyay
SuueO6whUXs/hfg6jra59WMVnP66If66Qh2LM42Q4nkmgV7/l6/QalI6eZogV6/E
McF1znjEHjjLUQQR2qegMZhDTaoZh7zzkujPFGUW2c1Og37q6bhYDyK2d2IP4KLY
lAxVQAObWB1Dmf/+HvEkPL/n6eOuJcUUSbMuUjqVaqNKSgB3VHeb9df/TzBvMUo4
zg4jvvmzgXVcRmMltHGu62jWMHpAijXDouB5twEjrjznd8y9czuS7gL2CMAb41pJ
PdnoGFeQj2FiHwgn0RlUpF5YXt2yO/LYv4u9wiiMaVuzkNOxYs6KB4LfJVP/kmLF
G716Z/Rt72/ywlkuEJYFmr+MA1CVWpAE9nFB3c/Ey6m7T+vYaUs9MSrnKL6xHV2L
Qha8DpZJmRiC1zNtWO69aXZVG9NW0NkUPYFfgd+oKb3zyh7TD+FMLbnFDoA5UaNj
xM3RP4lvzTXZm+suZIyl9VL1RGWRVeGgHrTisfbjatF6tmXL0ExsrMePHwJyWmZ/
MCX2oMWS9BpyFt5LztOfrUmz4Bg2Eo5b9f87XynpvqsUd/fyp1pFFABcEob+u8PE
0ohmF09YlWBUZMpbposDMD50mdzZgTxhBrHcOuNFlKpoOgPHmgqJ95IM4/rSsd0O
8+HAK/CbXhHrsLB5Eg3t+DqukBbYAwLtOA3FAK6l5EQyKUGlbrHgf7ZHDp9yXLw9
xbI5u3Qj6pLF38IY8w7cvhBc3xyV0irllExlPYQFV4StrerFXz6zZ7hKZGXTQm59
K9VGEr/FGt7gizPE6EI678FK3GV4JjCXa5EDa2NHODqnYIEyA+xA7418y9GLTZPa
K+vBDFASygHG0qxI6SoFcrS7/dkfqIfNF4Ye0wCHYCc20BhwUBbP0IH2fVQqGAkQ
21ALPhmp3X838z3WgXy6GAyKbW2zx0aYyPrVdkzfFrqz6ix9WSiJHRW46tUPW0Uh
ftzJSC/kNYS+lF0FdB2MEnxs8RwjMQYiKw9zpJKGAvopfoyvdja5aFvwSUwkKZtU
Y3GSojVdqoEX1cw6RTH6dw/npQQIIAMTv3XOOYUq2HVYoZE/3oQ81BQFsjT75lx0
hbmXg9o07wjMCSY8q0tqCfPPp2mS6gFVpCRk2+p7hat8NHs6AuIw5LpF7bu5Bkjf
ddSgFJ6bFKH8fo0LJJ5z//bOsjEr1osk1rTUzBdWOxzMSJOg9y7te9TQl8wglCPE
48VUxN2FZadlN8azlCO7wK9fd9hCcm6WIP2yjC9bDV4NBgd7bmehiE39+2+l91rq
H2uY9jHXy1xQ3V9y2HbvX4Nk+odAQ5986fQVt8ArijggbKrjnkQHuLLNxCdjN2iB
TMyCpvoQnbDkeLtXs37+Nht0j+ZId6sHQB9+3BHNpHyF0gFMMOzXxBlT4kDwxqzW
/wDAFw99yfo5t8N/MaWwbg5NkVh4pgkDY7d6b2Pf0M/upHCJRQcm67I+5XK+EK99
TLF0Jf1P2IqCfTRgOhO5zbjCSHZeVLF1gOurPvFdTBa5CCAmPeVG8iDvDqvAZyc4
wWjnxpsNT/WLVL5cGY3LUawxnfJ3YkmE9prvvQXRGuxyq4IV0X1ALSQ/OlWLTn3G
/qxZkWXfE0hQsKLud88/2p2NcNkU5kNCaPC3COyt2VME20smzrrYbhhNSUAT5/sw
iZ4I4PFyNgaW5JEiurrH7TcMtcajmNz3eyI5u2tq4CxTkTzEWSKbFMqLJjE37K5d
NbnpX4KpVuXeNv/A1K9kDjfyqPv/1714gDROo3Taj4tKOPEWRPVU9yPm9lOj+JTl
aRqfLVFPp3J17+cfnvugaQPDtOtpj6uYf1q1j0I1ITv2pGxNSrm/1MeifnLmOVYz
VDiqwzoMUgtWrtrY6sGEcLqbWeesbeXez5lHLrhbusLRoZO1F70XIP3fL3CASHvw
rK+eFWk8MC465Ti8aL3WR5PYGiecmCk0H7ffYVC83ztYrLdzQ590YVmalzUbIyUJ
3JTGRwNu4vuriLCXECAyZhVOaTPkVlRWjH5tTuvmvHINii2x+6S7dqOKapyykAL5
8K/VwSPyEPAMyEIqWDStFKzoJ5GpRoitfaDm4l3PuBlv0S3KhP93AthiXA3UX7nE
50hUqCpVycN+S5GC05mlvFyaigg773kQs8ccAZylUW+43z9lkY0oL/FgeA2udqT9
N37U++XbUNXLCql4kDcKyxwxLL/tkhIGuFhHYCEan7/G8naA3OVPjqyilifaCCf9
zruK/bP4VVX5QGlJ6rz8Siv6GDJiARMBB2jOuqeZJnNtftJJK/8GSHYEMjl5kQmc
DScyvudMouT1gnJUtQruFDqsC2BDYY+hHw4ETjLFdgLWdfoTArzuPNGZT3Qb2uIF
BcvMrRFz5DQHAL/r0qc3eg6pvo8ovpkmN7GL/eb8wbD+tThGwxAvRDPxLQ4ztTeE
HvXE5gGmHYNVZYU9IyVTXwa3ZRhBx4zSS6vAkHRsRFmgnxaaiPxVkHZa2+yLpmlX
wtfV3YeaKXgKygKKYPCuooWzin/AMWUkvBTzXT8/ehDJBq07iYmWkkZr0greEeKN
T5Fg6ZNKPpMhAKXvNQB6H451YRfEINZbgUG1zEaaojIDagdP9ztDJCle2n57AwLt
idFEZwq5WDEdFD+YHAJgLDOBEyaKUfTIIA4FlQ1FS3NKBaLVffpUZegSbgNScxMc
Z7vGLmNlxC5RlbEcN/jem7iIff9XcP8W15CMStmO1aSjCw7V4Xz2cmfZRnODfuBV
m7j9KeZ7xJk2i1RthJqXMSXrjg2H3uD5FArRGEs85vq4kG2zLr/sWp9dnSRAHKHF
gm8bk+oquN65A1//VuLk5l0utxdWK9bLe8nyk8CmJTNFLAwGUQcOp/DAG9n20MKm
sXfNicShbTGyNJp0OtRPuVW7oE2YWy2bZzF4WzCNZPC7MalSJcpmBagSG8j8ON1g
BFBSNshosXE17DFskGmW6R/i1ffLwc+mSQDlS8CbxTjk8gNoFnJqVXejPRWa8KSW
8v+SSDWfvKNn3Z9IBu+gezJGtvZ+nJzkSkDkyqbkytmBp+IcGDpo0S15IelEujIl
voA6D2RqfxgI0uWXQPP4YBo0/HUXh1c9hgwiCNqThnLVixqyzvXv0/gR3AWB6lKJ
H5d0/3u/zchQJMVgHGRsZjtj2w3gbmlYeEphXkHqjI2Xd/cReiSNKzLkEaFMWrgb
8xMvY0PA2l80gDiCSHKzIwHq2z22hFQxDZO/tCoF0TJSBp/twvIp1pOcZewowizZ
+DK7idJLyi+iNsFOBuBzXtmOXBY6Z3CvJftE7AXKBKXgYISUG/bnLsU/V68BLRCo
Fv+JYfNveqpc3WgYnQWjNaeNX8KN7JYeqOZxlvTe3G81ajUlNX41HHXzLrCCFmxd
mamy62Eayhuf6WzWzPL+35M5VIEL0uhuil3UKhaB9/K6lBIx2yLmIQesnVCS38nF
OopdVYIEoxQPgs8jKnJnhhCXPE909hiDp4kDZ9Q1bfMd3itmUOgo3QkcxgFkhujM
Vdm38Ax7sQwrtUOfwSiyoLYZ0G4VH1JraqvNjt5KpnFUWF/N8W99luUsOd3PRLVa
4+j8lQ+Kz6eYhgzKi7hgRHznaEWqf69KZh6V7if/GfyAEVS1nYU/4O5ar95YBAip
1kra8py1cYpVbcPvW1GSygA5TQlXlc2EBA/Va6ebE+YJ9N/2/k+0dSOe3drr6a70
M/LiIvSxctYhEl8xvd5Df3p+mmDWEth5bZdbGKMV9AzuqLaSUDv/nOr6xiM2/j2Z
xDMgTjC31skg+G0Z+gpcDcmsEn7NlU4k0Bg3W0Lo5CXhuyxfChhIchu2AuA8LED9
UA57OqDjPoD45PgQT0oAErTT8W+RH1oWQcyd5TtU2+fIY7NVXKXHQwH8bcahLFYD
GT2qD+rN6mrEnaVe5PJTmAwY53Isx3wMb+LYlgzbWO+gsnhKJHqQj3nju5annrwp
3ipl90y7B/XgK/AtYbPjlDd1IXvw55Cg3H3TfhI0iwRI8Obwbx6k5Km3t7ksUS7a
AhtB2YVUczC6Nj065p8avRvtsSAjawxPHK2g8TEmYLxYEOjrjCkjDbsYNZDju950
E+uVFLJSYiraWxlo9H5Z5VVUfXmgytqUCfy/B0PeDtG4puXMPQHV7w+iywXgNOAf
4qcJTCc7yJrhohiIEPSGBu0lXaEAFqybnvFE9JnDQlphsNlI1KvrCZ8+I2V5HswP
GLgTiBn0qRvZ7t6W9MkScrTRzN9f8nFp8GCR8yU5LCCaW7uVdsqT04Xo3STc5UCi
+6/dE8Bpx5loQyziD7ClM9gZ5QbQfLYgDRajNZEPsfkokcvZgpsCQUeYJrpR33bo
iZ6GrEwp4+0yXJBQacG0R9LPn8Og7YvVWcHfpg2QHc+B7NOS7GycdKtVnE3Vg75U
GMdm/+OXBLXr5yItz3FrcDOZsYzLWCaJik+Rnj6HootsB9b3F5+BZpiVfUTJhcgw
HYvgKAQ33foRbAZhhr5Oar3FlLqysQIA0mB9rG62/+y6E23X1HU4jj2RdzjKHGR4
Vb0gw9xcUd6hCa5enfMaUpr/8Z2akLR9ih7XSALMAhUYdBSSgilcNtoXyJHxrmhu
P+PJrhlmndZHKmlsERej54ajGFDzwOOu9RCM9iHca4HjtS3RNcl50LitSntYCTR9
Wa4DS5y+QUbXvCacUEno1mWIYHtEKoIs1nG25NxcKKOrUtUs239D9lymksUd7QMz
OJx9FwW0cyV4YD+csFH69JSgdKP/17Jjn++TjNAw7xmnvsp6kfcNHp+R3KfaAfD3
S3AM4fMUhCD5wW4grPthNIMjDx77twyGdPpTkE5c6RdhUv+//++2JMMffwlOptiY
+cGpZHXLlKvPZOwJjAsncN94Z5RIqolmgWVsIl4hqClS2iv57xy3HMF8sMhEnmx8
uJWXoZskVcZmLdnV6wpfFv7RPwrtk/phAJcpemFxVCv/V59f5hbT9anP5QkPj9Nv
Kd/VCgkJEYYm8XL3PD563BDfmXY5hJtjwJpKl73kfN8+ui5Y6hNb5QA3b/kes1Bh
o/CoK5daagSLeUrF3yepSSLC405ltauLviLfxzXMmpTL3IveR7uQSJrLhBxgz2iY
C/Vi/oQurEkix55rvttdud3EBmdCr7BjWbItdOiAozt/5cxqb9Fghpl07SdEWoF6
WK077vZFxI3coPj52TMEwqKbDwnSVSJCvENizSdWv8D9ssKHNKWsmEk5akt861pV
DJZqV3m+yD+TEuhLahpTsgjpliq8KqzGHS5Y0vnwSuSxFnIOLMtzRkZADuzLR1fB
naes+pkM0UdegshC7SibLSbjH6U/z89och5sVRdKFpWTTKsPrda9UzioennrxV0W
KQz2qY0uilM7zRMuL1gRR7+gx4PBQpzHsVe0IWulcOViEAb8JUWXDmCdM2bRAl6V
q12kLyKUGC43pWIPupdFOD1DDHWvQD5GAyEsAAxlSwn0WzEJJTsb3ljo5/p3pEmc
j3FOoPpwOAZH1OKeNQbzwzazCn0x3eZQFkeBdqb1fYqvC4oBarTkhfnz7N273GD9
q/EEpiLfQVCrOS8pOZsVkyjRfxMa6jhibJpKJKnL9Eql4NIsQ9/hc+2iVcHgVtf5
AY0xtCuaj3JlgTLkJveViLB/fQq9yMEULsCJCGzPcHxbgJQ+1kSUK5qDxd6AYqZ5
UHzRgc8A2kt4UtoEx0fly6bx46F6ZcVVUM73d7wTW+iHJn2UCJs/GThKmipT+F6+
S7xVwTON+SOv/GEUhqyS8qIjxouvWHgRljr6NGYCTN1/SD0D7RV5YJ5zw6WqVv7z
epDzpmRwVk2NH3jkxNLHo6hceGMvtuT6V+fF0GQ6WM3uRqxHoZC8H4iNgNQRNkLj
ZMevbMf+T4O+71RrQGJ8+CuIVtUug4Ejn51WRkTKNRjjS+bZX2wvbsch5cXcqoDL
6dVYf0vjCdfiQNJ246Da/bqQbxyUtbq3H+NQhwt9cPdggEuO4O91KWwpUqK0GKbr
fx+P2AwN3DRnTR/cbvlcdwWf7YvKrF+qX/JDOTLQEz+PuFb9afxqckWBAoYBIq8d
xxv/3WyaSPPmD2qHI0ulk9D8ip6sJUq44CjElMcsEqNuVsJABz7bg9EfFQvKSCwf
C+EQLvDmyBs02e+DCyIaSTzV9xfwEfGy7IalfPc/nvtXKwkJ6fkDXfXMp3dQNeVI
jk0f8f7RUHV+xS74Ggdc5R6+aN8cGLHaBE+Qhm+iJ8vIQ+MYmE1xXA++/3ReTboL
PEhzQVjyccTw6Glk7wpUL+y2Zt6dFgeViSKPysFgo3zaXEE4GBHFPb97lPqaQPbW
FyXmTTM42sRaBepfXmFwmYSLdJweVCHFM2T9TUmNW+PJr6hA5vHsrAguwhnURZsk
ydPhsfY0WkhZbDdpI/g/13MbqTx5KhdK/kGhywaZ43eCKDTnYAs31s5oIE6DJo9o
iyPDIxb1FVwjUWdgc+sKLUNUNn35ZFkEDn76GV5nye9qVW4MUoM5Ui32BwuqC/9E
XcRwXBy1VuwJap8tMdnytpqhtwrIq33urKjc9sLXo1LTJnQc52GRl3oOlM13MUV6
+sHwzbgSMdHF+kCpDCsmYpuT7inogK2o/fc+s94SojHu+nrkTDePUUKz1zB7kS75
oi1pq3zl2ZfAFlG/+SHj50ZjRYuhrszqIbOAcLwseHXvyC1Bbs8VLa/KzhhlWH9C
S7UJhm5isSss38h5d8CDXQokRfC24oXP1lgKq3N9DcyIbHJqWUp4gFue3vXYjfnE
FFNaLi5q1q8ixWPPdWIwczZS7+5bhPduK/9pNEHGqA/9AKEXOPSsSSjPaCMsGpf5
e0yo2QcTJ6hZ7sAwDvF3+PvjvVx2dayzzuA/heHap7F1tp5N4FxetuVXmYYvPT/A
NY++FnEIIJCBwhvhprrCN5Wp2X8kwAsVzd1E7wz+ahD6nVZTOjBWSqNbxLJrd2sJ
DdITLcQHxXN4vmrV82b7gvxishhvbHhQFP9HiJbWSuIcxvYuJkwtMKv6dKwLJdUq
1XIb95XqPsQNeh6bUc+/zyf7fTFt1a86b8HDM9V8WbEb8MUauPdltmWCTyj0w8hJ
zjqye6WeC4OMCHWuEkSLADUOTYhXDlcH7JHPP3tAMDJVNMdOqiHJcMImMnB+YSUb
2Co2takVPrqdzsTP/CMGY8IL0Paf18iRO2Wwzs63O7tK/SvG0HGO7hOFBYECr++7
e2WxYLRrgeo5K53ljctgGn+j9IeXHkV9glByfXQEM3ZfrcTQmiZBbHRK6PLtudZa
ZQhmaPnxsXM6NUaMPMGv6cI/pVx3Jw3iRNVYKPY59aV6Oyo6rdoUex1SGQRkL5rw
pzVGVyamFi1J/yJaixvKRpoFhhLU6WVNSLe66LSqoC8kAvxqi/LzZvMHqwh7BHQI
QcpE/JgkkGgRTvQoAQuRYbNrMoCJl+c3QP3ytsxyCYOoZTHoBS8vo8ChNB7OZ0Sj
DIGuReJqZDI/wzXCryZ2eR1UA7CvQWuA2Kj0CuMaxkoHBZdjgGSKQtm5ncrHJIMi
c3g24YQ8QKUqp5jAnh+kgPDsnBUGy9o+pa2hVHXrEkZsS0qbB18hBUO6y5PRkPXW
9zNpMurm5OI4Bzz6cfpFOyQH+oUAafVeHY7Ayi/2dnROUZgssMtBIcyLN8J/xqrz
CLtDCWcVkn2MDGh/18JGMw4cDI12M2/IlhC2WSVElFBUus5SLqVxEclqLm/lXhMX
r+Z8cAv1tqE9sl21YofYkbpbVxR7GuVsHOpWBTCNlpoR4dkjyFrX2VO8uSZkcjnN
+EDgLAV9ZGOVbFgO4dxSdB49TJHmr2s3TMeR5mXrKRtnyCBLhACgebb4zUX9u4ot
tdeD82yQu2njcZFlrNaSD2ex0HqEXrtqqXnuYrMhNKUSx3oaLrVCWdoFKH55zRpv
KjjV1qqNZrqGKA6nyaI1ufjGefzPz0ZdD+AZyN+KP/AJ+xGubrhAGcQLr/D3gqWW
8ST6Gmsv75mlzMhbT044KEApY7U1oAsM+9fBUjG8wedw0mIA6LPOrPf4G/+rMcoZ
DuAwKXc0VaN88AimGM5QdJQVvp6BwMxIHZiqdf+598dbaxHpFjwPZtHZuvZ/KUbJ
ZrYcOZZH9ASog0vSGJBZ1OrV0m7PDyx15dto9YWhI4yMrbFjJ/QHiv1d3P9B7ut2
FdqKeCnRWRgt3Ayc+gl//S1SSfP7ZjxjsL2zOoFvJSyq6h3Wh4hpN4Vo1FpY/uiD
LaM/bNv7t5RNjGZSz/MDVQ4v6H666NtvhpDe84Yc4GUjRYkEGYTAyZ+lvWfHx/vq
S7E2/wWzK0SOz1HeCLmIyrH72CiJpq7bXEQx2/RnPAAUg2GmARjIFLgXQ5xexU8b
bgfMB7igh6UcNd6LpCz+tVjJzEosGyBS6OMMvUmozYCbEFsN7peIvVm1hDW4smHZ
6mUNA6K2/YE7o0D9rF4pyOWnQrZLtK2EGtC8eMCIO7cnOmddn+BLGcXd0hPF7PzF
JxhrLuQS34HckT35abqGm4w3NoW+kkjF7/9a4fXieno/oYMDAfSKzZ+asiNnREKC
hhfV9B1xXePetqroBJhpw9O3huvsiCi8VDyIK69PEwdLhhTlH14kY6hWvvgD2399
vocl/9T78rBO7yLvZkY0FhIEpa/4Tx5TPLqZwxGYYL9qCNY9lqZyzBGO6YigJhW2
D5o65YJjGbEt+QxoqG2Jdd8IsAyBbArMt7E2sKIQCr57/iuHrqvrQa+eJOU4KVkD
GksV4roGTqhbxmHmidkzFG29SKyR8JN8jTQHtGlJdyiozdloe4R/U/Jqe1Htp4gr
AD62MmW2s+U/7ts3VVVFBU43NNmfcSkZjpwBlt3YOSpnoPYp0nKZryoYOqQLjlUC
6KWRcW+ut/E4oH4jj7HHgJ3WuMkTaINzozkwXeZ/NPgMGLPq1Q/QzVr9eXeYoZQk
WK7pHnMEvvvrM9anPHeMgo0MEel/k7YzxinQviEhbd9tlFkUGcpdjc/Jjf0qVLLW
nu463Pp1ZspDVrUeMhrsk8Ior727HVU0z5WkNAcCb2TQ+Vd4U69zfhroiB3EJ9gI
c5oocADeyzgOI+4WYyFCphJIiiT4r/zAdPGKFBAbovAy4Ogij6XB4AIKauv9kB7m
DBUQXzFsQa1iDaNfiF2oCOJFTdNWUqk/BuM6axiR4pFOsoPAYlyIH5tfNB9fjvBq
cbMj+/WTNS/n44/YuuvWiMIeO87uc39RRcaf/jQ2aycQboJGw9Q3QUFaemhPFHJl
DdgcDaFf9ryfklUQ0UO+Zj3PkFOs8/mLjI8CDTaetM48ZauzgEefJ9uTC1e4R+6g
lqYWNPN4QgkCwdfhhIR4+J/08/BnvHnCmHqq0dhkSQgIgjLNDbrt/aZNJr4KOgY6
oLgsJ2xdPKNOFq11Bo8DZQvOSJE3ZtBOp3eu1XB41pkel2iC9uBLU4Ot/wRA6PJP
woHVx/pCJdta6UjUlm6bWAgO1GQGyByDivfnnV2BqMJWWC53X68BlLVBElntJQ0k
Ung3ZU117dZy/z9EG0WG8jOHyYfRZ4twTb2IgZc22uWY4eaNie216G5NJyuVNVnB
hWQblAPBTcCiRe7ChRxGqQtTO3wuDprDHJPHP5aPJvEiov6NpwcT9by4z2KMynTg
vyDw0tcwfI/fLUHsVDsRP8XAF/hntESSG2V99plqebgbslDt+BnEybecA//75Wd/
pKdVEM+pJn3euYpakAUvRXiFSZY7Ya9RfY/K24EaVbavR4k02ZPhnjMLl7yRCu5N
0ASniK6Upa0imcA7gcVVB6xp3fx5v4g2Dsb5XN1kWng707FqW1dcjMEY+ZNIOFm9
7XS39rSdXGvGW8A25HrBHhiBWAMLhFIfWQyYQO1CfDMeafXBdGtUeKSTtCgL0q0k
nyKltFTNtQy02zlKXBksAbmxYWFlHt5Q7fZ2Y9KkOwKdg3Nw7oh4FwO3RrdJoheK
mJSWXtCTnCojYVaUHTnXO2t38lKxSG3j2yMVKC6bmilDsOQh+USlubluNmaDJ7Ql
HAKevOy9ZiqHWDImNfirlA05ORYGWDPrbC9n+bW4FzsQWptuUqBwjXzgp1+/pK7g
5YBVNUBv9aSzpL99zJBvmDOFyctJvF8hag4zvG/FD/KsIncRLiCsSR0ZA0FCmdC9
iGzn4zal1X4e+9tMI/8ksEhuQZq9r4fhkHkim8wfqeZvXmWzUqdYXluj6i8C1gPP
vAkmfIZVf/lBaBdEzJT5iKMiYu4hk1Gx5r7kgQ/x8g2EO2FoW0+CPc37UZwH9NEV
OAm6McOOcafJ7Neqo/ZXeS/Hw7CIfdJOrZMBHGwpqpAIEbncAAkUcEyH0Fhm1SAV
hOoPwJa0asLLsMDeOJN6R4og1Ug08KovZp+l6t2OWIsN5KgFq77LR1yLAz8TO+wf
ynvujktl4i9tCnxLQR92uZwFhoGLsRaMqz4tXR6veg5Nm1eiFfHhXit44cgDR4H6
+WrOfJaw6X0pH3sVFs/8PLq1yScFzRUlkxeRc04BG9xFM3YEu0s7eG70Zscs69yA
2zjvIyGX+w+hMqC2zv2w3ll+vRZOTexC022ZX6+yQOySeNf1X/tRtTcnE5mbrwIF
NGSmANixz0lE3nt/Oy24buXv0EhDSPFU6nacJzg6rvhrexeQW7oyJ+IfjBaEIRwM
ETI6ZkvMoCf/y44OYZyu5ziZtu5iK9ML1WIrsBuPYV4YTyTU0KK87lE8tDphV08J
T2nhCvA3ntt2XjHm2D8xsq0iFz7ugMDi+KJfpd7KZvJ/OLls8z/YabFQcFs8Jmpi
C9zdxfNfs1wQ+nME63AsEiROkDHnNgRYhBXHHV5YS92dsQ9i/43a9aOLCt9+qNvl
8QDx84QeG1P71v46fBoWOcZ0fZSn6T5ax1iNuBZ0fKN27Zi7UgIUdSQN72dGYESR
nYgD3pVKmw5FkO/Q7s7f9tvWbmKwdPVlBrerOvQvNlxN0ZBc0QG2JNaIakZAbyBh
zSXGDwFnnMIJgzY2I0bmsUjC7CUxPBeQP8mHik61/XyWDVhPPAAcNNO0yyzAAl9A
bri+jOf6EyCkpzvJlxb3c+auXltq5HedDJbo6BSEMfs23A00eGf7saunMHE7uySP
TmExJ1oNR4EXN0fvvWbO5Ne9AfaWlpaXShI6wgIJQ23p0MW9wTesj4dG+s6rAQ+b
C0DizlizmQxHvDU0qvVgntP9Ul22gIzJcIfVVvkolUUVJEWi6QlE9gTinvoa9EHY
vqof6yyTZHfWicgG/yWpC/w7lISi6k1YadA8g+celp8A5SMygKUalodTWDqHjYE2
qe6er/GnHZl3yzojFni7y13VNImPrlf9r5d25J0dLexMQDUXKrZXLR8BFPkcxgQb
lpCPV40IxEA+Yf9bHpx48ho3d+6Wdwsct8DHgoLkLuCmqQzx0O984+WBo+8vLETC
jkctPsXlDhmHFXt1RovezwRJagS3QOtPyDLLtqgrACERPi3v+f5p+ki6NBAKBH8p
ky94ladtwPsYpFrNOx9Dqj/QsB9EE0nGwuk4cE/QfuIx+eXaMa8hZ/8jP3iq/wON
pQdS/IjlZ07uiZkY2mAeNXWx39YP2NS1Nb6/3diCMzKATivtzUagqpWjmxrJNMFn
RQQ/AHddBCaU+yDjLgj5Smol3y/DwQkFWfxQ3FP5R9Fe6bhgK3ge/02EM0KpdGlb
ndMcARpgvtnwkDSeWd5z3EifACRfHIbyBc0q9eGdnqL2mkflXpMiQuHanDOOTHw7
IarXp8vm8ThN6vnVz6/9GF4tpJJgzk4rBiLybdmyfZrRyMMVpS0d85O4M4BMur25
P38hKyriycMXEgSFREDNZwihC+i16pUy33OuwNdAkluKdmPWgTux4RTB8bN0uXHF
eavnsyfcNIafg7a+xJknazqfsAcx7fw78qyk89Uw/YrE1bcZCfnpSTolHpdWgS+h
FZHik4EsZrPACtkmLnMSj3pSPX7dQhGHo4NEPTn+IXdka6kgUvESrAhFYzvZMZMc
NwG7NlwKoMzMZk314lOosItS4nViijx8Lw0nB9e3AjnmwPQSwI35J9KuhMS4Mbn+
9UXUblt4l+vmYRY3TcGBS6BD/nlF39vr7RKgxfiUT9UrwL2kCjtN41+Ynl/fBKOU
GdzRV2onC+yCaxZg/TgdiBnP3xH1mpmt0IiR1VHb4ZqWsFN1ZqtEFf3imQ4m3JUZ
35m2ykbQHFQrnZsjyvwq1jUoT5MknWTFd4HdwMGWp2za5BofY22EpSquj2IvG1tm
9/GKef2GGw7v5Rze0fkyCbbmDPmlPh98jwViA3O/LCg2GL6oekYO0frLDYNxwUv+
uAqRZr8dq0X5ReVYlxn3BpO1bW7ozK6iJjm5iUrye6jatarRDmUo0tXkIG6KWxA6
JBbNHC3paVpJGXakxg1wPGakjW8UnrL6EjcYne/jsug+y6yy/IU4RJ079vyMOv/T
sLyK+50sOCKMj4I91ztAVu0BuJROWiiz4JaS7HP0/CFKCiVsVHmd1Qx6cIb4vgsF
XudswZ3XBscZHQGFNuqWmH6DEtypyRT9k1PVem8UNSCwI3h7RwDmJwS5+DQSuyEA
mdWNbrXf+CqFpc9mrO+r9Q6VKdDxs0vNUb5Pr2zYX9UKFWsRMzAw0SEkqMYuZAcH
tTUJ9nXT6WAp4PqHGmxiSGD1dA3j5VMTtBcYUFCD4UwzJodU6gvVrkLUGbnaLwwH
IPKCRimprPvDXUfETyVIHe/+QQnsxezIDyP4x5AkkolZEbX6zBCzCddXoNLAKGPB
bFQ/JgFITdrnoyTlI8eFUrqcLYpwkPncxfW+f1sCXt/1cmcFSnTV7WN6xk6sqafA
aa9xf6hUYEFwty+3QEsSiWDM7DyvNZ3FTK/qnFLAfPwTwBPfFcWAUHvyT3myyQi+
+UuIQRY0KKn2RsS7+5zTE5REDfDmCPhcvr8vzQdRYKWBhT8KCL9nK6LpuiAM7CXL
CRb+EuoKbHmFjWBmqUxzRIDVD2BrGU6CNVc/DkTKWg/DIo4UiRck7dTv8N/FmAol
3J5Lv293yuDGPjWSpS1ZXSQKksx/eVdVqj8zatluTCRHDgBBzaZWXrJaHZDTekwv
JU7JrT553eWr3flDpo7aEh61+kl9gcz9bO2fMmeCoFMuzkMRBMhT6j+B1zef/Ce0
sYbsxt9p39wBEVFSoJs3vTgqv88N2eKEatrJMxVlkqlyw5un4DsLbz3JmSRNUrcd
1Fs8O5c4P2dvgIN/eia/DnCP47k/pfA33wbOfA5xnXkqzgHgQhAOnRr8egZoFScz
SilXHUe67RoYgMUR01tZ4LVQkIsSMR2S78hG9lMPowCY8J4crvGc+yrgTwumDd12
u8edhp0tiGH27XmZh3zSXgr0bADOjjCAdpra6FqoUu0Fziqsanhh804DeAIZbfgi
zTBP4GUk11fzar85rLvjeyFNRX+RCkkGufA66gkWjXwMIIFuD3jksVs8hdGU804y
xyk5kPKTA8b8p83J6w5e5kOdy1AEJuu7Rt9/E0WW6xHJP9/Rxf9G3BGEExNmbKwO
tY7S8+qPNWxmcuxayoRDInI0q5P3W94KkQ440t39ArwTujAGDxSvCaP/WQbfd7tn
vJ5F47OZMTWkRfo4QfjsXZTmJZu1Ssg/H0k1Fn+5QAAoAshZSP4VdOGcIeM/BN+M
zYWIAXhDKryZONjPlML9lEzd4T/EUCqtjMZUC4eJEkI8VVw/daBVcc4SKqwOwTFZ
3bNnah88wi0YGfhomcwBmCsNS4iC5q6CbYqg+GZXZjOAIualOSwrtWSk1tlRi2ta
8o7odhOhGoqTFO3t4FAze0mfUPcI9IaRtq6Z7guuk3zBhBQKJosFVUB2WRnMJIB/
lYQm+SmxYajh2dpLHDoA55AkRhvuRZzEfkps4veS66YthBvFFYZCpinFfRV0/Mkh
h5Wi/Bscktr12RO/XtlmlUAaIrG8r93rr1bzerxH6rC+QwOcllb2j277JI4USicZ
jHuPbX3P6GS1R8i3o3/P27/KiNSZQfLCD55SAgBaKYK1KM3ILKTSDMbj6As+7dE1
JkFpdEgHu6vFf0k5tK/17SBDJU205E2s4b52nwciIMa7IfgXgIrkQGq8Efk1Zn9T
sKxjC1hv8conyf9ckzm0Sr4gFjKY2ESbHPEOhDLVlN+p6USpdn/LlCOqG/UvBIEX
V39UkeYuWyuzmI1y+7MouV0AqtXGgry2qjz6rTxElrpMJD4b1twCxzZttDz2ud5I
S/ctCqnj8MIsWcG/vKKgtdYkDpLDoV1BOL+IwutMfv7zV0qlK2eU0NZr+TRjhGri
Q3MIJMVZG609EFBr2YuMqiyn//NBj6RAL58V7UpVCPdowSzAR2ZNBiakgGw7bKA1
j9tBB7kMq10GY3b3k/EsfE1tucxZZ5tAtXchl5vQFMIEgfXzvjNK7bYONZYBDSxt
u9+mkGVwqEnJqsjgcyX7+4UrAGprcgy6SmjGBaz1lbvC+l3ZqpZxL56plTzrehul
HdGF9aOJARgzvyjUlVA+AubOhBua73EgoD6SOWs7Pu2zq1+Sc5hgPgzPa7SILqRi
/id7G2rcOBGV59ddjsYr2w4jYYCavjykk/jk8P/UwZkAFqZ27DXoPRELke37RyTK
cyl3XFa9jexUweDF/culy9AlJ2ojakLcmm2m8fijpNZhKd5DKpawSktgX2fGI/A2
NIoXUNRfCKl11e/Tj7INOwcWoqJnKVX6beYwuLWKAJo5KLAix4439XXa/LUFTNqh
JE3IH7m9n8SMFHtd41ZLCDOIiAxhFNpR6TS+PYkfy0WZGZuFaBAQKq9msprLl/oH
xUtvKIdDQyLfvQ19eq7SPtqk5Ut3AIo25iv2LZN9Kpgnzj0ZS6V+fFp4yYNeSL3z
rhwbK+/CTBGRz3gQpGzvQ2xuA5OCW7+5cnTG/HM8Mxv7I2sa4uYViSspAc1vDxn/
nah0/TpD/vS3xnmRQklcZWkdrx36LxDln4OJomyPXWeoyAk3MaPn+UyPXtJJvc47
ITK3SthBaoWsBD3F/rHEbqtLGl9xPQ/Y3qP3TyMA4VdnX5tKsqY/IGjn2JPLDGwQ
noUzaWGT/v8CQtLBZOEuHLfwsf//b8rL0cr39VgBaNliHHho90k7PI7mczwEaRDp
LijI0tWzjE2UbGF8tNZKSGblfCE8u6I7eYtXb7qQ0EKxFAgKAbJmfjEKQrVY5p5e
c/YhdUNxS2huhQkCgBd65255/HJNjqTarkMSu3vB5U9japdGjByCvQNu33QHG8Cv
mfSzwQYefsg7NeXNjWnuRatmSfmGRQZolPzWvPH06OESFWq98AN/SfjlP4wQjxDZ
2jtNsP2Mg6JkVkkyjhI7UWUBnMUXYdFJuCxjuQoYJlB+dcVmulVSMoKqRNS+vZtN
4hH0gzVEN1Vr3lbnRmAKJL+WycYYzWdXC3O2/Xr0cyKg6F91EroKSq5nVvwGxIRm
d1Tx/8riEX78w376QmbA/YdVHgqqT7Aj2BYJsfrFL1g2p6vLybQnHMnkbEs1LodM
MEg2kGwi6cp65CenqDXYYeymm3F9FN0K1GVmj6EFX92fIQ2UND+OGvK7HDcfS5kF
FYNzxUYXQ/8J2dzCLW1/cjMs3hIUCHrwsF75hUwYzbuyPJzck6oA9+Y6R+u8nwOj
XcpJSvGNb38jYzhjaoq9UmO7VTxzk30gWkjqOiHo2/sCelGoDBe8Jqd25Yc6UmWM
AtIJjSEmSlRYT6kTXFmq9mQV5/yLS0edyoxPI1zLXSSugOlHBovIyRnhcEH8hErD
YYo01nC3qMHZZcKedEqMJHCVK6N6DiNdgNUHCAryktbDVnPVCphG17jCWaoej4wh
Z0/s25C6DOq506joh+irOj8ZrZqsP3A+Mc5K7jYHIaiz00CICJ4VLyCI2tz0F1WH
kEeKfQlPvtePFp8wYgn05lS4MlMM6/0hoSiOZu4+mJBgIwx/kG0UO61wbyiobLYt
dTaiOCLLodtiVvCbVv0v7rLa/R73RD9QugbUGE0UlCIjza9wILNfgbu+GvmeY5w8
OsK5OgVL06TPA3OTzAUGIeahPMx1KEjifeZwYjxrpSuKaEGfpCiMIityU9yUXoVu
3pKEhjTH04aSC6mIVyznYSWsU5nFEvl/Rf/iYRO3HRDREAnnCcY/rkc04thp+uK4
qRf3I2GhE9hTTV3Sw/J9HEAQa3aLsKi70Vg1VANnOGTiIvOMooDZiKd+OD085/fe
nYiddqi4zL9wfMHjvkL2OesTZB8yGxldXfOF4TL7toFhoTNI4aaT9AZTwnpwyw4l
MEAn3oXg7JOFE2qU7X+Ib0rYlSJNI5cAq0/5v/k4Dj55GBy6ojDJAvNUeUgQwAxd
tOR49eNgSBGtckq1mT7ArFKFjwwKDpyGUcRZLo2z9rcBCBftrKMlj6aDYt7XYjjY
egV1EPEEJ2PTePdzAA/N6RxZERMVDI8KcKvNMkgfwgz1KykQg9SUM9C+0JDcs5u1
WGzmvA7lM2E+GoQyYOGcjXwDInoMSgh1fJGi4LMMinEiHwHrPBQ7A0gjBmfZRjY8
VYedmFy25KXhUpd2dS05SoCpbIdpr3SZ2P34OnUYOTPi7yK57rSg29rIPrUFgWz/
f/ra3FbLX6Kt+G5BN9XjQYnaRryj5o9VzR4xsmoSjK2tOQMUzMzmJNOArpE1omMr
vahwFCIjuh8Tzo4nHDIdyyBolW+lm07GHhzxivDqy4RRNWoRdp3U1gZ22w1Ftq/v
u3NzKKLciSAOjeZBKQ6bjQ/soQIPAeeab+XSrcDgw2dKVoKBYUqYSM4pj7XduU85
avXXhYJgVld+6wz57Wvlx3DoS5RnrwU5t9xxBPjDZtsF6hiaP3slooQV9s+A2AIw
YkLDizNuXPPoIiBXcR+QzQeatkvF07ostPm2l2Tcb5Kuk55vgdeL/cJq2/2Z7gZW
xNF3HW92Hwr7ec4S+luIe1oN3mM3oD1jPC78hyKEtQ4O9Pi/wW8MFcuSrHkBiISz
XKZ3Tz+8ZDBLVvNDSbui9k+vw0Y7mHl5wv46LG+raBhAaVS+yUPyizkVj30bhXYA
8/R6018xM+1SnsQJKdVzdEY9d+HN6Hs4oYpoyCoYoUA8g7SGCmuUlNQLH0nM+uty
J8WyUoL84C1mjU6xcH1sHGlj8cYjjdOXNWW6/TV0qN6zqRL/n9e0ucsx79/8KwKW
9mKKZI/8EIte969k34D+H3Er+WoZGL9m5vss53mkaph6TNhYTPqJr6fXGI6Gh3dh
vXk9ZDnCL3RQhLEGW8nY2NyEg4XGQZENbZspn1eOSVA8fsxVOUGSJwRpxH+IeVyq
BNHM5izFGV7WzpvyfFcpp0Tgy+8xn6XJQut3YODmfN7CZzqflcG8bg5NkcINK4KE
HWUJnjh0n+PUX8VDIU/tMF594gsKKIDPXyFSPo89n9XR01pn5dFVRueQpe9vGUjo
ickWU0RcWHLorhlSWjNoFpT8cpYuVTYtsTRX1YTVzhA3AR+5kww9ARDbulWBp6ZC
/2/6407ceEFeM/Mk1YKNH3HG0Wx9jnRBS6RO+DD1DsSrhmLA8VvKaMiww69i9TTj
XiVIHS46Bkbq08C3uwFmlRIst+JbkDgFytEHtlvQ1x2NqCsH7SAHiN8HyusvEW3o
16ISoux2R8m/47xB/SPif/HVseMoLKTLBkQUx3XASKPyk+lMTRY+5tkclgEgI72U
p5MLExLKDoo3QN+Qx3fqiIoXyr0PgM5kcMzg7Wwxog3wv7V5R3EbOUy0/Fu+K8eT
Zf9dswq1+3oubnFpS4AkFA0D/QvBgjMvqagV5Imu5/CMCH746yEv4W/ovKngS5D2
YV0Jy+K/vl5kaqRRSZROigLD+XmqYyIaggKu31MK+9ICVAqO3EbmZTLu09QJTIQK
vlfLQm4XS/y4Fzoa8bzQtIixDuviEf0auilI5g0W5orDDOSeiFKoVtUvFyYgbexM
O/bVfA3HxQ/6vaa28e6onX2f7m6R6PoYBlsa10zMNTejO1LABT9j/3teSuBisnKk
6bTSqOWli/6UELFDD8B8x7DJkz4w4nlTJX8Y7NyBDIs/vAT0KfoDKPv/rmp+oE+t
pI/t7nLzvwUbogcpWXXa2BNmOOUWElrnXbM8Uv9/yYJDK/SeXK+LcNC3FeIRRVD/
tlcsM4K96Mgw8nFIHmkN48vjfgI55KqsMGexmbciFzhGEuMYbG1CKaJw6Qo1o4YY
ZnnjeZWW3bxONzCKrcF9llJENAoBBzCNBPXlwFUzV1hto5ZyP9q+Wsni0oAs+2In
xCg8Gz/ec0ei0jiAVXKbcRW5bxWEexxLwaa0rUgR16EXyxalExJTaqJo5UOQKqAH
zCex2wkG8fwQkZg7M6KzS4fUIpp1h7E4woNFFHwW2jmTYWPHnjaC7DJuPX/sSARg
a7+4Z0x6yotUe4pdvOxeEs0+GcA9sf8/2oEA46QUoLbLobpc6jbJMX2tk0XXa34B
jF8L/vw+lUAqtJieA3ZxdEHoY29/2hRnV6MGKI7c2E/xqEp4yP9wdYSaeeQIuECl
6N3qQdjQ7iMm5cQlg/laDlY+cxjCnkdH7fbEUzsynqcjPahkre3SeSjVM0okqWm/
UMPJcYr5yPqArg9jCSD2sbBzjjcQCo1GeYcB65F6VahhXBF1TavhxPTuH6faU+ek
Wubr+puZdAV6MesGQcusQxiicSyUkJqR3VK3DHpNBrtYXwUOKsv7CY2UuINIFZxY
OU/0dxZUDcWxktPDomA2yHk4ZIx44YXsoxprO0VIZ3Z5GtKIyYQbufMgc/Q+ah8W
72pcyKDA66WEjM9kbVuLzdDGuJbErbA5UAm6xAkuJhzp6ePiKFFoeBPRcRZ1HYbr
ZSIIQtKg4COTsvYxL5iERV1mQifDRPQ38QfK7KoxMzTxRTHfMvU3+mRk4J7GMvEa
q9XPuUbq05YPoJXf0b2wtk9cgHrVZGmsUzggx/N3lYbTNLaio4SjRVG5kK9olRp8
A3N63wkLWC6IsG/o+/ayJxZ6VQ3UkQTd4KYh8Muybm+7+6vHioxoEH6Y0eAA2PxH
x9L60EiFT+cyNDUX3nZM5Z02t3jl0mrVmeJnUqcy2qDeJvBULvGIRHClbVXbzZiJ
nk7+flW+XbCa+zvD3lOSuI3/Z50LgUngJU2aYpgyXS0BSA+/G/w/qOTo6wCUQt4B
BheDya+J/yiPT23KxIEmigjq1XCVRJ+GAAugXMOMdXBbhEBqwKKtcixLVFdKvZqt
cQ+Wo7Ucknplgixj7p/8xPUwcltDNSr/tjb9xu1RfJUahWpoeMOZ7KPvgSkeqw/J
Ek/1W2shcwRL40/vvvQdyXM0rpOlvz2Sk5Dq7qLVSz3JRjf0Mowhp6Z9KbwqE27i
BeIrCvI53c+VQqyZhjCDg+Y+ROPjHphWzTzJiMOUUHE3sGKhVfd0fzLzTs6WhgWA
7I43g82oP++f3ByBW6l9bU45kKrqZarx4BLZ44DyzKkP2G1LKYSF13PNinNzoC5n
JaA7duBpWlUP2awuaV6yDQyg/lfNkUPLhv2yu0sqp7rNuViCM4wJisOaxXW9Ncrm
5//cY15sCgnD/6v4QUrSnSXpWGitUe8RhTYTKwqzgBfK7BcFJ67ioFTL+evXzW20
+kjogfhtOds9dg949fKMU2XLN3JkH/Cd9ebR03WsKeuMGECPd8bNYgP1aQfZzM/h
EbcpLKOdjVMVZuSqyFryq+BQTuTVV+iVwi5JdOt/qjHheN5MlJpcnkoQsRRM8Gcw
M0v6ycOs5vKycBAmSy34nw7W+U5FSBPxKmT3lEY5MGoKkex9B7un0mAH8f0sXX3y
MW7uB/EAPWRKICFcoyyc7MKQC9YQDVkTU61LtJK7YG8CBurCl8fKHvZRund1HdB/
4T0hs3TrkC6H3w572DPQAzUlu5O9sESx2e06EYxiED6V3TJL/FbaEUdw/iuvJ93w
Xf+S+UM2x7DH24K+I2N4YEh3veO1AQbVr3OyIqfxyi9QBEvRfQCQNmFoTm+P2pIX
qHwbSbSgDeVE9GnMV6TeyMLfBqzgY8QaXyHmqc6Yq+tk7oWU0tq0EN3HX5iWexLI
dMcwhBEvI3su7etJgcs7p2+r/Mz8PDJPz3D0EhsN3EoU/8de05LCYIsrK412KitD
DgYQ3kxY1pC7wRB8mfJRPVJEwkhmWAyQ6Ehnv7lUfhdC0YBorRUpD84fMAiM1A1z
oGANtr98KIIG0oeHHi90xwq4MC+CNnW3nnZmG0XCxgOGa+zIV8gIMSD+i05HIXTW
FEy3W2cj9HgLb7tGipVhWOpZN9JiN5o0Bg2KTLP4x/qnjgj7cPEXryy5E8R02a69
0hLRIRpAmzmJoEg3w9bfqlv+MixV92R2y8nci1r3VnNJwxyxRqBCjKzPr3TaXMYK
MKinJx57tUG2XAjEur/txWuM6CnUu7kG+ZDSt4B07PE/cnKKSc6sJYcGJh4p8yUR
Wg0r1NC/tDevyMuufbkCpD995Kn8MrsIpj2RS3kWVaPVcVmeJeCKQYPLZpFCpa1F
GxEoGKARNRljyng3VnFheS6CWt/cSCqGo7TIcXmdGP/RPHUHe3hj+vo53q/fVERw
POxFJAajbMcHyMatablQ9g+4tLzKdeZIePKAJbwR/rq921gmXPTDCXyDwmZTu/d5
UZY486iiCA/Zy2p4jdyx39js/wfz/STvPcRdTBhlhpS3TcW3EN65jqcL8IpPdWO5
PS18MB+XOcdIutQYcYIe5RrtMu4mP2Y0h1K0WMdiy13ojItIBvBHbSRytYMPjFNs
TsurKgQou1i7NDRB95QyulA9wbZRxS/UiMfctEGUf+scQtqPFmBga/8vfPdng661
byjTm4AVIwVkIk0b3X37MjyPqvzkoLDPH7n34hihcTxQK84YzAiT+McrEiMjTtDk
+zJnmKjl9VY0LYJr6ZiUGS521dHOTMSfsRSBSvhY104qqVHY3pr1AS/G9xHkj3KV
IAKiS1C1k/ECbf0vF1EAE2DTKKk1QOZQChz7ueZDyBGimV7bFOLeUcJTarVcU0OH
dGRJmUYicmGKAaPOsBfIfyLnB3NgdcnwwdLqkOx3XiLl3eeFlZUNgp90+X5kn8vH
CwClt1WGyx4acX/1q5RCPyfhQlIkqS3Xe+X+YQwVo1vXXd0Av4lYJRcfrq/uIZ+P
Dwuv7Epg8U/VFn0RKQdd0xqMB4s09lCWmuXWcaV1nYvqP81e8jj9FWb2XpujN8gG
mhkAHGt6f5ybBkMFq0Q6sNZHoepVNuKdG2aoNysEyrsSzJ3EfxQzcU0lSYn+eCob
wouyOn7WVcvT2EHJeco15Y5Q5DKM3+RmpH/XpCNpzOawdlF6BwBqZ3G2LCqC5Nkc
mRTowKEDIA96U5aVyKUPiF5SVO+1ZdVmgglNFxlG+m5VXI2E4DIjQvkTH5Gxb2KH
4VcoG5jZdzUDR6Sln3gqiZNHaD5Z9jN4Fye/tigeybxSUBMCxCImHz7IbNoyLwQ+
vrVsPcUXJ5ov5ooSEDg9z/k3+bFOw+GT+ustSSiTDIIkn5JnP+HHPtxclFX8r3B/
RAsAMYz4j7GimYgmO0GY5ivdpJD97S5nK4e6tgRk/5zqqdtrMw1M9zraZQm8rd+N
9xaBBjJQ+b9MaUN7EcUETyFbFUc+hK4I/v5V71ReJZkNaWQH+c9KWcu2Qogms7vl
v0pJOZyi4nDhH0qAl8VajdUP1tIJGU2TQjOAAeHXhz3V7FlacBqFW0Ocsnf0khsM
ePt5X1UAvjhSj2eIxKkSR01TjHT+gxuPHGigMmOaNsry3XdZNXJi79yqcbYyt7m/
NEJYxG4X+t2TN9DH5X5enb7Ukrm7NZt7jXBVKP94sBsirNNvtjEAlos143kUcGUz
rbGRKJC6v4JFtTzSorEYFQ91mumtFbti95J9LpBdOnn7NsFRT7ABjfvjNDgOQj6p
CTunpSBQfVfL6beRX+rkYPfbp45kzogn4sUIy0831hFK2+jwXxvlDV3YWe8+Rh98
RmwiiwMy34onNMrW/ja+0X0z2rEClBUZ54OmJFRrlg+zQcydpqUVKKWCVybSexCk
A9E6iyHWw9rNS9pt2wZ92tp85+njc2q+cqf99/NaPEC9GDM+84mABgfi4ZL7pBwB
/bOZLSFbA+v4xPUTpkkIxsuFA1q90sEKUYsn0W0DAZoM+lC9psTG+Ud5pOisAAxd
nR397P6OQga7Lv/iL6BWQg1nMYBinGKl86PMv4oosbyv1ITqRI7IwmF9XP/+lOlv
aMXlDYOILc6wbKpj/dI62hTLfwxDVxnvvH6D+lxrzHu38P70vEgZgfLHzNfeKISl
X9wMIbuZnkHnnoFLOqUS7SU4zMkPYLdpLy1jUSF580Q2jGF99BlqZEkt9BRuSjUE
u23Tb+WD1gkQgeU1eVNHQt3lLf6Jej6QTTxZrA5V7kocgTYpw4NeruocR4yRzLNL
HJEaw6j90HEG1PDLSfuIbtH+A78MNShLtEQ9iGg5q4rOZFqSnyWWtLFL4vJAHuHx
PWAAfXD9u0LVtsPbZMpBKZCaCBt1pDS/ZGgGWVLF5fIEoaEMnSys1TUtN8pLJ5+f
f/E83hnT8UIAyTosboul8zEktVSclCXU1RSlC6fF9Eiqr1r/DcKNSKN/LufubPmL
LDRnwd5VjEBeqTZ1rfy1VUxcq2JK41Iwo96KaqHaH4D4xf5PVeKBStOTB2gTaQZ1
FXYcqcH0v5ONgwcJktveKugS1xIACpggepPUxWpc24s6ffVXSC6eQyxopCB32ibL
EipfysOO5CmF2DlPsu6IUOIS4GPoLQHEFkQRUdBwrmvVi07zAwlRRLq4GhIJUdEP
MLMHZ2bY/HArnJyj6nGPD796E1AVIgz0WPYQY2xpKzRMXlXyrizxD/MJNTbSIaZc
bB1NHFNuuAnVbRvpwNApK4mFwTlYnGDraQnxyzpxuq5XKYBBMee5WPgYyXcRBK1L
KRHjgSPvXBQ4mou6z6GA6w6ChDllx9PL9uzQhwTkoYQljdog/GhX306bzgkTRNHp
q/XHPCPas9HaBMv6lRRahQYQQds7VOk7RucOfn1xAL6GP1hP7p/urf1/AxuYzJUw
hMzp6iTxZp8wBKcQcOc8LnaMwSY0Nv92USdoTFVNojzAd8r+dbcUbOm/NOW0NO3v
76Ms1YjQoTt4Qwyjo3TPS96FmMyfVs1ga7o5ReFfYbJoJuuSi/FFm1gZLLl+D7eX
6mvS0/LKdvtpAF9gOt7RIkrYG26wGiRcH/w4HWRIoMCjpV3j0iS3NmB9XB4gtj3Z
2fscSFlBg1xya5sYgGFOzXu77ydDXEHOhvnXiPWG+APMGas7kPtf5+bTWg26bSM8
NYJjsAFFzcKBmt0guJJbiWbspL1j26Q7XG/FUb8SdkTuiEkrcJ+ZAIrY7VzgfmUk
+DeLv5pZdBjyZScwc0gv3u/qvXhd97y5VaY5PRtbqL0xPuCJqUyB7y00kBsUWNtQ
0hN25FpxqpnhNqoGkkYcQUvGK8uVZZqmHs+jjNmrG76rosD8B63xrn6+G43mkTpt
UKOybUl+GPtSzVjKZO4dnzZOyXFQ2aFQ4THsPi3ys0q63TBD7kOkBact/7HbAXf9
gOLPKlh42Gs/ROm3zyR2yp4I88lJYgb67qYBcz0smBCfebGez3V+YYjoyfm0uMNh
zfIlcQYeKyf/kk25PgFmj54WPw+mnTtHmi2nHt+iKN0U1raECSsx0aSQR7hElwkk
814U1ICk9cuk/VRLmsA6bEaHLnx7wI8lTK4iOraomQZD0r/13m57COQDefQYYv/Q
Tut51RpWvKFLyXzajiH0J6PBr4NvFZDwNZZfgYbVuF4RNGleiQgEETOPAXbxaBG6
L+/ZyW2BVnb8036PoC5pK6oQyaRzPH072E3u1BfXJJDYkARBj3jZE5Kvm4pnw0Ge
a3bHSfA7Dd5lmMABCETurI6DU7bl8gxhfO7btiz/qlW6QzvOKZDpOLLovHCLyxFh
dLpHuznjaFasJjEu8q6lNL8DrkLpP9GM4zeMF6DFYxA3jLx0b796zhPoKErLLgcq
V6VaUjNg/aPdHT6Jdd7AXnv3ZTkH6JMbJfUf47lvyb1c7bckKtFDqvm2WaLk0q+Y
YMpNnfcUdOMBNSU21RF3scDIQjjykG3+0UGZ9c4AaShErmX2Biz5D9goI9offaR4
AGTr4OLUL5eP7Z4lTYAohtuKApAZheyEAQFvhT5HF0rsGy3NfQWCAMEdTe58AxM8
jbZREQZhh9vLEbxyuAd6NUxycBwCxwj6/NXy/R/VFQcxb7K4SgCmnLl5kvnGj6IU
slvBEuPKMnl6OlhfAkneY7I+nz082WskR4GIlRsZ6a1Nn8tN3yKKEaVzLz3INsuZ
mOsdc1SGtwj5mSg3LzCfGnzuD2vIH+AUqkuQG0m/rMau2lVH/nor4hHFToV9+L9C
HS5UPydEbtl80zKzMnnCxVOJ10kwnioHFAR+mCSmzjXxjSkSpkt+fmfdxNJVK81t
o8jgLrWM2tCAfk/MqAxLpnnGqAkzg+MhywWxqEeOvfOsCbTuRbIT/YHBRZPf42Mo
zAH0rO61rd4Vjxqg25Hj8ri3kRZBGHVTDebZAxxmZ1FngD2UmWdnC4+/WvzH+rCd
Yw3Yub5gd8mtcOchA3pgoOYIanhEsPVYW3VtJdFAChHA+w7uyKsLOKLbJLm/efLT
Un2kU70U2Cb26EFeRwHblDK3OwNWzVoSgYsHAND3AaSfYasitYjLGvSPPB0GONqJ
/7wXVoXDH0b8Hjt/UtY5eUdxWkVxCnsMvtK2orHhQ2rs9BmgC3fl0lMghOIedc8c
UtsmRdJHtyQZo2UziMt/8+EDNLQkJcwNnVYKK8fZapTs0c7bYuthwopE2qWHI1nO
vBKbjAOCIB6f+SKAzFSC8bfl3BsFdkY9dqS8tta5Ln7W39hR9HvItYmqBaEolqyb
xBFxu/8ohbs3BNvys/adNrjo7F4zgkFHV9YuZmkBr7akkdc+kCaQIDNl4voFN/Hw
SusuAEYMykaWEr8tHE5Km2Sq+DqtLueOreHz2JZKOq3lxUYpo/v537A7ACgMa475
wmCufSf7RPJMlArrJz015fIgiEvSL/OzLwEMp17KJzc75VZgUj8kfcncS9W+nKDy
ZiuQBRWA2NsEp5rpwOfqvTzgR22virsvtizoqSTXZLpRItGcknjCqzouX15tpKcB
MV0ebl14/Hh6u1Lzng7PhMsALLzi8zFbY5pE7GtXppJcW7yJn0yuAI2lOsOYYr+h
0rk8wKF3cVyZLgwGDChjLwfC8PcYPPwHw1kEr2vktaMA8dZ3TQ3Zlh+EBo1zDdHF
WuhkIJq/oCKqETHvq2fi8LGLMNlkLYyySYqoYZ5rCJ3m7ZQjuoH347VrHdQpD2Fa
+frqxU0OczuGYKjB/XjDlDf7/F8wZ7Bz4k3rX58FUFP02z119U9qpy2MIsNSFNUc
mN26miGYtRz7A57ya6FbUqJrA+Uy3z42JaEUNNXB8xPLvCP/KiwKEwrqCbx+8EJR
K0Gbvk2L50SKQse7UIisc63k/GGEvnvC4IKhS7TRHVmrBrKjmjEzh9UE5sPV6ne7
4aNz3AHKNm7EHIvkRE3svXPi2yc9i6DLiMbYH32ItVQaPkoLD224F5wf+Pe8SqIE
oJ7r+s0Mhl3iCtrYxdf2tlSE4Ybbxj30rts0QzWC0S50Tc8MzeT2S3HyafutDoZU
aS0gGanTrqpj3GbWJNU2kxyPqrvFh5c3GgLpnIXrfvghu0oqluIoYxvPLNHduF3+
e1ZwLV/JmnKa2tfGia5gDUXjeqfKLqFwdmLq80fjU+jh/cJvkB30qpYHfyd0ea1O
jJqZtF3OS1vRaf9ajU/IUr0oaUPwrCoBKXNpqN0y9DMibXGrvjOxIXv4+LfeD4B2
b+8Xo1520WLZCARGrVjED8pLhZsDhOc9ON/4jU7UbF7ZNIcBE5Z8qkI2WXt2luuI
TEMI803Lye6SyNp46TRcYz0FE0CjktOtXcE57EGJn/R6LyhoZ95wZgt+aXbMBtBE
Bnt1wvChYN1KoHmuGbrgnLUO1UYYXVPPeHU+B8r7K6/DGkqQdClhLbajmO9Fpt2R
2kIu8N1mBLQT7qCw4aU7TEDp5YIoXH8ZFtKieUafnjIx4++Ir27ALZ2s9KnM4cj7
0v0H0z5Zme4r1iC3uBRaE4EiycJKlv5a09jo1YnwqQSd8woepU48VC0Aa9Er/UA3
wyF264oo7bwdpcR7PAJ/3aInGOEIo4Gij8hkz+5yDlfEao8Ono4zdntsanvuVa66
XCMFLVaLqjpVS+ETGPmK+ICt/k3M047qIya5sKYbGi9f12cSPPj7Dy6RZz/Ff7qN
sXKgZNVFucpXEjIva3VkAbs89Fv7rsABLrGv/6iP7nj6ircqCbgk6h6QqgNf1oTH
XPbyFvVDINHkcznUNBwAqMQELt5gTZaxAVdU/4QFdGXfyP5OrZPZjb5qOloAdLVn
gbqyhekRxU31eBxWFluxXeDIIIG/LPriiUeSukWf8P0KPnz1Qqe4ltycmpIKhNru
63Fmi7y2eljP6grHFkSiES8xSCRG8F4mus2h1FBZjxU5Oy5Lz63M983e5/Yhl50J
582vt5tbbTizU0xBERtKdJEJ8NCFAPBxXwl14bU+RYcgg8wB4TJPS0XmrexaOqDQ
mqSn83P2rgS7NMfJlVWbrTqDTKID8VVTrea5zJ/Mw4X/hy3xKxQl34KnVAJRrMzK
Y4yz84YzzGvVKEpmbtssg1fF/qwGMPpkYFmzWD7nxQwdOGb5uh3mV7gmpSQ36EfE
xDHP/6k1TaQ0KuG+8mWokLtoZxWEK3DhpGBKjA6Dw+CeSlTAQDsnkg7wB/TBJPFa
6A8DWVjQGM/RSZGWe6cTaXR6cwSgTKgAeYaGwz+wB+q6NEy1bU4tXioNq8Ye+2Qr
2KPjMuY+Xx/wcXEbnC1dCNeLHz9blmW/H55NX4n4fv3VAsJjBfQgLFfrWbHzFg5D
Z5/0LJ6IsrlMgczNKA2VFtCMXmNYsBxXIFbomkumJri5UV9i5OSHfEh9jyMcDH47
oTmQBAymdJcA+hqPq7CtIXJbTfnui/L/HbqgUz0LreAiiaM/ygkcYzOR30oPDQnP
kklhQS/+uGMNDr6PY0Xg+q/uuSR7ydQXctquB9dM1PRiGMXa5bjhgnWm+Cq1N7gV
R4U/qEbxzAgETkJxyjleNOV28VfFZDV5Q6eQ+wLWXiq64fTeK0N+BBcnd8FNYduM
PIZ6F9sKUr0hz/X0khSO+c00mNRxIOufZYx90Enh7XOB5JNfyZmyb4jOvK+W2ciw
ub/mfGAfllSuOIu4CL95k8SsH5gTVB4TA+0+kmtlgUw/6AwI4jLoy85K/UBZUlbI
MDIgyypdDN6K6ct0UQXOc9uVnm5xaMhi9SQXwvhPgzNIAKUjTFtTaDcjDvySELYW
5JyPfLRlIy8/catWUpMtGIx6oLK6T5sUzTF9qBvWx2xs9J98nSm/sgkR+mH5hIm6
tEcEJa0qh0e50+DJXW9ST6UEiR5T0UoCOKRyPgRRJICQdhcGNqnX4v3mGb/4cuNF
H1YDV8jBriZB4mJC85N0o2c3gT0pdP9XNO53uEnR4qLVA4NQRMDhR9JoJxpbpFe3
HBCzJu7dELBImqRFlR8DVBRA7c++vB6dfxW1ePJTxq83zVT+lnayY6GFPBLlQg1A
tRu3Wzj89U9JcuYf/LSD9s2evrIWb6n4BqBkSMct1oiTNJb1NKniUe3Gw2IBKC44
0W/JHQB3MlUCP3jY1ueihJ9f//gtZMNGyzOy/g8YzblUhOmcOh9uW35oVcib2Txi
WOF3r77cPp9Ii1ahOMGCOdY+Lvc3HedFDO9xhZ+ygbmZDT0MmciU3LmicWr+CfLq
bZy++hdxom5tULkEUdrh2uNv5lx0ApW6gqm4c90HkdiASe63eTyH0pAXeA5gvPA1
ioRwyTtQQEkcNFyQOclXOAIMtPhpYyb1eQT60o6BoRkD90ZpA8dx8GVJHqOPocY3
YE5FwEo/C4kZkM7Qz3UtjkJgN+2/wTRhg9YETAn0R4tBjssHQrB5EOSt8+7TNexh
ELFvwIruldSuIH30ZKwgOl2GceV6KDZxJVfZWCizKJIei/h8QDZlzj3qNUGUfUP3
PTXIpPcxtkwHPSu8vVPRR1ObR2gKNey2HMdNj35klMHLwxD5TrTzkh5xOytPZkH4
CDrmf/io8kovB3w52FvNKDwFqc3bxhEOhVAZhMOo0CZR277J7kAKePo9I7FA18Ae
EWYbrlIl95EwF0liQLit+2duUB+fI4m5U5WPSvQQasYh92m8ZnfstQzidSYRFBFk
RfjHTJj7Fbe1lxbWg3yWDAoUszCSSOpuIexsQon2MyTeOYS+ZEUyBDNXCeXSxOx4
gT46pEERZhifkvkgXpB2crKrbBolRl8xQ88Nd+cWZ6TdacsjZrjIF17lmpliyLWa
YfcikjDCibRnX9qrdI9J+YxX7ptHkSngc9JiHO3l5W/rBECb4PThfQt95nvvuEKv
5+caUq8ahaNHYGxGe6M6RHbSCnCaO8x43lbmB9/SAnLdGgXA6raQlFpr+50rft6p
x9b9jz7UCyH+jV0ivifyyP5QvHogtReRHQe8j2C7987XHYhkEhZ2CGNzgtCZH6Qy
9ZP0ketVLlEuKncZGgdDk/8PqvTFwZLwPiDuKqOF5TMmoKKa/lvwOc+WX+pNPZqS
t9QvXjitE+fP+1yuU3KdOLAFHr38MMtUzkQdabBOcj99ao1lLb6orlo1wkui5gjB
Z6ygiLKBv1XAx4Hhn2Vb0lUiVpTu04JNOkAZE48yl/wabttttxRYaXwGOgZ8PBPo
7AtpM0iluhZJudaw6MpX/7ArHDcuv+VMFEGoczua8koJ3W1AmDqI0G8MHqhhvJhH
SaJi1HI2lxwwQNRkirq+mEVDtKKvAfH2TOn8ubqbS0r8J/bisnityGkYwNrPYQuv
zcNWOTBlDFL80el7C8pIkyrzWbrj8qoYS3CLXbPZHmlcTFr4aUCxdyg1qB+7drTn
DWQhf5+OXoYOwYF2E1Z/W7k+w6MHe3rpLkFl9oxOvMWvh65jgeCBSVs/r2QvTUFa
97r5T9DgvsdOgT1kJMnys6+E10RQOFk4YEF21OSeTQ0ufHdIWh/a0bb3ClcYMybg
Tb4PNeZ+A9mBpevTA8y3TFPSVUkMaW60KU/kun082hzYJeVVkoSRtIzOmPfw2pOY
/fYQHqzW3SRal81d+EvTeK+CK99HCtCw7+PSRTiiuc9lhcHGB5o0Ilz7/1vI4852
2DbTdPYb8V+tR+rH4p6iLH+bh2qfeYIswk9bpGKUjKo7jnMNq6uK2oKHMm3Qubb6
I9USQAYnzi47QwtZkeRiDT741mxtpFMcC8HHPzzYs/bfE+Slh772DrStOcXOwlhs
oNzJw+1YecA4O9DHzJIdXpX5gA3JSqNdQ85G0vxJbiRhQixR4UCywhbUqLC/IuLT
sfg2cGuKcRLss2i4J8VUbro30uHUNImiGR7NEpU91hgTMmZknUCdZAmK04alK5R1
DU90WSCZIjkLaVwqrHIs2+/OFs7CywrGJ2MKaWr7CF7G0T2KOL/9K8LlBU9gr8OL
ZaOLr+k6TkXWNU7fPv1wTtOgRWN2rQhgFqD08aPdPXK1goDolzxcjUbP8H/YJ7s3
aLOPST/rWaUsZA7X340aiws1ZLzK7lO0xmORddWVu9k7fZxmPujUpZ+6D0/yefKO
MJHt/Ab7lArAs6Orze0a7mJz+mSZAdZmQ5br7tmMNiPi+QKqUBL7T26kUb8d9eVA
oOQyMKhmeUhjRjeDXUxaqWhf6Ncp9stEavxoZIx0VuEfwMc/RXlsS6KNScNFPFrM
7xr7pe4imjpJNPhppXsj2BVbAQ/oxtjtDIoIm+waS9zWqdKNU2so28AZ289MSpwh
4ZOLAmZmx0xrfQlDQsEsHgBN/VAfbkNohGI9sUNvcZm/B40rHiQDo/OF9kXt5uh+
VJzgdg2fLvbY162bBvniVdoH0ybt6V+MvnuG6aBqYrkvppPTGzQLM14vbdnKocuH
Os61QID01QMiy1/HyETb7QxJ4OzuK3mOM3whMW9WiHDBV99EHrMRCtZoD2VzDic8
OT522fRv3yBENVi4oWHXrYYGt534sURizIZnky/qdtzKAfPfpHFveKGoElrglGDl
hgFFJY1bu0+iH7yoiPSMzOd1YhEpmhl8wSz5KaM79LeOTVTFTEWNiglVOuhdVYTf
C80Pqkpe2b1ZkAtrc4K+5qqo5TCQVCgh7TLGUP1O8vrLJAzoQX5eBecoWO5drT8M
HjP/CYrtaD+Yd9YkqllLpGDFHAkJO3OiFwcrIBTMhynZfwSHLOeyZx6WQrkFT2u6
7zT0WLnrlhZybIwr3gKUPS+9rP3APiJ9YTmnQvMg/luBzi6WEwAQwWunoKqWJbyG
phGU8WKZD4aJy8O6ea5Wi6mL/Jey2KiCkliGBk6ybN13pvuJRK6QOohu+YcpeH+R
mA2iqhYmYfBi2NkxCg9Xr4vXwV5RlhK5H2dsg2T+4SzdbPDMtym16nnIurSOH4zP
V95TUjtCkRDQIV48uixUZV+Vo7ipOHP+8iIoIsteInX2QdW0YNXlhfb3Eotnd2yr
DFVWqKiZi18go6SB5Zz1UCYHVw+F403cCXpvqQdgS0+fvTh3Xgk2DOxj8Bak4ckS
YERO4F2XzCRAWYF2lwEk/zLk9KZOF4KV3uNHm1Ov4Fv3FjFzZ9xZjR7aWQ63Q8Ph
4caIxfBAM1i6XYAGzOArahV1Tu2ePmnia7k2txJnOClyzdFNOjvfvWvHD/zUPyCD
4gOhAus+iRKTOukOarxTBADLiQpJIkLb+7HvoP6NsOC78IqWELrm3HLJVORgx/Iq
oxL6lcNHvBLoG0GOcGQgmdk06Y2dDDIPd3DjpXFvIBr4WLcePHapnQLqRFAYFf7g
GOtWibB96g3Yg4cWpB3nhhSfpkm/TA3V3Jjmd6v1yr6EHtoQounyjdTqEcPMAtf9
s/b154yhc6xUex0gC5i5PE2Mc2A6a72Q2O+B5wJAq94KifS8HTs6EFYdCUQ5Vd3b
Gv5vuSPsdtzenG5iYd2h2dxsL01zTEc1Qm/Yf2brP7m07bSw+VY7aPGiX1/wGjnb
OlI/7jK7eLJ6gAJ8UNu0amULLZfaZCXRQo5OE9yvFabW/315/NRgp+IL/3fjj3BE
/XA50Y/FuPx4JR/05/o+bbnydq7Z309YRVZ9yp8MZYb0aoUhL1SZKVgS4B9uipPj
y1h+SpoyY4p1IJtSbMdW45itLLcwdPFovR9unQsYZaAcL6xm8gRE1YXn4nHxKzFP
rZX9G6WSU/zvV7A8JIK8e7jrxwmX0h1oBKFnNgezKz2+8QrQxmHfBvtLW52I9Wbl
OHwsh68JMPqx5Wl7OwDjmfIzGSmPWbFtnCK1ENQBlCBm8T0T7Hv4C8yItX7Xbi9A
nJR83FoYig1FufGaTTVnw5SUiCaTuJDGI7ewvMkt9NwD1BqwX1ifRXUL0Pv2H+Vz
JhO/eeGO/RXH8t6Q5PEBA7KVnOwN3yfchhd1/PcGge5ExVVOwJaicXDtmUsCf+/S
A/o1KcbtUEEVk2W84+ybb27ZCEbUTr6kXu5vvdwV7hwpDqAN6xKE2scWCStFpYlS
frrUz8+GsxiBDKNo6VgCZali9QQiUgI4moYje1RJAJC8TbfZGvmde8GxLj/CBNdE
GqH8L2TfwzG9IEmigrP5fbEO1Vw09OSg5HXGFLZHr0LICRbD+RcyeIyy7AgIMMRp
taNbl6ho+tYEf7aNrePPDnL09UfsZIWu/V4y79KUigJKKenJyk9jxuMJuAAb+aEt
qH9LZ+ISNLgSuqRUzY0t/Ng2vaJH3W4VpIaQnWMMg4GMjyH61WPvSOFYuPVDft3r
sg8JJZuA910H3Inh7o1MOmeF3MjFI+Dzz+cIWzdb0dQ1Xs4PHh+dXSN+MT0DrF3I
25qtqCTEkFlauGnWQElC4QiCA4slgeBYSiDI8g5kBWdxRV9vw1R4xnYo+61BrXGW
suj28R1N6TRXTqzjnM368qOYc+a6GHCfiEfcCYHh6ZyBhAzQG+TR1A1WnNt+vBhp
MsuFTUjiagUCMXOEWwfNb+iV4N23Vs6RMJYrrIRMhSFYUxPBO50CKvBdlg0rDa0t
ypYix6t+vsoLg3KpE+Wgy2iWduirwoKUChaI1bP4q5tXt99vSJpCllrbS13aQ9fh
1BGvU66JR3Jc4qt6Oi+l8WwrXZHAf2F/zwBXSN66XHEjv5kMlOw9lJnyiKLzu72o
q0C1uOklSX7rO3D2ExVaplAB6a4bTiRvB2jj+Oc144f7NShHDP6cmu0Ubee5+LdT
nM32go11iD3Gp2iQ9NWk7sQFyi12daR3YlE85bWhbn3m2SwLKRK5z9dGIojjbpPp
mxViH15gwdBuV2+puOyw9xtQSoy8qoQfa9ep2FOzW5Ea65GQ4aRb7OtObXcp/fDh
wY/w9ebO8me0hxKizPosfazErKniARunlUprKERYo7BJB1IXG+Vs+nvMXyqdy4Q8
ApM3JMysRstus+j/eMPuqCVNF/uXG6kWs/OfxXeZQwmXYY6pKeXdU1XCUFShWbfB
XFGTW9gCKFx07W6g8LRkM7P+y/ZTVGN9yhE+JUkDYVhbvywbAVsmKooXPTlBmDeF
Y7GpxPsT3nTrh1OTtsVNyzV6UrqsbZ4EqUEOdc9OH+8ZKkTo+AOupotWjsp/UQGy
IJG9rnh54x6FiVBl6V9GLgoWB3SFay9CTcZXVLej22wL3/FyBzZx2D7ynl3cgsg+
c8cDM3umzHQD+lbspMeWFlo7BgfaRWL9DnIBGScLWo5WNEajfN9nMV70NKH5ezDL
IPGrebJvaO4dSg6Ct9qujvVtdWa+SJ3KOj0QC5FO3CWPJN9nKsP3P/58K2x0So6I
uihFje5IyxMpfxWKkaS3iQ8cG8VtCD/XDPAgvItnu1R6h6/tRdsWDQkHkbuej+UH
10u6Ni+33LrJYbB7UjM7oGYcF4rqfp+CM3Ftk18Mq0zhJwSWtdI+aO4Q1CDedEgl
PeBuUnuDW4VuYqb5jZ6iJ8ujfOJ/GlAL/taa/8js5GYB2rEaObJ3hH4JvMLia0RI
Dnd2EIWIeHhQM121iPevJYB9lIU1AuPS3TFBcqvrT0KC3WtMBsU2cvMIyaO16NN5
Jcxf+9dcnC4DcbOsq2b5wDVc/wtJmlETTqDSAqtQ91P/ysh0ewMgLtwpJxUWVmrQ
TXjelyhRvfA+ia5xR2O7P61DkVrilfsQVFXsE8CVywBs2/yS6x74pvT/vMePsKW5
5F7THrgYTuSSPa0tDdJlzc4AYGPBgRCNrpaqoG84+9+WGUZtyTmBskCjZnz1IL4O
5hiyV0NLrZ65QGkup2jjYPFuJw2p1annESg8puJug+BaoW4/iv3ykJX966LgDYty
S903yidUtniEBbx+HL+1LjBUdN8yYEZmKtzZF86VQDff+niO54AP7WTbX7rMh1ta
d+DugPhV15Mt29p4vXwDda5JpKV2Gr1wmgGzbS0iqKp4TU4fZ+OQfItkIBN0txxP
NOcYAqRVkD7fYF9/aE5sKQ4ws+TBvnRmDhWvocWI3uM9YS3Eu2btIWaCsXwlyJ0L
ymnXNf0MJMN12rU4k9BWl9GE8nK/pmdYIrUQw0KsGS/l8iZm9sVg6X6GxhF1unBT
DuRJKYfLdzVFeaL1MmRs1JlAHR1Y1dClHX5oVzFKm6eJCB7t5vGh8kZ9vF2N6v+o
xMD9FNWA4xMScwpfDQhxpcy4WGT1wB4TcBvhzF2tlNkI3iAfKru8exLwwM5dPguS
oleIqBYm42NaVSrV6q3rhCgzZPhVloZ8E4kz0lfstw7P3toPnH2xbmy1qSy2lpT+
o2IXMVbPxRsazI2Tm67nJdqot9lIKiY50+LDglkSqUyyaf6MA5/TtBcnHTJhvRX3
bikqF1lvBW13GcdvxC+GfsJwbd/dftVdbzZJoWdmfCKYUT6NCmV715AcZmSkFN7J
wgOjBBnP3zfUd4Sk6pa2upPdCKTbx3jBEfg5iU8HvKzzylgEmCvNjK5Fx2QzuIf/
1RPOc7bsOoWc/8+mmwnV0Gbo9/j7gVHlb8JYqZNqUHkjrH5w6e9WcGhpeWwOk5cv
DvemO0NdwgYDARG27hUQqtflhGHsiA9BnwJLl7xozGU3sXhD2+QyV5RtYnwOfNBz
2NnW2gK8aoWUx+NavRT16xQA8XBtr5wV2Cv3XysCbyfCv6Rg11L5CeUZulzx3eKX
u66NpKDlSQIHjp94R7mbtNkMVAsD80wU5ensZm5LmL/JzAqUh/tcwMStkCpG62xc
lqAeOnNKMKy3cGvNOlpw9+x6Gkd6lEEg5/gWJjWHv6h+lr17RSFs5byJltDZgcYp
dW2dhDmrfz41nwaRa2oqP3Ud74fky0bi/8rmVTEGIAQ5ii0IHdnpxfNANgNk11Zs
pfU2koyCxHq1GQnjd3GRZrHhhj8JdcyM8UdyFf4PgQaOqTN0y9Vrd8XAxMciWU09
2UJ75ZDvEwNGgf5hRf3+ueohbG8Et75gZpA5dU87wjGaSDdY+fwMlBpMoBeJNDAH
n2mf75VJxh/yf3rqd684luSJHhLi43DiHXv/hF/DfRkZcrioK+2odALKID8f0hhW
WwLlifRDysqegXTGZ7b5y4lv9jICbeglNKVBDhULNtQuIsmGnt0ZIMcFsInGEWqN
CrbpGoSZ+ej/n3Pqcoy5csq5f4ncv5VBvHaC9GAZSk19hxSHbHPy9kyJviXXeB2I
CpPTLmWxBzyt/t/Yc/sEZiRHAUzJtA9GNXpyITZNUUXFYwQWQnxkFoQhwonGInMI
txGYATgRddaBYIRGNj4WxfgE4Jt4hzmCwIJEE9VoaUHlJYdlSA3ywTpjyG/skymS
eec/NfVJq5wWNT9nRiuklGyRvktR66Flk13VWy8RamneBBT2qBEDV4ujSDq8DGGi
sdNBSUK4cVMJEUC135tgWgU9t01b09dvUoPs2v1UV7WndLxt3WfzmFnvzcIRwd8/
S47HNBlqI3NrZlpyDkX1bOb6ybnrAT672uJgjZv+6nBPqywvBk2Vd+ZlxFr48FjQ
ZHP2muP1iVhFKl2d/iVq3Q4UFwiX5yJme0yPz+1F0vLJpgY4jEwmTiBvo2bBhzs7
zm4OQo2u+/LbUR08p59+a4pxyeyOkaBqD4se8VprGv6wq8kyqpME458cyjcSZVmR
RDnnaWFwsrkYRjPx+D1i6s0TDsf7AzrYER4z+OQnmpRySG4bBiIdV28a498I0107
b+okO62eUyW68xSvPpyg2B/dCinNwT/C8T7I8ZXnwosSQ63OERDFlCS2cqtWczU6
eOv59p2SYSq7X+D1EthkLPRGsrWhfsf496OWZMx9vTLcaA+312e2Lm5YDWhKjXPw
xl4nUbDjDGNsndPmV5uoIc1iU8K3lYEPcqK6JojoNN1U0cT8+VNdC0MXBVax87+e
OHy0biHu5Ogk8gHpcA9x1kuj2g3Z3j3p1sMU623Ge+eniOtd0PRc3zFuWW1CRGdI
O0SCbv6GWfG/zQw51NE1SEWCx5d0h64MXI8EcTmA4F0ksMHVI/PmnPt8UBEBxHT+
4uqxg4i3DiRWx6HmXd85eMtDVy54t2jqdZawUZCAPpHrgJ6+2Q3JwV7iiJu6jmOK
JReGrRLcet9l5iLhhh2l7UK0PzEGsFO4awk8hbLK+n9FYAhc4zOnRYwYFxAZ2C02
0lUwoe9bSRPbwnLrFwJJO9FcvIKhrPwrdfGTWJfI+PuS4MFT03/hQqBYlwYaAI+h
O9bcMjEVmkmFv2pwLtPotCPDued9kni9j+UTIQM3PLOQRqz3W7t4oRnb6eDIcE/9
tltc9kFSCQFeYh6kSlx57CmvXB7F+n3pz1iqRbGyzs3B7JQiBoeRBE8VLEdmq8Xx
+nWUIO4kRrSJ1Y7SIP27NcV+ETTGBsOg0pDeo0Mn/rJGPbWCrwq8BshNdHxd6hdZ
IOD2Zx33vFhLzz6y2YL7duzfRWgWvFs6wlZBeA6cSjbvakKYHjGtWrQhT5ICT7jh
QQA0nLOI9vXk70ncGhFOKp28i+NEe2BinGJiWbqhaQScnMt8KsdWrEQ4NrQzzwG8
ZL/m7rw3Ot8xX3OfTkjjvM3lGkai7tOTG93Qbc39NqbqqHHrsoZ0ENszKPO0liXv
42s/rWcnPvfEVMtklLnYVP2DxRkI24TaC1+urdJsW3LmyEU+MVhdZWcK6hNRnm7V
G3QtZxT3xzfKVHCTgJ9BFtKfemTndS8J++Q8x0V9Zg/0FQ7mHWSqCIh15uCF/M+c
sz9YfRcVbLIGgc0B/hh2kT0NEI1IGffBUFvQj5UVTbjc4IkIHpfhwSDLg7boq7FN
cIIv4bX5WDwKJJbTMXtupWNgIS9SybkKcBsHuozWaHVblZpW34mt9iK2Ztfxy16n
4FHufMw5EZaHM8CeT6N+ZsRlf4RNEoSmuC0dirwgsNn68rVmZujF2CRWEcnMsWJt
k8zr4nEXeHuWDPS6B8nfVePf6kWmwic1oitfeonwu6amlorZZdqdEC9Bjyn/KFnZ
gFdJD4WbI2i0i/bWLDS3WITIJ8eZ60znDQoBiGwFTppVYyqjLyG+xVCBlT8zf+ac
lToOKQnIiECSv/m0Phq7e3cySbH8EQgHNtohOyKd3vuygxmVc9HH8WMEkGYDwecg
4wSA9oNRHWL5DWLhL01+NN7K+5WIqC/jTR4e3KSBslwEST5hj8/zvcWUOblcjukg
s+6NKDpj/rE8tJdAFZmbWS4+0bQpK/econHcxkiW6B5d2wu67rlhxWFg0i4Qxfe+
xfvr6satFR4KRZZTJhMGW+f8yOufRt27Q4e9kQczP58MLcWUEKHvio2GDHzeyOdW
B9q5U4EnRUaBdmZ1q1LqhYpg8mnVal5l2sitZnhkUHxjP1TjItgba6t/ardVHuax
1TaxI66WiiXL2+JDmO7oF6xDCk9g3/4rcIjCNQYviO9jGtgW51fy1qHmgZBVbuFP
crS1iQHba5vI4eeLwz6kHIXzPRT4grqoEAwUOL4VTGN7jT8c0vuRLPzwyujhcLq7
nHRKGONBK8r1LXF4YWK9SNlNKIjOvibJ7gJ8kdUXSr5JLnwC1qGKKmbFzs+UHBAw
sQWUMH45oPa7Z1z7DI6s+mp1tsaFpamn4fu/VqTo+bsDMuSIWyMsRfgppJrRZREt
VhKlXZpMNcJHAdN+gapNWZn5ps45sPovpiTfqVbkucT1/10TrWnw5Isr4pPAX9of
db+DPb0/6VxRsQpY5Z8J1wC3pIRQG7ucRyzAu61XU2dDksxPbPKt/bSzv//pot7b
+NSXp2RispG1z9qXKCav0gjrV8GNxr0Nw1Dzi2edOlMiynwwrs4j5/1Q7TvcUDoq
g5q7JUkFK/4FUH7n8GfVZRfkxcAUH5Tie5k7qzWN31gSliv2kZoMSzHkUsFfZTxk
rzV8YgO50q/2iFywZaVK6TefI8CzAJLB9WN0N8Nt7fIjtcCvc4aXFALfXcGEIzYP
oR5WD34JEHcuM7gcKeIEPYi/IEm3+mfCsUNlVa8HYAu8I2KgFIaRtsobUDDTU7Bt
2FpVG4o8/+JXImbPOBBnQHDLIGFQuqtrhCFl9oovKier+bKG4llo6xmT6GBhwecB
fylQNk64GJ+n6nWYtcG1mPmDLWuV2VGFwINjvRB2xk/ZTI95tR2U7DDTrQr1/ia2
ZUjP6gHUA/iQSEsPx/tAvQne+MWo7Cw6WT21xsPqJlYEJW+CA7/JoVgccSsshdZy
+O/eS5fBPZfuwDK4ooExfnUg+k9TBHitpplMu/dtndU+drrgFJpAzf9n5+lVrBo3
I45C9KwCD7Y81SQMf234R0QPC4EPmQPFm6hG7VJqvWL93hmG0uXtVIcMaiwUakhw
U/csEYCv5VNy7kGI2iCJG5buMbrIYR49ZzPHMdIdD0wb44Sv5WH9pwcsEY0sJ/jk
+hCeH0UVGI7JoXI3RfEAnGzbTbn2s6oWqUs+kAD2dq04R12DyPwnyXp3tP1iZkiU
/y1rfXkpctXqJYW4wTORqGyxF5zqbTBNxDRzkoPnB19r4peSyb1htMGvxZh2rW7g
X+lQN50A3bAzIjVwzUMpdM5rzNUK0Ia9xp2dQAze/DQltoURNIZuuF2NFwcqIuGe
a0leZiHt1JFPFJmCBCS8qvK0TtCQH7ve+3y5u4xbRKsvQuSOw8PZkLMaKQZ3IN9H
g+DL21+9LjctbvK2qm+LhuHnQ7KpS6ZjVjcZB+De9Fn0qXR2PabdhCj34d2u/ZJY
108vzfOg3tUNOxZT8EoIv0iF07hZ5db77pcHoSgCPqNF4mLbGp1aNucnwvv2DVh5
Zvpw50gKPFoJfveQCV6QnVTzP/XXR40OsijFNP43DT0rVdbcJq4OxG2KxyUFOdCX
DppjGP48zE/SecX/1L58/CnRvCk5p4eOSQ2+r/qQbGtkHLeTas3eX+mUX1v+kHmh
QditkmxcajOJlhXUkbUjsi/1et3pozIwnlvROdEgy2vZPKv3YykITTxzTw0CXZsg
hIwqS6+am6uwYdRziL7mUJhoYMXBZ4ZfK2tTQpmfQ+bRfast35+x5EL3lM58DlYy
VAmTKCOAntI7nJZ3sqZEhuXT61O2a0IK41rQ03HiTEszCEdUFwqO2C/5cb1D7VBX
jDaIY7Gb/MXEZnkQVEY0adisDISD1oNxfxhkuNiEXpwAPtKfC81HlyY/MWPNkNuE
QtMNSoacQdrBBjMyULIdKyahR0L7BiWZi7OXH71blrQhv4DEcOTWDB852w9Bmyb7
5hoxIZXvIwTWGhtL/kXzwoNdEuo5DRSd8qcqQ2YWb0ZGdZ2wDb7U8heFD6NGNJzO
qWJU56AloJU0NQhLmcSrVSBkiDycxnm8xsQbDlRCk0w3akUYIvBM2q/DWWN+0OQq
hNHfh0U6Wsd2jVm1/F9sj5M3Cnw71pzdp1z31ecOnHu38uLLvqWVl614j6/ygk/l
jeU2mQzEiyhZ4ioJJcf/gm6hYWQvYHpDkwYbfRatW5sQQhnAf4jCRSv6F05mDk7J
Skv/OKHcKPBMT/UiTHITPW0+JVcA4TzbWj9ezXNOYyACtChF93zs3m0ebYxOuD8/
5SsOVv8+r2bG2/3i/gLobYiKJnI2rizuf3jNKSrdJWPGoTMTUU5/ETRs6l8cULBr
i0ziQbWsvasX9jzP43v2JFCa+3fj/pOzlgjqSRuu54Ugs/UVkIoB5Vg1swXFEI+p
/jUJ0+NoOcp3QWX4CVEN0yWrRZDd1ToBok7mwe21NJ3p+5P3Q+A07w8J4lvA+x2D
sCsIzKn85PRoiHAJWCCq93zzUc1JzMJDR71T8hhNrI9NA386qO1y+teXMjV7lTIc
duH9eZySZKFCbor03450D1P30UO3f5o7ER0bsMpXqJKEXtyttTgZQoq0M4bc0yjb
pjvC2il8O+1efyaQpJu70pEPuDo1d9H10Lqt4lCBYYswOtXVBdVawy7ioMV4b2JI
OOOV8PMs/9HUQk1EL9ZPwUZmiYfaFlC9znedGz8tYuyHLudNmdVELingSomcsjdd
SSitINwrz/n1vDZA4vJF/fjn1KeVO1gTO+gf0VshmZ6Pxwcropc+PtZAS6I3FrYr
Wm0U9PJiVyXdZ5QJFRI2BBPntCAjBW9cwdPNQVaZa8/nxAgpDknnjvE1TU3Ij2VD
FRg1RWjs5P2U/jEEPZTQyMV6tlBzuB0wnb/nKb+mmcae3pdJtqR3PRAhdAmlfc0C
C4ZZbweK3S6ZWDvin0epMNOW4y/6nF1yzc1qe1gVbs22J7Q1n83etZI9A6oGkSnf
qP8FOsXa5FzdMI4ks0ELfl12mPAaDE7hXqwk2+MByl7xJrHoOqH4zLwn8DSragj4
QT8UJhpseBqc9AtLtdJDCaewbGRGbz295wDTa/Vzen0WZ7lvcLJU+baRDryqaoRf
PCj4mYd0DeYtgc4znNO7XiZIcsvEuxYUHcqHGppcXIARsUzxDZbPckLPH89QousH
CO3v9IWI7V7NjSVSPs4iyTr+uFnYzKQ6tF53J6t27fzLcmyvdnwlxNhgvdcDU+GH
K8R2U/2h5ssAL5JAVehxdhY1GN2BWG1P2UiMmBB/F8ArY5Bnp9aVIjHHIn0/xBkn
bELnfA51Uj6JfjQ0XUePEbT5g3YRPOTWVjgTh4aVnQbgIAiMPZHcArVy5bNBTWbG
i9dooXrzrhjqgjxeFa7ix385wl+WsOh8PbrofzXsgzvmM1Hm+h63w/XQTeW+DWZi
z8fuT8pYmBJVKvFtc49HFmSDo/X4LSKv4W5jBH+nzYl9SRkngCnGk1tWqdCPNraz
uPIXO8eQCHVjxytuAHUaHOgItbRhZ3dUFPtw0ExT9lbkYSjS5hI4K8VF5mNwN22L
qyUjxyCfb20p1D14w9sa/uMxuscLmywJanOQEcAoEIo8hPptvQYAsHONdBzjEa2u
xaJIoM4mBUhiljwaKFm8kggz9KFeJo6eyToUyBWvFXJ2YWpWMZ1pt78+IzSpVwqo
ovIyhacA6Yd9+mcOt+zNkqwGiVKAOSflavFAuMWey3l42pKLj3nbdUkmclzvDulY
nxC8QNzlj0D+SdgIQ7387X/EHbHSe7usT3M7KaOeSQzh/LV2QvELuji3D5OA4AFJ
SKXQxm9FeN0ST7BcTfAY+sBaveVsXinJtdZvq5OAYTVrBLpSYix0EDeegRsg/n2f
ylvsaKbi83guqDxgTQT7gW6CkEuQ2EaNaRedQ7I3kMnfClFpqVLg1c4RRZCz+ixl
EjH2KxwzeUtHZA9tt72924FnIusuQ1apknRt7xq/4H7BmMQtjVRlKSP6ihWDtjPF
gXFPaOMCtk07Vjul5DIFSngeYlku6ETbriE+m+XXa15bNpds/ZoTHrseScVPdysj
nc0R9bKDqU0XRDii8gRh+hDkGGMrrvOx0lX0vO+ZtY3nTF0c8ZjC6iiU8U9K0KyY
bWatQUnjNLuQCDNALSli8R9E0DYJWMU1eQsnlCFY2k9tDfLoS/0OG9feHjARQNjm
LeS5YqbBKAWhZ5fxikuYrS4lDRMIwvGK4zbIOX3ua0FlL1z8aHE7PJWZ4BWAO+D+
r0QNMYr/2N41loWgW/G7aoCc2VCFZX4rhKz+/BtcOvJy0LrHB4J4VKfYcMsKSdqp
S7peE4fQvpcJIliOOTyP2WHwGdOgYjHtErzukE6GJ5ZyTSpblMOozncX7js3GABT
HF+Aa6b0QQRkQ5+n9rOmhDbZ+vNrr91ZKgNp8CjJQC1ilTzd14t1QEoDndn97BPd
v6tPtZS8X7GIOdIpL+FCzNrGgEi7JaoES08HvtFUVSBVyf0GaGeA3MVSpLw7i8ET
0g+HlUpQJ686+VCGfTWkmkmn/nIGFmXZVaagEYnEovXKUDUDw6brpGHmFTzgatHO
lSXUy251oAJOkOudi1KVrRbNO+B0B5EybAcMrOhJbhuKQqhJSxyYladsui4rDbsD
vfJ1s5t5HSYjG26JcRwWmv7vmnauziY+HGzyWPfrBpBdLW0W0+Y2MSQcgHTP2dKX
DFLG8eq2XMD3qvrw2ZJ1NQTATQp6Gymv1mogwt3XtXvkN9W3pgPfCDgS6qgAKSlB
++Dd/s0Q1noxHq7ku1eORQ5zZi7PruGXYvFXVH0AmuIip7pmFmoyp7EuaNPa+du9
TQv+x/QS2Rc6UHXEigOAsisl6estzZYvzIym6u6WF/LZcYTorSjaPXuqdm6nenhS
MBGUzs4ksCqp+SoeHjjsVE9l9v5eWuZrS0A553cFX6yDyb469tVpM6BjFSx6LRve
Gb2DsrvdwJ9/6mGbY0icdRJzgVa5saH1KqcZOQy93bp892rgc04eMocjbzO3o2An
uXsHvVWxWqMF/OFXfCXobOJFY+b3H4AnTBA+1csEx2nKIEI/09MlGGbPWgGLb0zP
P3Hy4kZ5Y0tYYWQLlH7m+7r5iGJI1UsOUlFBEAd+fDD+eFSTkRdk/tlqLRG6gAfV
ADA/tYzNllg1DiALr4p0R2cDU5QgwfjMCMCgcdu3AEFtf+nVS65Qy3Puzg4TDsux
GLsgPDRa2Xu7Bp5hKlud5HBTsW5b6xEtRv4cUyaaRI/qmW6aW9qTcOC8c1HSWtv9
2jTV/F64pvJg7KD4LWRMi5EOSoM5IMmMWNV6faIio/q8Y4Vc2hWJ+zSLjtrmnqgd
sJWupnP+e/Qjt1BCatVT8ZzR9xXQeIKT4cz5tTLTTQ9dT+60fofhs6IN83prkqCW
XK9sciVJ5Xrk1y8O3Nj82F0C37ZiL7lDh0rdGmDlENK5hDngN5I9rjdMh1LNLcTx
wN/mABFpQyLoUS03fewMAR67juS6I0uHHsDgKn7z3E25vsTlgJjgS3fGTdy4ZXgI
hQwiZowTyKIKcahMaSMFN0z5slTs2+QfOqmm3IOZfWJnXo+rKxFvBY77v6NWSTB7
R8VVdqL3RLoriz3WzWh8Z34BhWsmhwrHSU5vlU169le8aTI1nKwK32Qh59xxRZmd
8PoTY5u2sAMplVhb3/8pYYcPdzj1IS5uUiAT7BQKEhWHn1PqbHaGUEk0fsoMEIAn
2n/Nvq6J7IButmSdON+geNbCqmG6VyaqRu9woqlovGzU8/jQyuaBsyf2V/KLMjfk
2TEakou3z1f9mKOq3qIQMvszc+6r5EZw2JclTyPNZV8nDfBh2fDoOzHVY9PAsOEK
427CZmjYSVQirnqd5ePJgxpDdacV4CpYRWja5EeMNGL8hi0D56UUBYFqB4Rb2EWi
wqCgWe4a43DmMI5Kwk0qLqdMbsYm01FSKzQ01ArjaXkvFasYhiZh0bZrD3e56jTq
TqEDhEm6PLErDXV/wrGqv6eXlCwKMEfTMF02quXOelyXortLIDlFOTDmN7fqLSSH
/SgwiTw908jdIOWS/cK+STCpEOt/dLbDyZb0T9e5VsfSABVlvHyCUbTsR119p5K/
D2TEPrciX7P9FiXtWVEVNK7OeoVne44Omri4jF9yi2x3bQFMfQutSBe5DG23/Mn7
aRBs+RNnKAR+9uH5aVVBdqpi9Suvl/wq/QJKf8eCozerR4YJwoGN+3cXSfIENodp
5OvjU/TinsGqn1rilzHO+XBxEJ369fpBE9XuxBnRVKGx5/uaYrYd02p/OWWSf/l+
zdm2ou205ZbJIPtncakaPQeMo+nOR7oImJQSRUN/x01HlIBv9OCU2d3T9IXqMNbp
dE7youPtqpgp3DSJgWoX+h3oHi/f0O+/LrpoCM9/k9TNY+J9PgZFgkGtczocFg10
EqbA+kgSNzVEpTHavz6w0j37P9EBcqu8ULEbuINM8mPY+JLlkVPVMpuYGqBEEv7V
389oOT6styM8JW27r9AvMxuMCyELhZHioztq25KHr4yepOHIgMcJlbSIACUPBk0E
TCAWNMkWj+9Kxpm6V4F5EEcn0VH9d+TM4OpCqOslj7voFpMtQNUZzLDtDke4jrVD
ewx6w0ugFWpkQRtv77CyA7Q9riGQi2UaD1NM37DMK0KbHq1IUvcU0CCo9wkZYOlp
Y+81JPPgGIA9D3uqvkFQqADDjtFugty/OF4m3pS4+TIR+nz+KVHuilLNq3RTzDuW
CO6OQMfsX/7efOsrLbVv1VFVQ/nd96l+UUbaV7MXVQqzf3SuBiq6x6fT9CevuspR
87UoOKJWTA0uqhJpICivbS31ITzx2MiWttzB/dJQG+TsrTMQhKT3fU9f3iYvrjrP
l6b85NK/T1t7QlkOAvA5lWryecrWZhRvh8o8V34QQNtvQM5RQn9WT4cZB9Qy694p
wG9Un1lKAkWmAiTd+XMjBGuJkaVpJx+PNqPwkvsRc981HnIxqKLw/ZxGxF988NXd
WguazAPCpJVdIzBs0Pjd+E1niAMUh7nLjKYlGoE90EZfCoUf4aYq8UcwAXTRwi9y
sqR1+s0yJ0hsWvAfd4i0vTcHd7Y2H2B6mWNFH0ErpFod37FDEPVBOrHB7R8rfj2P
PSjRkT4yI+m7C38ngNcLraCDTt3eykWsB7JDRtu5NwoEnDqqo4VOIW1Zo1mNYyVU
Mo7gOXZwEJ/KBfhwLwfxTy2F+ariRpuvqiAFVaQ0wYO/B7W/ec/39wX3vZVmbkyF
nXAniRzLECJ0+oqepWrcJ6mtFkvRZkuxT22GauxQpQUbsywFSeOlhnfEaAo/XvEp
S1xVZWcIdAhHyvDOHwClb66EZGoHRteGwzwGPfO1ReyFIti3swVe1uXnT+qkqoRg
Y1uK31ddlffKqUo8S929GdFm4ANZ1Kf0F3EnsQVr3v8ey2Hu89TbYizmiwSQW8Ia
dEcLXt3/oz/tWkY7nCotg0Dq3pppJr0DlP4BRR2cDfdhtt5Demkl3OEWsiwF9HSu
xfBGuwz52LOlhecy3leAXJ02XFVZ2LbvvXAyzD07K6vRSLc9mkGQUgIRbH0OuN+A
2wLm3zhZP9JkcGg6+GvpnYf0FYDGbr6Aq2UkmoCDF1a/uNHii9HufBdkoAm2BEWb
sGQ6GJsgGtLlx46707sPFmJGSff2jpxjC9Exvr2l49R3BDKUK1UJ2hylNBB61l8U
jdzwf+h5RGV8rlfVjpoalkJ6MRDYZDijgrEEn+uLbqbx36jrX/AlZo+b8S9SI87U
l6Sh43c6aUtJgrOQJh6HxrRW4KD1JFkmKLESw/+r0ysYu8QQzgjuRX9mBrLSARb6
FaKwyhh57fw4/uQQi2QaNAZpN7FVtod/OlD2UDwz04/yIwAjwN5bowCA/c7D7G0W
YWsbQUiHxR8kC5Pa860sPSgqGB/uD7K1sH+cBpHAtHgGX7whlG1CYlWB8Lcmlt6y
S5S/sHuH69ZpSQq5Hf8rsmLki8R1dZoX/BmZ9n2pMBLcmvNLQaSe1RCj/L6Dgnt3
qBUdgqzCn0wxOhnpM/SxFdRYcP80GSS/Cxu3dDelu2sfMz/KTpHfbAFZN8aPKDyC
EBMbskENLW2OZu7GYeMyiUsk8KwQGzx8zteWKyyN6ezCTSQun1Bbf/gBqVvpdZFd
b0zxR4CX9D2QPeLuyA8ciYTDG8D+2589q4QV6WwCPac0Ls45f889h78y47p1sray
3YL3uuCjzNwjN19PqsEwCr6En629LIV3t8htTp5Ml14mU6eV5j/K1yVHjgtvoc68
rISN+4vbR7q7wDzjtQH7uQPGX7N16RgAfkgfISnPFFM/g+ybrD4GaktZXRwACC95
zG0OvA0h8X5woNu0JYpZjEp7xAnYp0L5K5SpccLISIvNZNquAJ3ayJYgPZE8Cq7Y
5RujxpLZg+0rKcjTq1RQbG9OpxJzk/lGsBhtIKd3Y/XNNjsSY8i8dMfxi2d99PXm
TJuloaNQKGLlYYl3ZlYP05R0dFROaPOFOaONHA/h9NJ+uQFcjDzieOxHJYTmCvGt
6HXw45OwLK2yQrPGRnkU4BBbqcOx9rG5gV9kIkRl6qaFPgNh41Aqg6ASQgObJjmB
vJnpFWb0+NYH+jSuiHdBb3WnB2egJJhB+iN5LiSt8iSNQ49LE6iQoYtUlDqtZybH
qVq32C2l4ya0yOd9LQal1rcT8ljwvSjA310X9ZSiMH75XuXX3PQNpAo7uzjlBrGX
QkbzP8Pzc8j6CrhrMPIUmiaY1QS740TS6YuwgUTAG7YBkCoNmvNnIQ+2Jib961IK
qsvQPWmjFesAUFyXGfASgF5Y7OHurBGBjamMSOCGwrmksXyEjUjVPxH/pEKlNGyU
uLo1EmL9ZlDfy7NZ3ZJoTLSkeJhAfY9H8iMcWzNJzzGkgmBvlBZSAGbkLpg4VeIL
5PsLPkWHfFAA6ExXlXyKpCfnEl4qUX/mrsPcV+gLdWSOq4dn9Le/GGC/GMta71F2
/QT5v4qnnYpArucXvwCRKtGM3+RxYRYw18wBQyiguywOMf0ufdnEmPc8f2SUy/9J
epKorCvGl8fUcZjZ23+wCAstkKxbCSPnVeJ/2eYXvQHabtvTU+SLcyvQmJORq410
CMS2TBXhgT0wLb6kFlRwOQX13/KKsGmegyijQbiL3m43EEV/nPUrdpUPZjDPJrQH
LVsnS0MYRLCT4ielrkVefMfxANCV2ydAsdqaS2VIQwINqbejCfakX6t9gwIzUnSU
ABbMCvrjWMH2gvpjwd153G6DDctXYMghub2ZE6nGC+TUiDaY9LYnzf6MFk2xoQnp
qr12IVG7/M+hLewTz5jmjz37wMTDnNjJd7nEXbf08amqpvMVC4e/2TSBX5BRynM+
ZHPZA2j6/zJmGFBiOQBX+BtCecKDTIkDMw5wG96iEGRzFmpe7hcZtD3hhTCxagPo
az1Rh+cio7991OOwyjWBduI2UxhUlMaXAUvkk1HqpnudLMm6YiJ3VrtP7Mwl8QD6
7mXy3xgqw58qzLiUPCMYwK7IimgpW12jNve1H75bdFbPvmP++e8WpODwOZ9z/vOo
NtkvyCOCHL1jjG1JPbRCSBziFSANXuKJl214eMu0dHXb8nL0rTOcMVQwVOVv2Jba
YmKqNs24ExnwvgDMXyUI0Mr2CI//RN7Z1/RoDZY15wca8+FMGR8CJp6Sr6swq4HZ
nzJyUzdAL/mX05sLpNM6IX7H916Lxb+gKMCVfrlOdLF0+RROgVtNLBcm59bJy39Z
RGjrL5C67dw9FxLWzyLW3hCDji2rgiX5784AI2qeywkk8lNeAbag+yaRyrJ8fgct
uEuhuxx0AtVYQy0k/ao6ylUVq5+yXF2XZWcqE1Loa3gAQKaq7YDea0F5KTdFJWIy
VsNtdBknT/gUMsHt5RSS9Km9yyRIuDuBogCL6saXRIMf+/r+eyCHHOCRy9oXTgD4
QnS2bR0nUoYp6/Dj34lw4YJQQkipbO/bpNOrhdoCA7c1dXhRACfHN70lA/97tug9
nG797aszoHawb/SAF9wOmkbCJMae1/3wt9pS/uyRa9K6tVpt2COQ61ls0vdMx7KN
6VuE397KvNxDOfU4cmNaYrdOEyABgiCP4anI8Q2+WIO/yBq5efioTUEC+cHpMEB2
yAXaJdRUDAVGDJSiBGEpquzwePFRkFkE+YkJG0F/08MLojSv3xn/mbTTF4lkyY0F
DwU9/82FjH1QdgRQ9w+cfxg+zgw2eiCcUv4bmWuZi8ZIOdVPdYloFrqPGVm5nmOG
ZsRWUg3pY25yJdCZlLfStYEu/jEfrSHFu+T0m6BaF3Mrn9v+tX+uo2kL879nsESM
L2x4D9YRE1sT+u1arvHL+TnGdScLDO34g7V3XJhK1BIq1SkTTDhHxWnEElX0rcY1
BlCENaNbNGKPQhPuVyb0nwmlN8zyEEftI+LBwCLA9tuUTd7GxE/R2asR6blp+PZ/
/VAS8YxGyLQUwBWqpNK8tCFHSwortHkQDy7BUbtXfxwMlcfa1zN466oOLsfVVgcx
vYLTIoEVsyeO87Nzx1Ry7g9H+fton6O3wEcsYmrPdDUQ+aWu1TwCLoDEjHld3oeT
3T2A4e2wHSXb3qDWPuHqBoznBIGZilyJNIR96DWoCgrzqy0KNIO/S2xwn4Sv2NCm
t+idIMhL4kCUHR8EH5TMvoFthIro2wnVVaklilbNaQHP3GQMPqX2rjRxejK03zxh
wXenxSmJwtCS+gaTfVhzzAsha2CHg1G9fM9Do1iil8gPF56EsJ8DyELGAsPUErBS
vhmsqT+CBs0E0FE5LH8tCyyBe+mTWqaAJWr8DWNNHAJ4JNXYUjS1LE6Uy6vEFsYf
hD610RFTY/AMUznR8SNIUqRGBO1iFDyF8KKiKGzcc8qyNEk8ujub0UJZyV+LlmXA
AIdX4qv8AjHO+u254FO1FDbTETMhy7eE5etkjASefHbV0c2a+ALk+etE0Su50FhZ
p6iqVUtMkMXyZ4RxWUz4d2fTWH04k13TqMU0p1DlYVDOCafBl1NOR751CDyI7SNZ
O4J6ZRx1UFdY9ckTAS4fPhA0U/oySyu6fHNVoLZQLA+mTbUMg8yxRvjQJCZpwtgJ
6kawiRc1etKjtba+2GycF4VAdCIJP1XYRWAhz9g2sF4XLdN+yJtdpXeA35mcQmEr
FsCfiMJGp6q+81d6MHpF5xIzEoz5ZLywEreCfuj9XbpPTaT1+X9oAJgRKZfRdFRz
oNsEh+vG2p4+eW7txaLFDhucLDvUkwwmxfFTcUsx0GLODHVxPyEY7tbAULhBT/tT
uwO2n3pzJ02541O/j9C3Yzxq5ZTXhYKqxUTlB1NlHI2xeshzfGlvqv+WJf4zGR80
WvxBD29NNbHP6Y/AUSsheLnictes0Jvs8sjG2vgbhh+8LZkfs7HQMVTMIuBEOIod
G1IwlNLV5qEDUY7iuK24+0kJcO6EgKYtk0AyMC5Jt7+a/X5PMq/HJriW+Lmm5ZZN
+LbwOMcGVv4tTl50e1SwMiec73vys6Y6igMYbi9Xv4pO79xD2DjzyBKVROThB3LP
sbZCq+vr2WKcOggEGRiMdceVEPZ8KFZTZaaG3unsIQN0p9GHjFOtLnTk2A/n2vmr
+gdpOpWjXfJjMsuzrq73z+KuB+jgL0KM8w/jstJFpQbd7+ovMRY7dytHS6/4cLUE
82R/KCbQ15nrA6obZc/C9d2wc5ZMjOBCGmvjaSaaHV0YDTYVNsgMqWssPwirOiMN
gkW9YrCRgkd+A48K8YdTIcGQQr6e5wMJhQWBBkrisOkF0+NZPOIRWSVbKPSLJL+x
5PMqolCPUL/x/7cG2P3Dh5LPO5MbtJnDK/RAb+lDWaMOWicb3pMY/c8p5iW07155
tzjkGIH4CRRtpGnYa3BjTA/a3Y9HcJvYoSG3Kd7r76g5ptVY/C235evnTb0Tx8fk
4uxhbmCwXEO9t+87EWBfowlmQmdnZEcwVRo3CakRqb5n4rcMejlEJV9qIwVbSQrD
sluwbfqu+gpFZhGhQf17CFWZYdUjQkMsb5r3AvS6yi6NZNSlg9DTqpPDq4ziAZYy
8UcGyOF6JzfsflA6jhErZGjplUdixeU5ThFKfIbQ795YAjdCPDH2ljRwhcnVoHcH
EVqA+giwCrTM/gQ8+3wVI10fAoAHLPyD1/W7lxgU8EsT77DQ8zNYTFvkMeaIA1sx
TA35NrSco8LA5l6LjJtkusyPJXv7bGQUy+T3HPGUHegfXOO8RFZeXLZlUAH00yPy
jcZSUDgJf2lU7jFE0/4qdgz2ZEVtrF84UpTEIdlVhpt5k1sSHNwh+QzrSo6OgUZI
NXQTAVARr3yORAAmPYhjJqdzAyuO0UAuHoL1BQrCSymDloDZk1X0K6E/QMiXlfJS
qYrpH7wdDQsAnBWh0jp+ydH7iuE/yx7hrsqJGmxhpavmdwmEw/C6wj4ONFWFOrso
3eTFhO7M4O4qQD0iu8kSkPAXoKmmqQl7AERIgkDdaweP5tqpkt8gIC3nc/3uYRSY
nilgCN+E/TcWbh8gDfilHF/vRHolO3whwRIMRYDSsB5qqH72idtm/B4IJa4Wo4eZ
Rklq5uz8ch47kynF38xbtfYzl5AS1tp7tMHUCAJ3yvR3NfWNPQfMHIoepUI9y2m7
ozvRx1/1lbToCTixxJSPzzaRw9PhMostFvagObapUiaR7Srbg0tevhriqg7DKmnH
L0AsnmAztgzGHcaB5RhwKkyqlZew8pq2X7Pl5V/fHqXIsbRNjtwvGlIQTocPHQxy
v6AZhC1RbKlWLmUoRpT+2M2l+mxyTOcB977kwkW1ZLqntq+T5kjBa+obX6wVFEVS
ZcnBU2xz/5ZAy5SmE9WPdFrLWfXiyBHGoVf453DfhJTvu+NSe4tW5Ey4NdstCqVD
eC0Ks20arL/VDSysV4H0Xo9ScbId4HxlQVJ73TUf/0cpCfCy7VAb9bTvUVUXmk5X
g/VRXQDX5OH0nTjvCUD0eKtcSUPpIf/4W5guiwG44JW4CJJjDS90HfEdv2oeU6eT
BfkThPeOrJ6nyi3dISM2JttGkLNQ4GL6legxF08dZS3tk4m7BlouZ9HYdRhHsYfr
FY6H4GwSSmVMCE2Uj1bvAETRegkew2m31i904UXOdqt7SPSqhWmKdX8DGkaXUme1
AXSzEAugE2Y8jfcmoZ0yiYYDV4jS6pLxp4Tn9YVOPz4C/KQ8oQSU3Lo4Cx7S/dGu
+SL7u5xNmqjBwfMwGDLJ7pcG1yG+VWe1T/CbO+O8JY7JCMbmORRG3OFuOB9qq/gt
ILXtF51ItO06YGJhxXM1flcxDkIKxelChYezSI2dxIEAGmRAbJYhgWBp/niTb+QL
9FC3b1xGBSdi5g0uzDP9ZGkw5krAXyo+CH3/C6PS57wYGuxPBttKk7WCpmIqJl5d
rpvlFzwMTeYgLSWafI3l/OJN4NHNE5ErQ9F2tvE4cjZ9aR0rJNEfKsBxmOUe6kvm
BZvw4oqry35+Rer/uEnumEXZZtyH6HyZxTGxynpE2xclmJVn8J/9yqh1RE7JytyE
CZJpKv3Iuz/wAzLE/mDfeQqdie/N5UTF1kQIFyRSXdLBzJ+L4WHHaTB/o2L0WE/K
M7x67qlfJawX+8MdmAU/lKTs3IQtcVOCbrNvdkfomtxD7m0vskXjo1kcQz4Sk9Yr
VlFtJ0JgvxteyXhS0fWnPdAiSDM3vJ1OEwPAn6i4FGiA78zHK6mW2lnh17FSq0uv
iT/IwzGDMcKZEL7wX/SK7e7WF4c9/WPfcXSzK8c+Rfo28aUvQVgFeVjUg7xv/yef
pncMH/kAzWkyxWG+FCFsSLS9MgCeH81SvqIgWOHkzq69iHoqQv5urT1jxuWNEIBr
nxRjee/PXqHgtWZrz2cTUPfzxjNyNF7qVWEXjTF/QSZD8qZDfl7nh0Yb2zX6qKzx
IgcaRjH8CdIoBw5K/4Nmn5uRwLIsaMlLQcJ2E6EB80WdmaBTEYgI/8HdqmZogOof
4TFPpAzw1NLc21HCCZQ4OuGfObNTO74QrjYtc/ffBic/1dAigHVoe3J6NQeP1Mve
RNPxOUgPAGEKESnC5l9tESF3j5DE83OYkJCQM8/phm6FzOlwJiZAu7TK6G5LZuOz
jtxXfbf6razY7ql3uUkbSOId2lxKXPZcOXGv613WvydGWodl8QgtMupkUCPWyILn
S0dSkXNqp5opmJOTsMgAzC1Q+BUfgQh4KH+4Gcd3foO2KMsV6Ei0+oRQ9yDNlnle
7HLd1dcAqfan0te/H9oCywZUhRkHP3oRDsDrWCbS988/8OEfl93I9ehPewnjUqn6
AtYO5vkbOEnnFJF7A4JQNPMJ4e1a1m9DF64E2eprXc6yMwB6gC78jz9T0c4kcUys
pyuALHqYCdrH109cVKblZcul2b8Mja0ovMOpNyDyZaf7fSDuaGuTG4UcoMR32shn
Y4nP1BKxhgQeg/bSjl7qVC43QQ2n+ZgYVwWpZvUcfNmXkIbhmLomCUsvnA3cPS2v
X5H+BLDISQN6CXbsbgVZGwtmkI358ByF8nMfphWZY0PUpHxwKBw/0Evz9tF+uXqu
HZfMEKLHaeE/g4IRojwBLN8k2R9Zkfo3C9Pozk4OWZwgUZkdaJf53SJQbNQAI78T
yIZ69x1wK/uxvzulKmSux9jHFRdUfxUSI0UCrThYRigOa6L4XqmoGmvp9LHVN6nP
GICaY5ypY3mWTix1oxq9tiohxIG95GPwVgvpVHpH9BcLowtgdSp7sThDhwKcdLHs
UseEM2fIhEiHMkuhNVw5X6DDFVbp9JXkh2EwodbVI+lUiQ6eRK8h7tJigHYh22Vc
k5AQFeijz9Qjo2rcBWRVOTjavc573Zkz4RiUxQyF0mbjf5UAmPPa0/3oVFucqYIi
58tWkYvmK4N07MjkVZ9I0bYJBHlYDMW78+JyJAH5BQ7MH9YX471g8PiiiLrHKCwp
hV3mXlb/G3t920oavtyh/Qmvd5FXX2zRIOpzEd/kKyNUkQsynHx2Aml0Kmi/DesX
VInHsftkwogpsEg5HanUttzMIqWYlrO89y2zVM8hf6Rg0Ajaz+64qETMTmuYpRG2
dsCCyjkTcIXSX4IiCXF6qgebPq8Kdo1/NMsvaMuZU2fMCf+aazPWkkc65zzNw7MB
/A+tW7wW5se7GP3Kq5i2I8kLfFmA+GHjr5LgPXZrCHEuX+nZtjdK93skXGSXL1t+
teArR4SUhzahRDIGxoMzsiAGOBWYLFV/xdRigpj5WO/xfpgQ48N9RAItUUowW6eQ
6uo9LGaTmktsTxw9bmkjBbD8p7NyYZP6X8AHPIY2qnlaDwO30W2z5eHfrJ5GL8ni
9RnvM6tVwYiJi+lYmjNDWYoDnAcIUamiQ+HeGmI/5FEr9YH+T2nBAvmG5OtWth+A
rEixfct/e55BEoKVytebGd6Yn0SIZ0isdo1STeLLmZtgHcCyfbDUe+uSlYSx578u
iGIPAreWD3fXPW6sNlvH97ziQoDZdw8qNOA0ny7/XyeHakGgakN9Hshw8Dbx6GZs
b7JZrSfGZioDj8Z1eTSFiU7AJ97VAoh6Fet/SWSXbUOdV+cVJoCy40D8nRHJpYBT
XA6En82UwZ0g9v4TXngtXkd1gKAAeAL5XjsbREVxr31oN+eEb8SJ6HUe017RLMaM
iJ6s0ffexBZbYewqcqWNAbNytlKNhRUI45JnQMn0cAFJnAGT+KGxjUHmCRNU1qx5
gcjRNmokpaoGSHGjuZHS2kbKoxOVZ0PB/DHvfYyWpS9ODKXZPOOjfpM0yyxTDTrp
qVUR189nzXR3tK3SZRtsRexXhCxXPWza7Z8+Fg4gxaP1rn/fJ+QzYaFt2A5TlXpL
iP/JVaWKZ7vGqcg5aiqTDA8izQFGrmeGqUSoIpLPowN2EQXKkurTau2kyJyYO/TC
YpOqfPZeBye8XxSBtPg14mzRmxLc3gx3axlk6iRPvA57e/nvtNPe39PmtHqrU8Sj
GsHe2o74uNU6GCyMz1x2CAHf9GuEpPY1BxYEFc88KfTeyhbtsB7kLlUshXEXfLuZ
w0NJxg9WIQjXdjB/facIaNoyKRSHUjdfWipbNUp7w+dsHz8Kp18iom8wQ3qZO2ka
0kxszr+2Tz8xbIbabHhih9DuQHyfLITgoy4952D3U2mWDyZLLylm0XpgEG0nTtwY
oi7Exf2BCc2EIgU2JmoG4CAAjoz4TgwIDqCtHCE61TqsdtiFuUEukqjN7nOrc0K4
JaXiFlCl/mMZYnaO6POonp4I2vxOjpIlqSOLwRRDRs2ZkiJoqCYp9585P/WJrdOk
kvN8rsQaB1AS9Rsey7ySJ+9QBqQC/cxP8diswJJVvmQNsIEJozgif5G4wMcsj5Jd
VOgkmNnBjQswg6QlpgB10mEWPl/q2lBMm8id2HrXkBeG2U10bxvswzHY83nl3/ap
AnuUF1SvskLcLcQIFiBMzh7LKq6leTfsGQTVt5hHLdFy/X+9kp2xPBdDYBPKkMrs
QCwU9RZykhD/dz4TV/rfDIryAANlziEaY9mtbAGU6VD8le4bnrEhmrDmdzISdtMk
yk3I3f3pTHGY2S5Ox/7Zn8U5kl4L6ZAq4Lmc8RUnVWAoNIjGeI9IA0KMUn9bkWYB
xZAndVMKv/wprPLtDZStVotCEdNQqDnGL84+nMh/YFGQKnGLQ+ZpHEOp30fHOa7F
GBjjUIzSKsiS+I9P2dOL/ccoJ2z9PCXP76Ql2+0QWteovNi48JuhAz/zMuH6ETZ8
HMQU3IPfcaD6qF+8yYOXIcu1xhDbO8JTJwdRFxV+IS+EZ2Mqm6hf9dtrnAdY+fbZ
6L4v2TYTg/7HWRn29/G6Jh5CboyvlCkd39HIrZaFcaASUAkiaDXL72yvuAs8ikFy
oENDJkCxjteAQmN29o3JFYRmmBBCjhb3RjsjqCIW0CX/6LNYhaF5R+IkLIKdsktt
5cMEol0HyIyPmxpz19w9MsYPjR/sCCvsS2wEVwE7KbYshZSv7zecpI/oQG/Sxd4X
a2dYVKV7Vgow5+XvvZE1FKdlJngN4SPa3FBoma7hg1s1ybOcSp+4GWjl2JTEAvxN
WwB6L9FgjWDKiooHASMAE7elgmoCG1sFJ2/3ACy8iCck8LGQUGg3Y6z4uHHQ39KH
F+8FYcXwvufIAHJ6k+ovropPKxtJKBA9VmYJU1eJAPKCBeuwarNHhAX60k6sDOo8
9GJTULiTGw3xPKJkga7qiuONIB/EeTS6eZQm1zNzWzgHaA00tjscCTDRspifL+56
kCacMIezIUcKOcfILzvoEU3yz514BB0xcfTtUVIvezrsTXO2wcMSosETInfbqFQU
iwFrvEAnGMlRcFaaYBuzmeqGueSuOZtFX6NBWQ57eMVyPKFlo+VMqi7dzvD73gjG
IHrpu0PY7R0gScdwrGezE1Gje3ZudfPcbZCfhIiE02ulNOfLButq0bYwdcjfJwi7
VCiTYWUwskYGzLntKeIFEqq3dDSLJqsfJPTS5SixuiKRX07am8cq1vWLwoDYwXBS
I5SKjbJDcjbLv56cAtefSca73LCdharVMhF5eiDejvGEy1hSK+46FKp+zFh/HTRn
Qnlhcj43q/bwadps6/7X7ERo3cAyPZ8MA5E0AIumYVOXnJIBk5bkgEYqYjqMUwKB
Jt2X87rsd4v5htoD8TiWh0pVsSgEAigEQHog3aa0C+pPWC8ZnOs0CpIisE1ncVTh
L1GKY1EEkv0TUy9mv0DgEJ3pHxjbtDOft2PMPjE5Wv1fGEsE4YpCbRpkFjUX+LB7
LutEV5iMG6ZckTYMTfVzhxhwpmHOOb6xnz/IkzbyWUrkETDsBHL6xos+xhOHZSsh
oGKKd2aAD6cXpZQQBYVnNJ7W1S2q4x/6EVOdXdWMcjLgfh/tJ7uemx0rhU1wQ/1w
KxgeVpoqgHu/PcXDkOXMyjnpX9u5UgN2TS1nbSQUkrXSsxyE3dDutHggKu4U24I8
NgmyxT5zXWxRBnn7FM0ariUyV44n3pe+cDSaQymaYr1wOKnrrU2A1sYdx3K4lOP8
ekjDj1IWrAtPjHUHaN/6bj5DPaZW6LFttfrLZO1jzJHEt2AN/dsZIfTeTveBwBcc
P2xAOfpL8/OUJCtokVWZEIaPWs3dJZhAkFhBNcsmjaOroS+KIlDP8hCDje0wxVfI
/c67SKOpDZep5cxM/WcgRQYiWSXCAVBrXEVKszk9LNjb3kGeJOFeESJWG7sIv+Zt
aZEdLnYyJ4FL5zh/HaxlbzJBn4NpkajieDWMLHrPyRs1HKMGYIra8hBWh+vz5QH4
1bqRG7bQR3RuKQT8lfz0xXsaoEeGLEa+Y/Fkw+UOV4DEpBNMscwGWwK0nndVxDLF
cj95X+Scktij5mse+KbxGFgp0wKpBIVHdqZ5NFVWcNXATPJPb7ZB4XjiUlnkbuHF
zYNm38Nr6ibAlNs0TqIra3pqfZ3s/cUWYSqfq5fBbVDKtBqV0uN9jCfeD7ufxEXA
XqdgyO55+g/t2xgwDwC/OwMXWKQiAYBkkRLNXat9ATmOHSNgMQtUQNyLnlQTwhtW
ctXAIsdnT5CoIQ2GXDBC2CW564tzFczlkQ1tZaIJIEt8ffVbnXfuigz7CUYgeyDd
KrIp8uco7Dn67BevRa7vgM+sU7PGhXz+5wjQPkeN+QNPUW/D7S6g0VH/6Neo5fSY
fEalb2fRh3VBg1x7QIFwDsj55HJVL6QCuWIS63ODak628zfDNPgX/ALzutgQiuT9
eP+ws8wPlfRTxXxDLARFAY2SqEgkDzH7hm0As4q4RD3lpc8+Atq2djYdTHsteWwH
kmDRf4VIoChC+Q2bOQRzNcotOwBmr8JT1iu5LdkV5nympqPJovZpOIpGvxfiRoHN
TzYHv911ygpDp8oeWE8xdDSVVdP7BXToXJIaPWhJ9JB4sEIt57T//zKP6ATfgq6J
XVTB26UnUecX/OzG+rTu6J7hY5PfmoRixt8TJnzHceLNzNDltGAJstwjkklIAw2W
vcj0eaiWAxk5TCbSGrgBqKNsLPaqwmCAdxanLuhudSQdAGgliqYfzDtJWRLvZpqT
ZXW3q/qVH7gwGLuYuYAoxSMqqTyrS8MJB+WTuwKqaL6drxSWqQ7FteoLwQsBy4QS
WUGvlb6YR0B5t//Vho0HgTPeMtcXj6HyWD3Brm+3FrKAdOymFE7TxGExjEtenkmq
M8LDC9FF3BFoNrdZ4B1HadVd6FapxiExa75snikApLGClx+EC8YFmG+MMAv3Fpsg
8/D4uovXKfZWdzogNvxX9Bl/X5a1m8NF1bLgc6plR6B5dzoNohwAXkYta9gUh96m
MjMGlX6cjb/L74gmid71Xr9HdAAyiz79TwAtUH0ToNvPd5phY/bRkzDKt7Rmn//v
+5bQOmXeeEIHgRzi3xFCu6QD8rNUdddVHFMP9LvE2lOhOi98JjRYec4/aAXDWMCl
DlXmYkkNci3bYfrMvwPHrTOdtYXmcI2l+jF92JMo/tRLJiz0Nm0tlgS8twnh1XGp
7mhAzzwlQ9U2MIdmVvpbs/lNR2loXPc/NCQO226uX6wCtSnymaXwgfCotn3rumGf
aUnvZ0q1hIrWUan7FVF/C12rNj9n1pn29517fEW8RRXwYuEuPHQnDCgKXUre2Wfy
fU1BQ+OTWvpMSFWMxRBcGn2P+qrK23Clbxzn2bb3x1lpkNfnI5W5xigApmA8D1Ok
UQiEnmkKUMCtMAaqWS+CKsBDVDUAMkj20UiTkl0QS0hxNYRqrCgDm0Xoq2qFhAsg
1A+mgJ9dXofDB4PfsUuTQ0yNOtCBavb0Wtu9mB25Mf8VZUhkmuFHF81lFlsWSPXx
e90pPaTsgmA37rKUxoEmY7h287j0GjVpSa/Kk4r7VTAsSXDLA/FerCnc+cdXCD9D
1caF9nG3EL8YOWaxvk+1a5dS5YU5BSFihGwKHROtHFe4PGwGYQYji9MsVWPR2yXY
YOxHp1DsfSPV5ZYL03IAyPsgHumNf0XT+p8tlYbgnB/KUHlFIlxfYJvwNYm2dp+w
ylGlbZT1aGpqMcn8XBVcIz36NHGh0DYbTtpx2lZ7dXEvQun3AUD9eef2bg3fzDrY
apzEdo9AgZn8K+4ee4hYxjFPLBKwtMQUurahKAErfQ4jeTxIWLR5TXpvhGAd8DO6
F2QnlqcxO3A5ynC3nraBpDC7GmxC7HJMtONGyy5BjAk3/5mq0Ahm0fPtRpn7vML6
eFu6vIuF1471vDxeN/q0mCaJiAgmMDYzfmESQuRPXaZNTWip/MsTyPmDI4q5PnOI
Jws7S9Td3K8am+B9sAIOptDhtRspMpNOy7kLgie18lDqBlx7RSzxoPu2rYW6mnq0
dJc/KUg85IAU4mYwRao4ZF28t+1WG25q5Nuyj5TeZRR8HJZmTAHOfiaqCncmLuUu
waUeg3PzAdno93pnwv4Fa76I8aZtPr/7Ghy2LLonTk6bjEkn+n99u/LFiPaANlm7
aVVNRwTX38TMtREkYKmLtpQ8rvk/7Owc1Pw2pdcZhC0rch3+yki+vpDgGrlvAl0q
ipkMFLY3kDZqjhGFm8+/UrDWDKG9xfuuYHB7tQe8PL4wPdwJO/QsJ1x8JqRsHxXK
E71CjgRg8nZMq2sCx0RB7L+HWK4lGWrT/hDUaUiPc2WlfokWNY6ayV3xjTwsPvE8
l7YMX1HQtUwgkYpaVhJEMAxSZJct49RVzMUyZcVGl0yUny6HxPaxGGAIjqGpSB/m
33r11lJTLkWOU4WYNz6rEOxLh4vSc3Mxpvuocd3hLH5gQ6hGoud4wvAzl6EZo1xv
D9DwAnHOYWrXp32KM9KD277KCWq+svQyaf3zG0gGP3i6NYIhkdPXVya6CEygsRWs
Ou7ppw9L1tU7g3bRRRsBTULp0P0nT6Ckc0qZ3jvHJYbfAcLXSfObF0RydW0ZoHQU
G8n9QR0gBlYnVDnVuJfwStilrd0ytpc6HBDR+l6bVfYLDo7iXF4XtO5rquKSi1ZG
MDAljRc4vyV9QmISoV55cKB/WKeq9DpnvyNvt/VrST1Ra2Twjq0olzGgfCqfBwGi
66CqwqJ+6JNzsTyw4GG4yU0Krgii99QpM0gqzUvSFR+jVq/hr9kOT0dm/k+FcN+n
jATv/L4qhrKC7akU55+zwu/PZoKpq9a4mibJIJeG8/LfTmGidRDtJHsOjOGj9xBi
l62F0WfE8grITpVQG8qFpdmJSL8NPg1hlV0bZ0xMcKinlrEBvHN907nibdSptd+2
ZpcIjeaHi2QlVvFIJlueNIgnJBnlcFtPo5fERYh5PlAtj3PaJe6L9s6Uaj/lIhH5
CGhfoDISTGCRVa3xiM8HRboRCpJ6vOiHzEdVTRbLqlTAZbU9Au7NLWZrrmDzRQw6
jvJw+2BmvS3sJcxp3kA8xl8dHZWvRKmzNabi+C7Brq3ROYjiAV6D08F8CNkDLpgl
Arq+Uxv3JbVLqt9Av5AhfN0hGzQHDyQPT3blat53JjC01W5eavIWlSQymRQWnmBe
toWUYNFVW0jLSlA8u2HCKdEjfsRimcK1ehb+CoLLI+Ze4NL+cZ6mjwu6XfBNRknt
pvZARUDsnzz2fu0NDf3ojqVnp22Dj7zB1TcWgAVR9ctODPeSiC9bjrR32zednSNY
CSrsyAtodz5IPMltzs3JEdVVfVfxaN7nYsBRHj8wAY7KpWHDGIt90XDYjdjSF7Yn
CSiSTHLsAepDv0RhByoR+LTRyDuJ3MPWOGGrt52QtJAgQngNZ4wRCLUk5kqPBNIK
ehnPdu98FShnUO8H5TtF7YqpoV9frduPKw9anZ+UlFzmX+AIu6DMEyr0GnizsYjJ
oTUVSd69T0Sxtpcco9O4DSQAkdK58lyaAab2GX+gT0vBgP960BaLRoCJhg3KGLIO
1vDZMqxS4YgWfOmOHatsyRYUjuUW3V5z5+qpoVO6BILbY5ZzbJYXyclmfGy0TVU+
WtFW9xcRVxwFEZ4/pt82cXt8bUv1QuL9TM1CQVyPxxj4BT1ESrw8tuqvdmFYaswG
wbp1afhDWJNRffQ8dHVCsodlcQWEsz7tUFPhorTHTzy9nRCuGMMoYr8wSqL/7BWG
QusaVw5Qlg2C/esw8C1L4ouT8I8fxI45wli5XYPS8jUG1hd86xB76cdyuA7uiwl6
2WtB0guaM0q2QEORHDa+Ozl4F8pya9E9WFTth2+kW4KMqeyKgEMmIw/vIVsR1QY4
1VwtqaRfnCmJjNBTaqLvK2AuElkKjUd2dH2Uk2aJeqRWVeyrvNfVV0zh1dRjUut5
VeaXXudUjdvT9g5fhMVFpAEW/P1Tj4g9aOZ4XkCR4AlmObl5tm4vOdIHWs8INfJb
YOQzRCNV0Knt5QgsY4QSRObIJXdnMN6+rblrtXaXBIWQpubEv4Knwp6CGX2dtXWf
7+1KZ8vI5/hL0aSFagK1OVaABl42SkPe2BTwxtWadjABnirokRowvRVXtLC2AKkB
mpeH3jWfrSeAobMhM5KL3Qtonqg7w55XiWj65FW9DaazF5iTBUajQRo70ihUm4+a
6dZ9h2yLMjVvdcDGKsWziGO/WI8DXFTtYtEBEfhBrzWLsMIKwslyC9+ZxlaEzXuG
iaO8nq1DdsZZ/OVHK03Ne7jIvfviPap/k0hfBbqaCsl4AtII8rEeJrgx3ao2BFjC
Hs9civ+qrUHXH2GzIHVPGnbpYARgTdKZPFQ/If0IcVIG8Dw/kgAuXf7MDSX0ZYNr
LIbAR0eoUtN6dJa6DecFZVXSnMppvpMgtIPH81caezYMsVNCHj+Saq8ozzc+8cGy
ET+MT9LwZrdlUZXgtbKlSslAY2+PITGgYb1qWlu5v9hq9fnUuKCJ+3Pzonl6D3qk
eKVil68zvoUDKJiCgOVcxn90nZQyaCI/kcS6rKKl5i7KBb8MY9f1qYGbh14uuk5B
rqCLZiv6w11dr4Jogt5A5oIOMmCVmONg7RkcYyE8aHuw2FF1E85S54Y9WLbjF+kt
fk4Ud5K44hFxrh33yj8NZczewtDWmCEgxkUJWbWtT8OGMa6fSHmhu5fJz/xUL2m6
MXGcr0nB5X/RoVT57OFAzCnwPXKdDbQzTHmWAkwnTn8ghol0rCimjm0J6Jm/CTfh
YxvZTi+YKTwYRGm2pP/i836bL0xCXI9AmVCL91tGeMIgVdQZlHQH3T4paliNn06I
IaAfCschDmOY1wUu8o9PVoa6JJWuvxG3LIdXFAZIs4BPKT1UjhWbnXOmWAQwkDqK
7wq8p4ddnbReQqXbQTKYjw0efx1OoOhIgPjYdKsMk7ORZuznqeV0yqHg3FHIrwEM
dhz75PTnmkS4vdldL5r3ZSWY9jEazU/+7WwXjkzmJos8KgdugDzxfCKpgaQ+2dlQ
IwcqkgD25UyFH1PF6hdidtS/MnjVdTZJ6eqbvEKoULlfVD2ByA0U67zWOAt+6wQi
96dN13vUFnacw6k08j62/0AClRTE5tSohJ4RPztt1U08cMVwrXr/thDQAs+HXBDf
Lw2bu8JW9ZpLgMVwbeIH8rd3EHTCccS6uokKdOM7+iJgIrhIi/Qeqj83V19Sqgli
CTnq1txPVplnCwMdWV4R00v9rw4VHH+q51JloGah11+JNvk+vNIJ9YQmiknQnTXA
aptx908MXYd8zNNxA1/DIUtIFilxj/2Y8753FTVhO+djHDSIjPg/mL9eWTxI3/dq
V4y7/TA2s7IFq47SROOotuvxucyq0cf0Dux3JitPLFriqXIEzhp4an1FUhPePvig
GeiICxgDhZ0PdVvteBtSb6emESpz9d7giOJ27CLnEJCmlr1R1V0JfOvIbm0wKzn6
zol1Vz2dMQOQbKkLs4bkADVgBpBP0uKu3kCKeNtXQheqlXueGBKIUmfQMb+/NVGf
oG0upXEi0IuO4O3HMiyAnFnjVwK96dHrQa1UPOcqIlRjuVuVBMiD7P6VdVLB8eH0
WDKLsAA6LqqfrHHVHCq3x86/IzGArIwxtVVXs1X47sMDO9tfSgZ81SsT0zYWB7dd
d+rGFvxGjhhmPABItacjgPkybsv4PIgqh6HD/0rRQ57y5jy2DziRw/auzDC7iF09
gmUUVzhbg9044wDbiQ3T4hOW/qVcUZIbXEAQ0l+h3hKcDcM16o1iRfffEudfl56T
GZUQb/ccTM/P+9vo8AKtd7BaHO9kRvlqXUfmKn87CnrBtgxPcU8aQ2gz48mp8fvE
/wdhk/d4t/CYPXB0ZlGJHk7wCyPPppVmWi2o47j3/xnU7jg063YW7Z62YhamXw2w
Upb2Iz2FDffP1FcCGLkVUnpbqZ8dyLrXSh88wrSmcUHWpO58vCh8XQYw+0npqw12
on4UgVU5ounQKPlpsfLxXt8t74uJDDCEA1odWQCeIJ25+lhEhdbgDYhxooRzGtaJ
YXp8YwbYuaY4E5rONOWm5skEhdFXu78K7jEsWD8oFOZ3XgaRFCA4I5OIBEdnFLR6
DVTCdv8kc65e7Lkq9yhH5Y3QRVNZP9Oi362UAFFPk0Q/Nhu9mVHQcbl+qk5CQBQ+
3o8Pl8HHJeHk13C5+55vhlhSOi7wMtFgKBLFCLT/VRKX6Sdu/JcH2xu254O1PIq2
cTWqGHs7eQ9XqEqNrvac7vUGORdk6mnJZvclZ9yg6kmEeZXSK9u5MgIAlUuFCbcO
A9uQgp81leOIpdLaghX2BnCclS6V6Zz8fPxNjiusw+5qQz2lxSTYb4xP4bBEvVz1
edyGgzim6rxO5lBfY+nQVTPB3IbMXVEAkoCTS6oRTKNL1KEuH1ahdKjj0kLGPM5i
Nr1LT/QgaYqy07iOEeAnnOEKlD/XO2SJJr7aK/1BhQi8dUwBjQ4u7PP4Aafl544U
m75Wmg77qf8FseGlwb+aCxNWryzETUsCKf+iPMCcjoXF1ptPcGXGetx4tZrUGoMP
8olvvo0Rd14m48xcSN7z7BvZpOQSld7di9FuUPKNknMdshEWeDK38/ardz+8u0Bn
c07Qc1K0xtErarF6iaGNVFRYQCmgM8fN//1cNXmEJtfrQ7PbbuperWNR4LqMoCOG
VfvXusF4Lva9Maz/L9Mh+jWpg1vHYeE3IcluksBvWb7xxKjaw9epf9yGaDs9vjf+
XTibtXB50eAGsBQsioFvcv6fJYPGt5rjE3yXbHh7i8KWjwJzIMTWkE/yLqXHY0eb
BgT/ggSDoIVhMVEOLORc88vj3htugbAo7L1Z6KCe9oc4zsRUfj5jaPeuGM01XAWz
j0g6Sy5pVnkPgJx+6tuCeY4FK+RP1XPrIv20KSnAvzbq2OJcLAwQxLagxaxt2Ilx
zoVfSyget0t+DuvZqmNF+It1QrVXMMj3yJZ/ntsdhq3P/cDq6SHQE849dJS3FIT4
QyMqdfhvbun9y6Jgxu1RxmDTSYLdIE+NYkkVesK+EYrlqI/L2HXFty61YcL68cKg
irxNVD3SQ0DbWLAcnVxIu1glQCJrj4rUwHxhswTDoBDnwZIqj5J9FhRJCUHY4id2
CLPhaDWwO8v2SWBgss97msd5CNgzYkPj4j7OpixBzJOTvzz16yy/1a+Il9AoHFil
Nf5M3rGn2wcN8esS4Nd8qOYikQHmfKQ3NCGJA88goeGMdrOKag9QIV1AzoBA2xeP
gSQsoaNWdWFGqzZk356WUg1viysqU59rwg7A0uHMeQ5kYZDPwoO3Sp40KqAzNuuo
xX1BtbLoXuNlfakoz5QEF9+Lfl8zoErdEsVpFFkqkhjym49nhOtywXxpP6x0BaZa
Dl+U9ASX6L5NyTyo2DgPQw4gPBOIO76Phz2xOCqc9r04SgqyUQQvAf2BX8FPTOoD
DClrCYyra80U7/aEIsEHZaNSRu2E323aoQQSb9q9UbOw6Vh1DUYe6VMexpPy4L4D
GthHYalbkOQlIgCZl/spiNA1xyMXmNKIowiDlEtGfz7J93WHjgdjPXlQExrv6xqZ
VfCUQYs8hXhJRyBGJTvJVeob+sLONB/Gkw508ZK3xZ+7XTW7JCWiXgGBZyg1n/wB
ZpG3LFklVk8XIsed1qq/1tisfbeRuvkCi5YhTKD1vYSZV7gUmpTF8c8tpjfK2KYs
HrxQ+uia1A2QDLH6li/tZScY68gymXMPQBj3yn4nEhNBpKMRlIGAWFi1+to5jdls
n4AZcP09n75TULbsT3IYXY0h1fix8SCLdZFFJU5OHrfnqOtuT7Bo5+TIXiSL0AuF
1F3rVTBbER5BNNz6WdOoBPKtrI4XwnhUdwfOD0dG/4fjFZuMIScM+OqTqRsiLWGE
p+s7W4jOFNvcvCEpe+4zaXyzYPoRtRAJHSgbEHRBxw5sxXvzM6sSdKvDVUapjWdy
2zbxckaZZyYyBoyDbt4l0CN3FAuyKxbus0QWFQX0FAu5KqtzTjVFqY3s+caVBGQt
igiKToe/R0RoujrB1/wcCtST6bpSblLluOhRuvqphiGcAikfjTDx+BnuzMYwUEtp
9ynxGKsDuTlnYy+eLyO75RSFhpPXu0m4DjoidFbRsPVqkTlhVTOa1SnRzek8P4nS
xoEfNU5d0fmibCwLOjc/UM3/hRTRh+cU9QnZ6xG98iQHyKUo62235bCWd5ECYnCk
DLx11e+r9kduZOV9R04Z72Uzu/WYgqV+RlfU3dHTsapvLbX0rzXAP3WoQIVI7ajK
lpY33eO/kOxA7JeXIx+inPykWBSLPFQHZd64lJRKvOrEyT6XPVx1rYooyq70bIp+
sLaHIX/lKAQK0EE9bCJxBHH879XOK/k5H/rMwv/Ss7Vnm4O+fC7RZHXTmB669W9J
dxFpLtmqroQ61mBf9fulQVw4CyV7BDmpf08PLxKDtsqorG8N4V77yqT9epJXL8GM
H9H1WZcyX4Kk/UO4gNpjXG51W6IqQqUMyMQipLTmaP+0XeE/0ohFeOwOOTByC9tt
tozQ1GzQs9JQGLDX0MAsiL7tE3zvdvkcO4/Ek3VAd0DpSqlpwf1LOW3d6N+/VWEp
VgmSozpa51ZL8enWdoUlaB4RS0wYOoItHtnB9Hvj+lvyYIWo5Mi1P5Yefci/E/ar
XqLpmBnYBIOT2KCvCEyfEEAjo5eMBjIKk6FS5TjOSH4jo4eEBnPOGpK2Y4Xz3YAh
x5vyPbr+XVsovQvFNKOGj1s11AEapM7QUjowwnH+zsEjQ5SFAhSJVX5z5TlWqJxa
FjEkMiJmwoRG3yiTspG6pEJ6fM0/7mDN/w2yWY+0rsh1MpP7pCNHMb0PsFVLWv5D
LgP2xx/Aid93q1ZstDvWvV36HVfeTOcpVdymDkyijzgduq+TgBso6NWfi9WCfZll
aBik+5tVoeCfeJi9/ztLvM96kcKIuGhx+WGdRn6Lzq+uARjOafFj/I/4hVKhMojB
q++Y6AQbamE8RZ+yDD+z3KqmABClFQQdjYseC6N7yM/07fBTQ8gPAoYK+vJnrzAG
fIRDMJO3MVDYK/ZXQbd4DB0f8kwo+Q9d3gxT3tfdGdvzBFuFT4RFd15jvhKk+A+S
vzvTRleI++7vMtZIiLJW6jQLCUgSAgl8Mxy3maxpYYQG1ABGrwEjWo5W+wrA1GAF
krrVH9k+AAWltmloM5z4lesruzD9NB4TAxDC2lUfLFl1CB1QaG1Fntxo/g4ubDT1
2HyC+6bj8Li4JVyCpyHNnfwqb+E2dc+liqSHPtSylv6hE8QG8CHyf+qmXR9QxGjR
DeFPEqgOd4YFlVj4gK4sZVLY8YyP/ZIAc38JA8TqhXxxtQ5NbjxoSmbzknXgerWo
+G7jYuqKOx0HfwIT4zEwJRYIxHa7MoipRq5euBNcXnWtEjWyhEaQijhH4rpTWX8O
pPpB7THxIXR2QHHws06K3OZORZAuL8o11x3aiB8ysMjOPeUYsXxB9Si/zkMDPlQ8
R/ZAMyl4goVpuFOStb2IYfbBVGQIfofC6UNqb1bgHJUouNMUHDsdGsgOubXeP4fG
XRVNhhK7shhDZ4HPYSc2vZxjeUuTNp8DwK+8KchSLVGiD/Yu0yGOfXOyO1r7ziaJ
AFiKVcZem99isO1KPYiUEyL6J/M7ELyu+OIwolS9GPCXmEvs0lkEHa+uZFBMWqhs
w4QbZM+vVC5n4+BxWLLGEX7dkqgwe3IM1ICQPB9cHm8Uc3VL/5VJIPgcYbZRLuM5
pc68YG+3u9CN6dR8Ebw3XkZhle6uaq9T6SjJihhPDJdwPY1l8NUTFnJ6MZeOiFlG
7Yo48EKhLElputRuOprK9rRsgDSOpiyg5ihnL4WDb14WUnTdTAyIl8D0KSjkDdE7
6LFbuBkAdn6RXvYkFYoFq6ci5lfwRaQFOMUe0iaR5eY+YCb2h2h0UqlV2m+C8Cr7
OuZr4kNdHsTmLc7BPOt1oMFy92MizshmUU9K/uIobf93ot/dlTmfnuqZJ+mRTbCd
Hbwo73kMZV+5h1llW0TEb44dQiqCJLRn5wKw0p4wNlaOaqI2lhDkez80QXsyiWdj
ttcpfmGHi90NpD343LuT41bEaUYt6Sq/AgJxoK5zVKMHoAd8Hb1KsjBWp0MMVP44
Jkl77DZaFmx1cv7xTki3NSU/vr4jImg2LXvP0i4uzTQBieJYMwe4+ZAE0eIWmHux
hsQA8r6iQM5hIjYLljy1K7fJ4tnd6x0+HIsGZEJtcTSa/FXWKHWJmHGcrKrPf8jG
lxkgp5veFbe4o5RzvP2YGfPjZdEWOFOINeuf7b1AaY1e+lrprJ7teYJwAQ05QPTp
exOH/yLo6hEBaQI+TNG9TGzHci/014Psn5HVGG7yntXi1NYAp2G2HkCS2tDkMGqL
oGGWjHxS34Nm47GuxN+xFIY5Pwd/1uXQAre/9ilS03aedn1ep7K9je31kc5G+p0i
2xSIfugb8Gch3T5UkA2dnRhd76jwJufV4Q7z7BaokieyjzFuXGNeInEqt6MMQ7Zc
A5ABoqshnB1c8pp5qxjoHLcAe5vQHZ9TVU8dcaFaGxHNPop7J3txgYPLuW/0B6jo
CL87E6DE9dysp47BjE6ZBiw3Uikkz/WrJYNh9f7bv2U3PZtuqlURjxC174vgcSvP
EZFBrpwJILg4TsBJtTS5WuC1Wf0r0l2iqfmnRbx+b9K44CMsAyfeaAD0Bb2r1Mc1
UtiTVQ+oZ8vYdp6o9vX0mv4EVYY9v5irB5WfOz41TJ6q7aBRcDH+dlsfU/jiU1uj
SMwylVVfeN4veBJffonnODi81jK/47zdwHM2DNWD4Iup+rcSYRisG0poOxYt9vvq
zJtANgyq9aOrMJmr2f8RGQOaSDwOmgwGXTaq0RrdceMnCuWKZ2nBuVTfoxbGV8FN
rhQ+l3ow84jBQt3e0OdPdp6ufkrpggWvd+o4BIyHgODTJrc83K2U34gnfdmmYNXX
4mu+TMmeOMVQlJ4oOx9zIaa0YIcN6mAmnP5uz/YaGHbZX0B6khbpJBYRTE12hbSn
ssgsmc0olohT3An1MxmnAu0zojdaTgbjHNJO6Oy29dqBIPLQwaI4H64JTHJyMsbb
9lSQb5UHRgMKnOyfP1JMUwMixwttrHDESAvu7fDi8TMZ2l7NMI0JRtR8fym0h+7F
XYIVQYLe9+YdK/1yXzkEBBlVUcXhG0plVtlNKbZMt6Wn0TgSL+ZZFsjY/1yZG98b
WhVFStklDFJiZgTF6HyY0Zpg5QfX7iToVj5u4WMPoFzv8vBkjL0u4lSOoWdUwB8t
hG6EPR7lHCXtQnWT/D+Ad8GfixUnSsjKem/lNuv3rpNM2WiwmUJW4ZKFYJ+aGhEn
kjm9og5b5Mz6TbEVucJGVcGtQXTo0kKD7lp2FM6eMGCA5gAZXep8ej7TyMV36hre
y4ALn0zi3PN8hMvdTaWW6pAJo+MlZZou6SSImT8Q8VjiKRL/Xsg6nDF+45NIu5jZ
haYNfqAF8Zc1QcBiB22xnByoqtufBbbYJNSAd+xwP/9lwnrjuuY/dQo5n4bxRwgt
B4If9u2/3UVixKbNM7jh4rwnZ4D8DWHdSnuzBlrlQRWYj7qVigDttFYIt2eFUgoH
cl+CcJcEtP9j5kOO8/yXYPWq5HBgu8RBiX2u4mlsxNoKLHxg+LmsORDegH/xWGgm
DIImlXgdfea6Qs/+Q7jNB+0wcxnwBl0ZzY9laVpHzYQBH6dZar7TiWEwPv3vZTrn
Ms8lOJC/qOJFAfpYwvtIZcXzTlhZg8udegh38prFx6UU529uMJ1ypVQp4ET4bqGL
Qx/wgBlWLuOUXEWQTYEr46ieO+VUfBHBDJ+VousLCBZca1MuJuEpd2JfEtY4diLB
f/WkRPh95+Zp2DqhopLwXLo26TdjO6yEny7VZEmkNwzQpMnODhTilClH/hiOrd5Y
T87RWfbQ+R2aWXAc/gA7pYjbBKEyA5Fn8hc/+PBjMXbvAPhxiAjpXMJXKihxl9cO
HwdaCJenrAkP/7aGYHg8KzL/B3hNowqpa4/XALsgROxBHHYwpSPN0YxcAdMJp1hm
1ykPXDRdtD1Dgh9A+EUs4QU93ipKjZt3b5r4tR5BugqUlnwjCk5dHXrut6Si4O+d
xUbyIjn8Gt5+hnh+wAPnYzz+7f1LgvTERVL1YnTPLvhMYjt+NhNHL9cus+NuIP0n
1cX5lnWrXnBmPwQyv63+0eZxrdkx3FRaM/ZUKjjyfIlDFFrBuCY0uuCEoOQg/f3i
8/zDdvPtnPJ7PIoPtOUq8XD+z3yLXaTy+2X4mQzC/QzhyzoLm3+hbutcoCm5zMQH
ti4sIiQR8Qql3Q/b1l+k/wrn/H91Q+B7lD8MRdDyVdqF46n8hxAnxtFHl9oEPa9G
MbXqQHkVR7CNkihc42TBtzioOgfWTx4GSm/nhsQhqiA1E0OoRxaflf+iwjz5MW2d
oHbsH5Jf/5JHnBnu5mc/6l+HirKHW14G9lPEi5UckBvcBSWy9cRJj6uxTT90KdTh
8tZwPc0IddReE8oxG2B8P6X2Sl2muc2b06pEgT42eJ3oFBr4BAri3zjg++UumF0O
YbRa2TPVeIWrSQOusUH5FPyK2PfiiPsSSsEyKYuzUMTRkjLuf9BfsapRDHX1rwNs
tb4ivshOUXCNVVCXuBPmP1jXcJHafDgXk92GLE89w+9X2H6sp+HapqDo4CUDVibe
kK+EyxQ8Fr8Nqdt0L6XxfbqEqL1lIJIZo1F6HJ7Z5h0oIvlAXCDNKgFapwG750JN
iLGvp92phjfegiss7nC3+kZy2nLQfHl9H4E/tsWpecJQSPw/yJQ7VidycMOr74X0
xW9VR2s04Ss466yxrKUYexaG3u7QAEXpkO9H4CSIlFhgVDrLp3YgnhuFY1aGDQza
/Pm8oZ6uvgUjVCiAE3/Yx3B224AM2ENakENXvDgJ7keqRZ0vo4UOG7qgybiTuK0I
AZbIBLCKneM14P5px70Nptmkxc4Tim08SHsdIaG3PXVNinD3TqYOspVwWa3qyAC8
cl4BYaErmp6L5zyAHMMfmYsrrqnP18xG1pegG1du2J1kq99Ey39RwkZUWUUWgKiB
n+Fa9Fcrxg+GB3K537hZ/EI+N34Tg9SnUfaGKe/E9FuBAmqI0sfeIxfDLbgRoA3b
pK6WD0HCSXizd2TmTwgKlOl7xruEjjkPq+xr/RI0bzGBDsGgJN61x5Avlnb5yzh6
FDU6pqlH8ubeZrfvAJ4murs+bOjysYxid4rG8+xwsxR1/xHu2WP9IEcexD5g8qvV
qPZO3VdG/s61VeZYSM4ahLHRoT2VKABxwxZsGqubczCb3ilOjRvR8sukV721NX4k
EZzXd0mOI0s54DxKzhp0aWDUB7qkxNyTvHDv8UC/fFg2DK01Tvj6j5wDnd2ojwcR
otIm7L2x1DU8i9iMJ7+JfMimXsYwDgu4cG+ksQrr6mn7H2FjPpl5aFS3T+Dn3943
K4qYmr/+ciYrZbhwXdE5D2pLfFhB3B6z0GOCOO2sZgmlJ1c/SqNzCZU/BVF0gWdi
aSlVMm/sHSGzswT8uRguI55teY7LfjhaZalA/tQywGZahzjtkBnwjOvWTEbc0gYV
FuhE47t6vo6melQ/9LE/ZBK+mu01lVxTh6xVb8rRRwwVyLHKtx6+8u4VDiAs0LVt
e5tuIPHAKq+RYYBR7lkrMUplUksUzCS5LsXCn4ztNS57Px9UgxpMNtuWCMdocgUn
1BF/cGMEpI/uDJ7vpX0kZ6XaEckFvbQzxWGcVu4f4jZNApHdBWOt8aMrz1fu0wTg
xrmnZ9Ev/xjUj9EiPjboWT0yaxATpaSs0X3lRGCTpORSjdQA4C1iOrirdptsKj61
X+xeocQ/ghNFjGIVHOZhreAUD5pl+vEy23f5ItjBoaWimzUBanJxtUh4uejWjTG5
V5FKS23GyqPGwdhM6lthjfS3aBU2xzjSLGEyTux8TYRwKZ3V+tum3yHie3+XpsIr
6YLgRVlcx0B5o8+FOve90faTEF0cCuxmwwao+NmovyrPHOtoUItQDf+IxgEf7EJ3
+Sd32AKaKeucWe4cFOuOBCYuA6xBnOELPQfEWXS+6Y4cfUkOAqaUrcwXNYDNxadQ
fdiYfqM47J1kZdF+4YQ7B2JmGPmNidJL1bbxZY8qTI+VKczxlsX7aHZ9O9lCPaFa
rP8rIyORrN6jBWbnuzhOmWz6tywOrq4Ths1OpVc04/afddmrLLoAU+3dsCmxcVa3
snczTnttgqLKl9Wfz0Rs352Wf5kmF0iq9sDwSi00+v6DhsynVCzTzZN4OiTvMky8
OfnZxfngq1RTk/0hGF8+WOHejhcPnXkeBZgTk/Jb1TM9uHSvBtlxX3zsLxawfvE2
9n02+ERndW0B2+5nJj0dXoEnJ2TpebF6zwacV+7zBuZV/lzDRaQS2xapLn/dTUb5
xDNOujU4L2hi28H9aUn2Q2xyYYPSbZa5D8NI6eA4uA2BCKdFPCb8puyeTkieEkrK
7fy/slWgQAU/YHTvcQ0Dj+qTOdSp+O+IK1MtyXdDzuGM9LzUkoybbrhK+PpIhwQ9
xgAGoLqSuNZxkFN+ZNXk+6H6VdqFdV45VQXycp4s5Ie6er8kL1q8oSn27hFotQ7Q
VBymNwtwO0D+5sDEFoukuvRc4qDtVKGtInhw2JdFfM5cySnu3zp18kuCD1iXfaNN
yYDoFSlaug9DGfAaokbZb1UtOpYmGfT8L3QfJvk+MSyXDrfrgGpdDZXoYklACMXA
ev8XMBuWaa7dsrovEhNoFay58/quoskEetNLE38C1u/ErnqgfCQqTJwFE8e6inIc
eliuRPEeqQdCN9j7Flj6ndX/4xxtZvHjg8yP2ru34wugxlu1spqJz4zOOx/LxL65
DGfa3u2FDaPdr0SczgB8pC3Kdonszzjabaf/Xq0n+0KQ4P65NnyzDym398skcbCj
t3u2gMuT9FKecLS4C/HNJv0Wmki0hx4UnFA8sDBQ24U=
`pragma protect end_protected
