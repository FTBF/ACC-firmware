// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 03:56:40 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bQfwcQExBFQSHe+bDjI1Nau2N/m+CdnYBVJogoh1/Ij+y/m1k8aCUtEyUT1lMAlQ
8NfgaKxf0YmH5Js20pfaAJNNID+H2mt7xE2uwzE4tWbepRiTdfxxnyLg6Lzq9iB5
2DPjij07azdxCZb4F5OcM3u646iaysXBGuiX4Gutzec=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 57744)
nQiZAoKNJ8ddfluqxOlhFIyNVEeINUy+6EaJ6HYm7gdGTnc+iwjub3smnOToImwc
2M+OrcZmCYHRA+Gm1s3rsgxjE+obMRtAUX8BiRY0bgYzLbOmZwQwPCo/iuPKzBG2
W7uDzchp1JaeVwsIf29x41RDUoag7kZWEBMVGIxt9a62855j70W5dMSW0Oz0leV4
IFs3nWrDIIgmAzm0+spvawWaScK/8NfOj2JcRBAcgqCiIzSKH6gWDbEcmrHLk9uW
WjttYuGevjA4X37pNIgpuEUYD9JWsdrSi5y+4QZwrENA1qxXXpl8V4yFe7TrCdZs
LwLUyFCLsXgdW2bN2Jk9HmKv+i59etY1oUIoslAmVRkUdlPhdJ0B2KjhnN3axdfO
orzgA9EHQZeE15b4WyIKHv5dbe02lUQnOUGVJ7U6MX+p0Z56eJs4FBZnHAoMBFQq
+1bkn/C17AuHIKaP89fy+vC9juykNO5za6DwsMi4e9P0HBOdpYB9h2z9Q5y3e3fg
q90AKb9WJEgmhbdeAFkS+KEw+hhaENqQSPzxteNZvdnXggo9xvp5Vi4AI5Y9yYeO
s9QJX69ig10mI6WfJLeFz3SlPZcvYGVKBtc0vm6ALyJsOUK+ULgM6vqg3C9/TCFs
bAZZJVwrGE7HYNV0S38TziqS08ctTteuIiGioopDTSs699zCMyw+74m2da9xvGrf
wUncJW36ttGVVcgUrga6MbrsICIx1xXk/9+Nh/zyb1EX4z/aQmjq0EEXCNvT2Liy
HEIcUh3tRQ3F6qmxiRSEJcnK6UPZN9dW3FBgQnW5e/QseBOlQkpDYhUkUK49n5pm
usHgpLbPjtF/lzGmeHfp3mUkziEhdDZ1xwxBeP70MP1eMoZOFILx1PfEjQxS7IxF
WEGeYEjWVNqHUQhTdWuL3SdZwkOz1R2WUeiaqy4g/BGUlP/c+aVxwOJW3dKmoWdO
UN2jx8cn3a29NYrUjIjnW6cNPQglvSdE/HhbaON0lJ68JzGNND0iqh1eB2D5TXpC
s2jlQ6HgxpXYrGUrn8McqNNrWEkXsTKHWtM/ES/3BzOds9oQlYksG37QNUTY4sr/
QP99VG3Xq4UvYHXSJCR1Lw3sHq20uKwASS0Pygg3LltbehyGGKfJ/K6vsmeUyimX
M+svP96v8D2dpYfOtJpV+0O5K7y/VpZIfRQVpQLVp9UQ0OlMpgkzK96x2UDXNxLn
jQXVWwFpQwHmpipm+fGnBcDwHhe1pFzXVE4fjbWgFBo1XFex0do7I5/OJBuTHAAQ
sYcTAD+UX22vStmKFCKHQueiS3yAjdPhuZXhxJlJ8s3MC0WTYqnaQMfGoBQK7I40
JELyXxG+64v0//1dGkVCozLSCYuY6d+i+s7SnWU//OecDh+XDzQHPkQ45N/fGQJ4
MRbJomt+/3GNFbAT4MgG90Z2fncGmp92dvsk/Olgz2QrojIZGgJhcCxEL9P5/a3C
hUllR9qFd4Ypr/BFz+WoSSIlv0il7s0NSjVtYkT7A4C5e7ItvA7rggZlEYaJ5Qa4
jSy5ZrG2t+jwGeqGO716rG9DgcZu+IfPShrYR4Pf0YCVp05J+mb5/3tXtG3jydUT
0YqXQ4vzmsLuo27PF25TIGSATwEil9eyVn8FDR+a4Ni/Kr9JA1Mh43sYQFiN58l2
NiBejM7o0AJdlCz9H+HBN/ER810yjA376CZImZzfPIcBHPiLiS1zOZurudZykK/Q
TM9eXgN+8sQkgjWao7MsXvFcmihDmo0YYpdI2RTVAgxyARriAVT+uI/be22+FKiw
UZT2+JVT0KNBVpKsHiyBdJ7Lgdzxu1sDbQO1zDD0S7VQZbSTuTMZXoVETqNdA5oK
juTv3Oj9e1xklzJp97TTOkCNIdyp2t/vZllcVjYXTaIJs+BnMt7b9II3Q7KvmO9Z
JUdmphZFaWgsI2l57O90Dgmq9vTQipdWH1Y9HPL368bAcRy0VQmplRK+6MRYSG4q
6cOsc6cV3Dl9YYX/x5ZRglctDiwJLWBL5p0SJL3wp5rfIR0DuWWYEz9qf5v7RabI
dLfL07OBvpTBB3tj+AqFXtEWpuAutThkGFpucLbNgJeLtuI2DWCemzobyTUJ2Uq9
rzGn1fZklQJ4RyFG2o4s/SLToXOAYJ3YQaNzRU+wrNMZCdF29ZZUZuwpc+0J0TJH
yCsm9Z83zoWJ7CfciVpGsNjhnpkDeYHAcI/SNvR9omnszNQr73D+7HytRzpQks3P
0y0wh6m2qA6B44If/I1jdNlYpsPC0Shz4ywozKmAMbq24g1RGpbbt0oEDs/MacGk
iZ+n9SWY3khDPNNrQ2DW3fwEwxYXNp9wASry+qHcrFl88PXLZSDx9xi/FuGKG2f9
DYQVeSf8cRkafrr+Gp+jSJGwgm01o+LiPtGpVBClL4PAstmVYbfDeTtQKFG+CO0n
IHsbuvkUPo1XrQh01ewhcSJ24Bih1hiiZ5c3lK4x7RyT+UflSe3GkbWYOWpdlhjK
XR2ZNF7KEUF8+mhxv8xofAC5YfxYMrox+ZWROMiMyNQi5YFVnlnrAW83JTYFLfux
ND4gyiRDsZwgIbDCE2xh5k5SGhAoVUMWEhE5p911Yh7eQW0yYJxlXZCmfgw3KFim
Gm8nCA2F/pkUQDyubh99a0f2nFekSoLnPv83bE0zeHKuOV/8NtrP46RdPWgjayd4
/gWeBE/u4b8emvcrNUJZDiUw6vL7xuIMlbEUNuvT9lpDpLlIt/lxMpN8tJYH6aCv
7trLnKxliBEfz5sos1/eze07JXFLrTn2wc/jXJTH2cU9kODy2a4U5MH8GxbjD+Cy
sJWiXxjzOO44/XoyKlWCQ7N9+jqwyAxQbHFR7HgL7qQMD0zF9+NK5o/9y4DYS9Dw
Yt0ARbDTHYrkvxsFHbZ4DMpqj2/T3Rvc8obGWiBoPWXFMwNCI3tYN1NSMz11XDzH
axnzyQ3iL/tfzPs/F0497kHMZp+BooloDdalID6n2UKEQAX8pb0WBCqd2Y0NPyTB
hvw7PSmOOSSVuXf4ObTUEo/KT/vAVGSOgeOyteS1PWoA6bMPwz/qNPz8lgA4gYf9
8O3wqqrTA5uGwjOHvFehI7gzE7ZIs8PpEh0F5Pek1loWe2JYF21EkcqgQnj7jk40
SgrTnleGu+qMkuBYWMAMrHB/QCO4eZoGioz/auKiHne1cgkU75T9eBDKQXSCZicg
l1VB0dy/3B0ESCCS8p2VGSegyzaAaYAaE2OSKVtAlZHeGu6DQMUdYV8f/t+snHYt
CJ4MFi46frhxp8Fn8D+vMIgVfyqpj2H25Yakk6jpN4YOoa+0XBVyX4Bc62OOxeuo
+6gw5rx5/qW22uhxW3B06w7BmovRIE9hEwtrRo/qgQjpVMwjnxGkAgt7eLQQQS1/
N2ZystKdgxdrY++psBstKJ1PPKcV3sUcsOJdTe7eXyrO02h1ivM6m5+fEzL7ZyIX
Ceo2kQQKbD0fs2SXDpvJkm00IlB1DkA+gAOPzRMCEbwVSIk3cFCQ8IZSAIadR/rZ
0lW3DrSwUpZaNmariTG+ghxVpIbjV00M6+PKqKRVILBYAGAsyu9DkB0J6E2Iu4L4
S5vfojAmH/E/ou2g2PFYRGBaocT8gXMnRUgjzEKfNAs8EMEwZPblKELq/8GGyBKC
TcNv9FJ8smkDZbomcvY3gGzv7HRsai8Hc/vlj3gsmw2uLCwdpieyHPi2PPOg4WlU
rR8+mw90rQoz8b5kP2xNN2DjRqb+W8+Oz1dENc2K+mTnxpZ4Qr7WwK8JdZQxJ2TQ
3U4n2WlVPlGQk4lfh/Dw5VtKFem+my+XaHJsTEvGxPTh81CxmXYS3UstaPcI1wsV
7YmM/eKRIsjAyf4/Zwbwr71vwT0jUqjtrkY+ZOVmdl1xyzEOkOGPdKCR1KW6PUX2
sc08kZcnuFlsSIjt/MF5l/buQRVgiKWs27uUk3WhDAT1VBWGhSs8VeY4kjzKoTbM
Muxttv6xRzp1f+ybDUcxTDtQW+4N5aU3CLbF7Ab0rDZSF8msAwqUbPbpgYj4Rk8y
T9QJ9BbL7KMl1tXOuZGBonUYpziynuHwpRi+zz29ge17i3f6Qa9Xj2SbqzhqYg7l
zHGXUg74oRMiRpD0T+w4YzIxCY87OjvI+ta8iOBjNnk2ZvT2sGJUqq6HvWC3NA9Q
SE3HaMEWsLfOCFZdHr4C2r9O0nrOXcLt9NFuI+CZmO+Pnql1MFUtVm6MHiBcgREv
oCqszPsFuxIZgNt67czbLcSI0AHlO7LIO4z5R1/K4XuMOj/6PKQOxL1MWOTELObG
UrgACPuTtxkUw9c4YE+S5JzTh2aDydOsAKs1PpOL4XYmUPJo3eMltBUFnRV4kaZM
J9H5MtUfU4MQgrcnSAoRJk5nncB9y/6yOvYabt+qDbwvE183+QLqrgE4j6MNP27y
TGPN+341waaNS3UJ1+XAKQDifOPnV28e5cIyj+/XsnFpgxsxP/OUkYnp5zMqjOiN
Tl8IgZC5yxFI/+DKPFHrUFhvnQesUO1kXNy3lpWlMDesyI9rZ/AZM1uVDfTSXcbT
z3Mqd6iZAe4KHRp0/gDB/zD92G+L2tppy32RNaf7CJxwUSqPnjX3hlJ3KLpeNXCo
lBzvuniqo6sYmgo3IGo7r7RS/BDixX6XBVOwPC4ucKveDpr36f93VsvhHMxjVCjM
VYcHLvVEteBSlKCh5zMZ1J/Sp2tgYbA1L7lzdg7N/MPhxrFYdA1tD7W5sz+Jpi6E
ZT/aCesUiGjoBxnrOQzPqJWh3zmQ2+WLvWaQt6bE4uS6nll2VPnHhAHtMtwiwkig
Lz1Pf3rUWt/v6fANgnPU0tTbcG/8W25/bbaD6ridJrKcvg4LLo8OW7spJLn1fxdr
T7zdJ6W43UQMFH/e91HgCCMSlGd06HPTrOD0nCfimJm6EK4UsdMvEy5d6d2Sroql
HD7W8LlHLy/5CCXxgDaznPc4HKhbi5sFWj8ZgEjwCJIfeNTlFQKKhLNukNGopY9Y
qlhj+9sE+aAeBcfwukhr+svPXrZaRpJaESqIAO5TV1iOZ9xYGc1NYGEf/vJwri7C
Q7g4TN8G+35FvfQKSk/m5WBAKEnKGvCJlM4oTD5Y7J3pgvmvtZc3jZkt0FQzEMdq
axWEYc+WZM6YzDdahW12dchm0/wW7VIL25D6UBGn26UZLBTq4XAWuQhUEUk7gRO4
KEKxUGDSXZiTw4JbM7RTq+i+cwQD2P2SK8xPYEV1u1ZMiMrokG6yOgUWpIMFzKJS
FQWcRFVGbITfEEJp1546L4oTk7QLauKm+YUUSOdgvFn5b75czE5hPG2KBsCTGaCN
KEPNVRac9KKxteqQqBt7molO+v1VmTQX7miOnzMIunK3y17xPSM5Wrz5p+0FGrfP
YSGrezSZuqN3gLs6UzrwRP9W2Q3qHU/MQHfCHoYhamWCp6q6FX6acizPU6HDklCg
YMORIVtWCniI4a2OJSMrG8q1S3z12Mt1L/rf4Hep2K8UHsYOZKVsMxqIpCUmAd5N
Z1fVcKs+GaUgXseHv61APnkPdZAcZfij4rNIho9V5kFF6D0Xr7XtJYGcMRMqjIan
VfCrStHN8weqnnM4VN+gf7oTO+86UlkYlJk3t6/oSCnH4fNunH2SPg24zHm+9mTG
mlp7pIeoitDPIvSa4aT1EuS4wpYKzJQ2vt2uRch3y5hWLWhHpwPWMzSgFLVhu7wX
Hw/VkiyjqUnFotN2EOmRNC9ylwii1TShMholAGPSoFa7uaMUrFu3WjCbjah+Vz3v
3dHGI8bIivFeCgFUNQ+uxoHqujne6t2HZZyzAEQKV77RR1DmsEz44tSlxmlauB07
0AEuXEEQyFB4V4kDpDWLfAifJ6UNytsPjVufMovRjZYWM+xA9mjw/iQaMXiJZicb
ba0tYNEdWq7FYpIj5SGkrWlCWVDOO9eTGI9goIoDWJv6jH27HGGpCKFNisb1HoK9
ekc8s5K1SyuJc6q6KgoqvVCAk916ZKtOzEBIr5c0RgF57tGApKQnw6vR4s5Pg5W7
Jl7mAZsSyj4SwdvM6Nz4J4PtaFdKk/HD0qkgAo8YjSxIGIL9rNitIxQOQSWcAdys
QlITYdLpUq+k4dSdmu8KJM1WSltJttO885gnA+/PZZW+ANhIS/GHRvmDYjRo100j
plaAbqd0wJIXu7allPzK0N9doM7BMtn5Rq0ITs2Kn69MknTVwDN4hvH8tEq3VwzG
dDe0blHzCcQaAHu+RkssUy9JeR+A4UW2uwsf93TLi5vwyvM+x+Q1MBQ9hMiT1AuX
2Nn+nBcRdt2Oz/GjnEPLjHLQ+Q8N7NK2H/Oyzv9mik28BjtEWT7ZznISynEXN6A5
Sy/HsyT4nRFfks+7A2rqSgIRXFgc8yvG+282XG5ThnSBBHRF3lvKrS82C8qrjY9w
omOlU8t7a12FdMj0XIii1pv03jRrR7KBaYcDcayMZXXjrLzO6sol6QpDps/mBcYX
A8vBzsKsieqCcqUBSBq3amyYoKQP3QrhuHptkWUgHrmZQ3TxSGCVi6Yyo8xjpw5K
pHViuFFr+PX1KLUDrvlq7KbfvV4k6Yxh2GdIZ812dM4LQcr/WREOtbuVYLeeq5nI
O8c85ggjeuTEJeoRMh4pxiKYOfN11hQ+lndOJ2S2TFd8kLFiPjcVD+d93g3JQsz1
NVEBKs+gklRoFojBIqDOEIZYYCdyVrBR+bMxt9cUvwRiohORHTJ9d3IrBQqvFTPu
Ha8uQcWIQdLb8LFK30dSDUPjF4myYH7JEiBlg1RtGV/c3wmJd5BCu5f9M5AMgjlR
D5eS/VBrY++6B2Dknd0SaBLd+5Gi18uLQzKuuCilp4vUQJe934k1VNaoT5vd2sB5
z/XLnTAZFu/2J3edZqxtniVtE441OtSe+1MY4/D+rZZrAUwtAQExPhoX4TIhwzSA
DDoap9O3W9DVMJNX9JLm1ZNU84aplLIp8h451/sTofrxVU33mKQVD4IczzI7BtWv
P5aSpu/ddc5qa4t3YymGrNmSFdZjjFOIZVQOvEnvS9HYSC8XJr+D9KOAYQkD1c61
+w0VtJwS+P2ovn7ovINrnhwW694IOvmEi2vH5oK7zjNWY6TcT9hb5slE/oicbsTZ
KxJcS1RlnbS5J71U9cU/hh8bjzEKFG+X4Cs/M1bkleKzksFUMK81lzvNsOL+g26w
o+OAxBrm9zCE1V+rgg4IkGP60qs/nX9g3d19Y0CVFu/gUbBo+ec7wIFRmgW0DSC3
/YXDet4Iy5o8A8hBBOELSqfoYKFCpbUShavBwNVIALLqosTK8wB1TeZt8FUX9Q8B
eyTj0D4CMK6nwuJhbEidxnN9uj4sIXFdtTCvEzz9znqGyK3nZ+W755ql7HzSj5YP
NKFwwQANES8QM5Or/ZpViTbVmydzbftejMbwFz183ebI9PUsDlJdV9gjX9ZE+z1u
xUQYGV0tSZHoccAoxRdojsc2KjvMeVlkoIjqqjDyH2vUXaJGnpYwSJLTMtNGoO/U
LSVHVgCQJPCHHtAqW2fopG71JyqewwfNQPYpi5YffNwQZnTPhQiLjDFSGwC6Kunx
bVsQjDST2cweT0USWTDj37Hr2jeDImH30//RCTzeBsqtZ8VM2YGRnXTyyfQXwpz8
jjLveA5f2ZMCftChS5ZnLoX2j859ng5A3pEAqhHDoP4TG19m9PJRqg5xsJKZAtUp
13UJ5vjCmNQP935CwcDui9bbSAMRKGvyZZK0foL5zi2RV8JnY363PSdrKgt9c2bp
YLFJ6f8T5lACEnfOnSX+yWmc+5Q7XlRoSNfg0Sut3ht1Sn+R+nPeR17uKU/BOrFX
P08PHp3Q8GKjB4N8bs6Wg+2++uueCUf7pgM2ajgxIfCk67ntt1Xb8O1Ij0y3eVEe
Ztuu/68aLO8I2sCfFqZbi74VMq0K1KIGYJebi+lgX6Bz6MJtlG5TdwqRtOJn+PBR
MDtlyR3C5P5FHKN9LjIcmFTP1Gmpso5TesStaUNo+15aXidTnvpncc0f4dWUSR4L
d6/lYuftX1uQR7DFrux/tvAt31x708Jd+BG573nMmo1Qi1vDkfcidXPPXOQ7DbKo
MjPb5x73JZvgJ48Pg4bnQSMG0hxjpbkjaeB2aHBdMvf1jU59z78HmJvISjaWPByo
nI5KxypnKA6ycqUgAZVq+btjrdXNaGkQEdEjmySs0xLspy8EYILdkWn4Z/HQHRYQ
pUNB66oqSHbcRjJrZK0GJaFmmkG2AyotpS45mogm16tSqLjQYivP+2ej+Flr+TMX
7gtNAJ3fGyX2j8DTraDFUVMhDmV1WPGZSB6czm99yFamBWJQoDnY7iw8bLkMDJGg
JqnIBnUBy0lP8Sq34BPwjo0N0yDadk6k6WbtyGexgW8/danHvJ63f+elF4k4hN4D
Ino+Kw0z4kRyuFqgtCULbxhD5Qn0VyGceqcYEzuaj2hKFlE6RwssL/IG+zUWBWCX
zQUZJtHDXlHpvcT6CXVpMLqAPEKTkk8A8taxGPGfheJkIE/9MTenKY6f3jdZkriG
i3CUQ+FhSEQhk2yELVMpvCmPzyc91djixGtSqgdcb/shcIt4zG1wnqFs7sqAn4mq
g3P2nX1cpBOuYYtIHmjVXoRhmAMIdslxTlD2D0BKxxHPKJwmWqDn03nuf8zfqxwK
snAZolsF7fuE9CSfsGdPHKi3HmSIzXOsFHhDt9PtWBV5mnioJ70qPjh8rSIL1Emn
XGOP047tojCCdDrprWNTSVTbFHs27a2YEUzbIYVnp9jAlC0x9hpmesWNBQj6Uamw
zCa0TKwlRDnG4e7vSj+PYOt+hw4cT4Tumru2DUa2aH3Q8TlUyXdPT8J+Tc9TecuF
PRVUtIRMB4zcU8M8Kw4dmQzMez/i11pTA+CvJY4+kri/osqnv59FQosYDHapYGyP
gKT565dnvkPN/nUdNoM3tiK4f/pMQkzzmeKs87LJdsOtNvD/vAPk+mUwtlnMlOJ6
svT1Gsx4mMPkI1IEfMfUqv5fmXkzAnRLDvmpmZN44jo5srGpoXKsx6u4TU9dSMFD
Gaj+zP8hZkMYyi6fkbMJhB+K8m6ZvTRPH1NZGyUU5otldJOeRP1OSyk+pKb0IhdO
OOaIeNT8GWE45KiZ1wDShYGUXsS3LylLSAxYC7/rL4CCn7Vedg3CHwitMT16QWGs
OA+aQiK0dK6YeCg0v9MEgv/eRgNBgiYf+L2ENkoGOhwN1tRzRaptiQElh/QNPJBL
BFXicCpXoLVcui1uWbeEE9UYnU2tpKkcb7qyVwhmYnRGrIs2c1gmgJclMeBXVbfd
CrqeRxJQn5fwDsWdKZZvx2IHUvYaaUzluLE4lK8Lr7vmLU3Mvg3GuXrZlxPM2Xfa
9lLZDf2w/tzXbt88xVmQv3nojQyuUm5Sr+/z2dwJIieUTRyLRFETwtAAhpAUBvDL
k+kWzgfF3ccbUU5gyFYIlwYNPus7ImyvPJngAmSHqlOyRboYW3Ver4oOpzAJ30XA
hC59yJIXbGLBI2IqJ2rBWYsv2kXhWOp5ZFMa09RgLFDqrv36pfz9VBYkPaqH0cUy
QLcS3FS6fmClUsnRO9oBOeOaGGTSrEa+6agUIowpMF/Yr5vYp3f/9LC0Fahlwpny
5bj4o67YhNXhjROOzKrVUgpy9kW6JEhXDZtWLYwfhu1eoi1OYQ5uota6O6wu4v/3
4nc38liz8EjqKXLIMYHuLtzkdg6LYJNoM6hU9nxPrnnxR6yZScZHnhdPp8GIb32A
yaMylGiGa9nW4iFm8MmL0k4YeVAlwFIiKAGLBaUBxi4STK+EIMHKo545EfKO0lN4
4e21oCYO/7NV+pSk0fycEV8oFXQK7EKz90NdaElBkCQo7RDMCe3mHwzkFiz0GxsN
gS+EG2n36tuyfpkJz2HGaw9guxZIEIXBpjAE+KYQ+Ec9tBbsh95dDBX4fLiMzZoQ
b/h8fBDCXajqGKls/k6Lr9e1TvFRT5ZXe/jX4ugQt6WLdmPRWwk9KyZh6W41KM9s
11SxrQBODaoWqisBhMn/FrHQV82id44LlEYfDEOK/yusdeEsVeAWqL7sVvYX5rNM
d44e0+tvWTIzTopXkzTQJ5kWtXoCxmHw2E3eFkTUhAuVKHzaj1GRGR+YHOmQtBz3
R5goJKlnxmlz1EnMe6+KOBx3GtAVVkKwPFp0vcZIPe0lZonxe15uSmqcT1Pt5G3P
WJCchUYO8iRVqz7icCDNnvk45kyvRZW3ocKd3+vzm52V1jvtTJK30vNp24K1BIDn
mv86i8jGwGzl/WlhUhUMqruA/njROV89hZRaoIMzozMuyENBj5kee2juOHzwf7dQ
3I9hxXbPPN5dxcc2ZoOC5bncn8v+5LC8xLjRPSiSk8a4d5P1/AzeX0K1Ow3yBhQ5
Jtcmt07TG+w5TZscXf388sPT9Wu/MExmPNloqYLoVw64o5GZL6uwSmFip+k8WNLC
tLwyXO7/m7dd6zdSv4TSGY0sG9LtzvUhlGFTdovDtSelJf3l+FsRSnwHWX0BgD4S
UFKFHi07oyIVwotCW4Nfot0zotMeBqdTvOq4Vav40baPspByLtsttmQfw8JYkgoP
pU404bSXpc0Zj1PcUV7RfFivFI97rVhMMpMFJ31lowBS6zxjtJf1K2ru6g/40cmQ
WrCFq+flBVMPcOZF0WFB2AqAUqNxI6X6PrfcO+eO5PxQRIp5NH7COavWOwhOzbX6
8X03P8lV9K8sowewwypZlA9k1WkKBQpN+vRRkMATAUFP3WKLOzMXHoD0Nh1Kdt1t
5qx0dj5/ytuRexcFchgI8ZCKeR6QSjS7zncTMphP76w43TZzDZJXBk+jxlccxWz3
5jQ93s/nvRAALff1PDVrNOjyK1NrckOOrTEbTQ6ZvxbwuPWmKX2t2zbuIS5B5TB8
ndPvtQaHXOuOqr08ggLmGoW7g+OVHz+9YJN4ekLM9QdkhE3ioAtY9C0BbKGQ9QmC
dM7WeGUuC0DFlSLJaI1RY8VBW5s3AjxiKO212Z/yo32J8El3C8l1al0rBJp6O9dm
ZYBDBOUs3D0KUsjIp22CF3dI3Zxqt3qSkzLiyOAMWvJ2X26XpMvMxsr9tSvHrD1t
2gNefrCb777/Wm6C29qpp1xaLGW5BOvmk0xQiItbRuAd1rAuZm7UtDMrSP8E+8MC
jO0MxPE/SwtVL59rfCB2DwmxHVJ+7csH4i9YHM1Yb+2Geh+0BdnEw0qvSingQdRq
IKUIODijvmnsIpKygVQ5hXv/OcASi2NHmUg3vwYO8ncos3ZXDMRm3YRYQjh8devV
cw+oX17Sl3J/0nn5pN1YlZvcCkh53Q8eZjA6N7+BBIGzn1z8Oj4mMYb73pJW6JL6
nM1LPXM3FBjJPjrTa78ZfBsL0pbnXzKMP75dz/wyXkf0ID3dmXfROUcKtUb6DpKZ
KF2SNMQOBeIga3m+ipV8SVb4ghxq6IMGThMrxbR2jhroRcnnOT4ET2hAoKp1Lgfx
Su0p4Ohn+O9DJOPvjtFgUGkgdkIHvuCkKMF+Kei/vLzgAqTsnjq0mwy6KKLUgr/a
Pv4yZ/jmkMvSzB4e8iU3y7NXnsAPz70rE7VuxdRqkyedQD0EBvrixRxiC7SH3v9W
/H8Cgt3BZGn9aYRLIHxmMtIqdj34BvaJsMg7LFiTRSDxD2ZJc0Gew48iJQjJtPOy
+l+pGi+lFQN+apg5/kTyCIw1NtLuMHBwutFqhsQSNwZgrX2elz/R3h2qY/V9h8QE
VB1cUfH/23VyPB0xXIRybYyu67K36VaOdMscxR3CcMcQJ2pxTObvnLZwgMfqoLe8
PG05ojQzJOsEmQHqx+8x6RoElQlr7I4ofm2WRRdEz4jUs8AOGs3UGq5YRhXRPX2F
adl6M9+zjUjTcSlEoegjzcqJs8eYVE+vbkqv9l6i/cPCdF7XblZeJXceXLkYwdfn
o5L7DBuXHXTysGx3k/qe/ScTmMovOOCzO4oLUB+neHpY8buucmj5Nb7FZKY4Y3P8
gLIEsuaeZMndzqs3I7xgaQ9TVyA31UM1EPvnhsj83uefCcRNuQ7slMivXksxzBdf
9JYEQCuKRjS0aOizOAsoc7K9Vg+MwYabkSs2zksJm61zUUX5neL1CsPzMhiWcQKW
K1KZ2DB20JNr8oDF8ID9cZc3oOg4LorWjbRmTK5BRpOnLf7nUUlulhlZkf1kFFru
XPSQN91H74Cy8MZOx+Y+m3xJ177ahEADfM+xDmf91b8qa5wBYEHarjONOvi1lpZP
GETEw66iIqI22vSm6itkT4xMmgX6REBk9Ydzr9/r85sRxX3YvanKoIZNlsX2luYL
5VJhQ/2HMB6qKo6u7jMzljrSPL9G+zJ+VISN5GW2QkAcR9ngFeurkYRXdtEA+4KO
uf3/FJg+UhRerqNv2Fv/CiJPpPCvWwyXihz5kNe4PFdxJSqdBi3dI/pn1EoMv1hY
0WlOs3sQVg+HeQucDDZDsHJAsKIj5J5MTiWpl0Nb2lJBo+1Mo3xeUe+WToB2rHxm
Bhuppfi6WAmZtO2chXVJAaNq2GDOr+fdW611QaTJrjpzVz/abvE8sdP8HWAr/UkS
wlGZumG4c6u9opSUhFlcI1MuaYk/IE5P1FGezWr23HQZNtODbdo9DPMJ1Ady/6kI
zm6dAoBdbQRvxixsyRyz2qEBbfUfOv0xwLNNVigx5utvvxJzvJjFlGkq3UdIPpgF
G+Nikg65BF3sZEDvpVFNlS6SxRX4NOKhUDxxVw+SfeJaYr6S6FmbitVtLQoRDY08
faBampQoK1SztoeyJVHXT4PYMUFPewO1UYdiVepH5ZbQN7Ouamc+K58Qaj41voZ3
XDdD9tRl+YmDxdfjAVT/82bCYRt9w/LJGKIQSZ11t3kooCJREecDzwEm/6w2MwBJ
rWnl49Zossde80gp9R+dCvnDGjdPDK0n3CJAgy4qi2tLKmqBnaJoCSZJxl0JO2cH
0QHXY1GyG6BzTTgvXSZ8wN1MO5gr5opj3djIOs9X3Wkr2JBJ+FQo5tn8eWLT52+j
pdm7FAjOANlDAfwRXqMnyWYuLf5z6PzyfofDqaFeizvbIvWnyykfnMMFrirfcoA7
ZHQN6fKGWdFPjIGWuxoks4tfhZs0EjI/1PLRPt5o82ShB9fiuxIEvycBkFcV+8JP
CFvX71pHa4kN/uZSz88lVD4okVTGRKXx48UDNZKu5YmrO2X2vNu/1XoRX7lujG0w
1PD3/Z6qrQaM3SiI+RD45bmLUAp4hJnHYWM/qorJusr5M/Z99eJ3srjcZKzt8FNj
wx3CbUMbd0Vc4h+/xgUzuyveRwe/IpHjOO3mvStk1z2pYv2GoV9R4Jjc17swrOEK
rbEGJizORGTXjJx1xz9+DJuDsCDYs+CuNPYsGBpWlZeLmOYSV7i3amiGqpmW+b/e
8boYsOPu2TRMK2TXvILvdWWl6KEfjUHXcBu0uT2hk9227fflXvURck1vUMCZWxpg
ntIWzceZ+mfdGDImp+gXyeCaSnZb8dycIWC4UsF61O20wma+/Fj4GcQAj9dmdDYE
Nw/f2AEoc5mvPsWK75gTukyC98qgoSxnt0949ZdIMsbCDHpf5fa5RRokUeU8d3lg
qeV90gnnD94tmun4agSDIpJ4o52Fkv7cnKJdUBCsx7bdrgU3AeN5xNPoZ2XGd0ys
mAHxg+PexYgLDZMORTe/Xd+GknOlrywsFUihhs4zm8y6AOONHhO3iMerxlTW4375
x4H3SbMQytXkdhFtXCoRR7s8Tby9KqUXiNf9FXeHXPNom9OP9IJom7WjNHD60A/C
+4OO7GCxWs8mBSn7T74M+eQfl8lSRNVQ0Wlo7Oc7qWosedfta/ZmnqB2L7slmLuH
1ffiLQf7IINLV4q1xWbRjNgPjVMVdTwXvShHYZtB1KyGBlszhsuLl6pSovDhtYMO
LtmaVRPBOvOdDYDmxu9meDQr8CXqUEIhgpuP4GIGWtksLvAJv+XiSx1DaCgoizDg
wssZCR5vhVHiVoaEF9i5THE8fTQsYmga/ysoteBluMuhOyAFtdnzbQBerFbnjflP
jxBt4lVAgiEFbOVbkR1GXjNtVbgS+zB5ihxKeVoH5csY6U1Dw+PCHXapzS4WMmp+
uA1jET/aD6FP2yq3hQGkpNEjapZAMw2koZe7er5672bq2qFzWnMiEn6bcNEA7hVf
z8MvTJeTlN5XDzn61t/hHyjWlFXQj+hTz7b6NaLSdG2e8rrG3MxvYO9O24H3o6vW
YP/zyEk/j5jNEVJYWvQ0K9RSHQAiv8Jz6OgrZiMVVVv11tfGVn3GDZvni/zZ3qRw
58RMSDe2Om/ssHZA053F4/t4yMiVXPcCUoejuiyvxDcIwYMWc0/krrLMELwJwpj3
DtK1FafIJsM9LR7JXKVFv/hmxBPnXRrpOWuRlw3GSLp3FToktOXdgiUsmJJmg4VJ
7xmeKII3H6tGNasH3UCinfRNq/LWcYGbXlHoW+n0AF/xzEIh/jTy+Wlu2dPXOUfs
LxeGuG5/3ldsq+TlzuCLLZycBXTlMArC5ApjAEWYTE8tTQvWmWLJrdfFC2cGPZw3
2KOWb2U/Tfd4sSVIKUe51RhHM1qGfw3ZVlrCEtZDTw5FLB34Ed747pTkt7IAuB1l
n5N1w98EUW+wQVwTc1k3ZP9Yi4LEmhler9yiJ05IZWsp4NtCrzc5fG0Z4oTfwhEa
G70S3MajSODvWOOv9CYqElfZt97H0mDwJyN6i2Vi8+CRrKYGSDnl4y2MRNMe3uQc
isKHQtsOyOY06OZRPUfKp2S+EUDl4Ik/C3AaWLGdm5Q3h79OCYXs9ZFsOCC9esdn
svJfidIPW3v9HYPzo5y9+R2ASP+Bh8i75SbjfIieKkGdD3nTXsYK7sPqqYtrWVY5
SpKF0bonJMhEyY/Gx37aiY41ItXu32NGQHCslKls0gB1YNDdNiRzf3eFARFoyksD
pJ2qTcrIomGnki0UIyBSfMKF8nyghsLR2tBBUbwXGJT93+z0bWCzBRSgXe+rSURk
ejEHzl74ricSpLfCqtyxYddI0sb7OTCl68ick8hxXFjz5wo+Rm0OEoeyMXSmwKdL
6N1sPWkw2p4NH+gLrJfp3BkL8jUD6HxG2psCCI7cTmrlJjoKxuZMQOZ3RvOSZPg5
kKdtbNS8+DrEh7IvZYsE0M3uls8mbM7BIh2FNOmR7wkV7VoDO9i3SaRlw1OBwuQU
CZRPDWUJ+WfkNtY0unazKSybK3a54xn0gJ9c+NtPCQhaTF7wzlvj3K6NaQZlh8jS
9Yz0uLsQcmBCo8z91V9Da5CrU75s411NccAEbny5G7MkgOAxHMhSUnUz1xomO6mh
/oUeGkhXnsEzzi+5YBMgbGl1we0QKpZhF9ZydqTJrUyfv9V68HfYg0rtjehIvQKP
WpOw9sUJJxpa10W7I0uw52ScvuTi5SQPolnlXU1Wt+JsXN4bzVpT2XdwEB7ATiPQ
ErX6b74FHhdZqvAHOls7AxtEkBAEmzkaS8aj+NlssQ7yfspKKnhJm47+yrEjj/5F
YcQGoeat1WlwAbR/RXUb3ugbTgG7v0WV8QM0sEBaRIcKT00BeoVOgNK7MR8OsLVS
QutgReeoX24t7mesmC2vYvLAZkJ7hZA/xjtPkif2ol5PYqjpozquKe52jozSyct0
ZSqWnvM5JNP9AHtO8CRruRd3jW9F/hMUcsY/y9vZS3nZeb/Kc+E3wNxx3ieTZZIK
vtENsh4BTerbkS6Oj0AY0DecbtpLa8Z48mhxoYbZGfLnvXh8AjMIs5/68YB4HYKZ
+sS3a/JrBiXKiZce2DUaoXbwd+MV60QHXIoY31ZjP0zZ8EBPk6inu5I8vkrptguN
OaPHPmZEW8fu2eVTUB2XUQz2MAKADFehvAToWA6l7PeX3khisCnCxN/+F5V8yGlv
bAQU/plH5ELdA+I5DP35BDdxOhoIG825yEhviRynx7LiI447BrRKgowWfewbuhkT
aDra61F0cES1OxI5Edox9kFp9nAlslnIU3jHtn9sTA54AG3IvyMHCz8ZVz7CQ0e9
e9D83PupTPBQmdxZcoyFFxbxF+PtHFXgZZVJM5mBQoCil6As11JFuEu3IcPwXyb5
vCZguqCK77z168Yvl862wpMgwwFD+ktLVtCOrFFeJch6i/LI2Y/RQ+hB5+qSoNFS
pevXyKpaG0kSrVnSzuz/5m99FCN5yKoUxclJrySdLLWWTsBroNRE67qbHcUbWEpc
DMh921LhcsC8igRXj0htaiMjp+7fb4/ZPDQ3PzpbU0ajcfRnfQhibW7Rn1D8b2UA
3hM2PKzv30ZbCdEUjlxmjzV+OC3NCk5dM+zFloh1vozi8TkHxTACF7aMzgLXZwgL
xO4w/1oM3TmJpd0eZfOQU7Kx46lJFdT5Y0pqS0lJC8JkPLmyxRfvGWYSb7KfrAy8
ouwn8hlc7W0Ctjse9woRkjeqyPXACZMW4ujNTl6DvW5c/8w/iVsTraCgbI4tM1JE
8zXrVRRbhYgIeo8O4chiVFr0ee9g5oqsFm1h5uE27gV90sv8oaQ1ijhWvspZujXT
xPz85cItRzSyKJHQs0EUEPlyF9apwa3BaQ6XZ7oxIbopLHIz0XB9pn1585ANyX3h
s0X+NORVz2l7YvKcyVletB5xCiPuDWJiRzbwYNtie8E2qQy0sCYiAyxkASXujLO6
GbXWVBnnLmo2k7laetes4i7hHblLF6uMOlKTR49wpv0zxYL/x6jQzL7EwJJ3vcA+
MDA7QIy2V+xR7YJxeQqU5L104PkQFAExzndQJqL9rFE7rDwap/WK3o35Uihkqpbk
9LvM2pNW6Eyi8RFxX7pfefI7RrCPgm1Ktu4kAiKiV0FL/oxqXzGITRtiwGBUD2JW
1Znx0OcayI9KoVgKCpbLf+gXg27mioOFfI3ysaLAmfSECjZuNaAd1BrnuvZt/fy8
GE30zjWgOygMTIMfO8lhJA3nifghEyZPpWXqQlp/DraIHHPXTosFyhEo8+9QXCVy
F26hDGx3+QW+aEf3zkAUBmTqiSInUHLx9b8tCQxQtqZYBhQiHlyet2/WMJPi9rIG
2CYFf/f3CFhrOTfvpNc8overv5fWiAS40z+/adPL8y0q0XUUTz1Rr3xcyQznVyJL
rjHnBpu+veD3t2IlW8ZfWpNAnyQrX6uYbwAIvSblPjWFWxwR20lUCKLzTp6GvI/D
OUGBXBWXRfqVSVtVYb/Ftm0H3IBeOfBUtsztOLucZ3sFMtGEVEWTZKM4WafyJ0RO
N9AGrD8oNoFLQFrrlFfI9yXXyBseufY1nMfzFVrIZh/DmpOM3ECFuK+I8CDAOjJ5
6pL+HAh8HcZEF4x3WDCLwFVuehgRYGffDf0DQdHOJscVK1L1uBwO/75mHueUS9Zg
bI5ZJudkuKbEf+zRliwc+siaftsVqY3Hq9OYp9T9LpQvb7Zf4W/3nZIlL1jiXMkJ
VnoVrqO/uktePe0hZRd0cOk9pRuNipzHhBUbY1eSyvsz3y4ZKexNhyIanz+h2raE
fGnt/xrXNI9nUGXZiSezp3dFgX7xnFRtNUPzBUd724u3wRGKnbPfs65h/KCd4xW1
yJ87dcoUgcRqBxP0LXZaF4fGsC7Hpgz9KGA8pkzcxILLUfIEFQEumZdgV2ZTeGep
NLt1TxNVcRpWk2BR1LZLue9nMsWugPasHcXvxyx9+MxwwTQjO2KiH//Vfa0tBgfS
f3R3Ta0trUyL4oixM+aNkMf3iJJ40Me+mL+g+0rdXBjpejxwLsZr5J9SHvN+Qtrg
lPrAjFJRRlYj1U3t2XRTqa/zbil3sDO/cJ8cGdBRvFhJjW1lECpUm/o+/olCqPtf
e6bx8UVgnsyqaVojdi3T81Dz6giVm1zY4SNsmHkO176ik1893uZFAO+HdFtS/V3T
rqstJ3T/+GR2iNaUcATHnZgbLpNyVW9abmjGlHymQ+VcypO4gL73Wz2MZak8Kxmz
nRt4RjTcjYtyGVrw9/VoH3Y8jH3lHIZWRUbk2r3qfU/Nm/IoJSUPS4Fc8aaRjhX3
rzELdJgCyDKNp8GeASCb/oWmtZCy/WqpnWtQkDz4EHgdHoE6pbOM/8n+W6p8DXEe
idBiF3E3teq7k8TxKYtX3gZ+6GzKA2oK25mvB8dAr0ReQQ06/yQIuI4Yn13KqzOP
CVj00LCVl8T5A5br2vtsacr5XHoza8s66gej4Ry1UgCSUivQX0CPo63XBisfGnDX
ajx/1I5bOyA8vaXLc8YQTfQu46rxJuXGoM4MAn3HwBobmd2PJK8QoMuvfGUopPJK
aBEzxIskynIgNYV+1iKuzpAv9rYhKYa1jLAhueragk71yQsDHspErNFJawdaDut+
5oG9y7xjqSszmhB0714i18dUNDnk7XPwzrtBzO513bqgngb5k0YkijIhwUCXAD8/
OE+P8zED1V5tPD5EbNbffT6+fWy3jC2tpBUy8nYKlj6tZMzqIsQOecqXqYmdTdY3
H+6DAshYJd5tHU1ZjCkA5Zy454rP2zh1Mdf69fv7hOgamipJlKKoIjsLslNA4xqb
dQzymrpKLe0jgPhm7oZgyJEb+MX3XgCb08ByWWea6aMxhMkWMilfnRFGJiDZfV+l
cmj1Dtr+NIw/3T03hOIyxlLfxNtQdoflJFl7GKQJi22IyE5+2MspRzNhEWg9SXXM
Y0YijSKALVWsdB9IVItO5kcu3Kw67upnqxVhJEqePuuI1FT52vtt6y7iM4xiGtCI
EBVTrQ6wytjYbQuxOjrb41KfBT7kKak7+ji+eGMWVTDHrPFgGJnjpnNqnDn3+pl+
DyXnxin+YEVZ6JO/ozVLs7lxEUmzwsQba9TnU0I6jAJEzwQHtbPB2tQJjjbYu3E3
MCi+UPy/6rh4hg6ZW8crYlXIrg8UmiHkYjm9aBoVmL45a207EzB5W1We6WN+Y9JQ
SWGIbQqc7+dIN7DMDVTWBCv/A0WKA4srR5TL/9YK0bXz6/wnVz7kBNvATgKjJnhu
amX8jnZyTNgQc43RIlF8xam1F5mh4l9RACxd+x4AY8UJhmCos/6VqC468afBK08P
ZwnG8Vh6DTy/y8muwbw4R7YZZLXTDWuKlLgxgim0fTAbnM6d9iGV7oyHpX2MW+8K
K8MeGPgnjJSWdkADXdMWSqb7MKL6wnMYdlbknH2rn5GEJgAldtpwr++7nxuUhXo5
mN+eCTyJdfe3eCk1xpvQyfbvIUaXxbu2Ylmx6KpMZIvgpABWy6WX/bWQxG3627ua
fhwX9D9IrxjXIjfRu2J4KDu3g4owLfVdFLKgQ7a513vdg8D+BB+KxRgoUAssZDrv
FWPTVWzD4GpiZlazcveMf4FcY1IA5v2yGqZ2kw+fW8blPQI53Rsmjm1fTnf84n8u
KC0oc63QHo8D83UCWsscP4B+D59FmK9gD6HvkKL4ilQMZ6ISzv4IsI4yNa9j+jr9
Ahl8jw8bN1VzQYnXtz3Prqe+vOtWFTKfXdRnpetj612QSJ7IBmc62uvniqhHdVpq
ae6i+1Euq57JYCEEPtJk7bDOzbjXLeXnzJRTMUl5EZpm1KTSE5IPxjUD7nF4u6KS
bt65U7SVoNcWiy5MblZIUlKAmRHtbC4Czn2W92t/nXYEUaASZTK9SehO2UFxcYRX
GjJdu8e1Ntuda5MgnjYlDcGIX9WHHXqpWiBKQC4SBGYc9vlWNyrBpBfdnu0Etzaq
MpFuc2Y/aui+1x6o6pDljtiFzWCwCTqfNs3aDFbfvfb+BhvWXzFSR73Nh4BSDKz/
h3UDWxXOuf2DPqEjZvdaKeqXY7pojrp83Vjj3KJv5ixttWsG6JnOFZML4lzl3KMy
wBthTN5/S4GOkvVE9XknaUAELNUSjyxG2CVdpHfranCsjnIJCS5ef8NUveEaZ0aI
yq5F5X8k86WtmQjN1zMvJwMYdtgxmtYY5uE2QKJOYAM2456AoRzDDQ2CP3ayWkic
MeeA5LmdeViDo7coScSIHs6eAn4gX12CxpaP0/c/4+BsMTJDazHaoqdI7+dQVfn2
v4lUiVRrd3pCRlO+1siG/0AD5Fily3tTk+9+F0nRKkH7/2HvFXty2vJNBL1EV+b/
jCg1y8/ccV6ZNKdQ1Ea0JULSDZ6chJy6vELZM5/EQc1Db4JuI7CkKe1AqILtis1z
L7/3/ZSE/OloQHKOufzagrmTtq0Kij6EZysxIMQYA74KXbg7eHIyWR0mauRslXwY
k6Alh42Go4VYUycjSmsIMrIXJvx6Mv2x30Qyxx675Toys1T+V6DiWZ76+QxGPyaV
WmqJF3ZGHCWXlH0XSYjoLbL9wR2P4ScmbYJPFNemAAWXG/fUGe7NwgTSGOCfwhDs
31zvDmE5PTQiK6F6z9yeY16yEegz2KakmE0JTL99cVuW4p5xaRbzp0P28jSAxDks
D3IsK4J6m6J5go1ByUmmVeEnM+nnbB7eZAP7cGIvwc3NToFHlUlj+KbNzof3plci
sfw1NJsFpOzlezl2xTel2u7f3+Ss1Rg/ovWZhwng368En8JZ0GYA7LmWowLkcs8I
BDz06oKEq/9lM/MD7Z8ve9FvX1EfX+XTYXPf3uukUwtzpeUQRSynHwVo304E+2VX
M2WvqBJzUIK1paJzUQLu1UKqm3XE6/XJT1ZvOH0lcXuDx48oj7pu67oRCAcTIaB5
wQgWO0UWc2vT8Ho4PPOSrtZNYCM1s0gnn/g/w0Mdda1WlmALFczB/+nZHCjvjw04
udawiv1z46dJoApB8m0+iF/XDjuzIuXQpniO4n56j/+OAGfUIZ/hBRxuSAtiiD+s
PNlN1H594UaRk2bArItxcx5Ljw+ftYxAtRNy4DhTi1mHOERxtkzUU71zYk4GDVEr
fPDAykH6hYjdlM2T4H6D84IQMDNa8kHjnUR1bo59a5fjZimyCZlu1ADrDDlAOSNR
14JPr+jWEFoQN7tMT5KtvHiC0awZ0+D84iSYB2fniz+/algIeZPOozl7DEvIg0BU
lmjUS1pj0w3bA/TNeON2AGwsncURyf7+7tFrfBl7EOOhEejnS0fi7UqbWS/e0rzD
/nuWetDqayE2T1Lo0V1uKgeDfkyJ+Y8xlua9XOEY54LtT5pOxAQRhDGY9wOXPPvu
PThnNZ41nVbQnynAHo382kG7NC+b/7V+TvHg/PWM1YQt210X/MKZx0UYr8SSkp83
GoO3IGA86S7vkgeFjCo2OENMbTOQOyKEa4hbc+rosSAMIBKBd+I/jemOlc/ri0lq
BT4MMgOcMnJ5X2K8hoTbViCwO9kQtiGo4iywxoqYtQBhY9MuV+xcpDEGH6GOMYJt
cYmw9phnI5e9RHqihae1Qo2WKqfLA8+diKWsq0CdZT40szUv2ioHjs6RcZcSupSr
tjBgWsUdCoYYTnJ1HHpeuH1IDbIJOFeyR1+1XqA176OiuISgvNql2XSgTnhPdSKJ
Bl29SBCwEGZtCa4N6bmPoqCguoGwHRajvmCcgBO2md7cm9tDdXxZ+fqk3aURogyH
UblQpttoR9+MACEL26hfkkuywdeQMZ/8WxA2zn6hWW0lbFp1MhVmL5phhsAA8o8H
leStgLq9EpDW5LpTNhwa80wpSh+m2eXrBrNG8Ze5FwiGrMXejEJIUmAXWahvvw+z
bkmTjis+rPDZhwHkvR2zhyowRsx4/fjmIRNOW3Q003u3RPkjMhqkb7yMX1v75TVU
HzeuVEsWyhnaYHcjK3fCAbT2aXCfuPK9rY4iLdre7LjBuG8E2G17BBFEuOr5aUR+
9zM5/qiNeqbZfXCN3iYp2RMjofyQyL3KbTXb+aUqA7/XuRnih20o9wHcMlmdi5Y5
kNIBUzgLT8DgwT2zgmFwjoxWgTYgmEHLOEwHI//pN/E63iumlZ6DSLMpoM2alGV+
0DW6tSONzYxu5w323/NsMuREkDONzJwwrnF6WaZQjW6KiXqxjNj+Nvrasa1E6R64
SraBNBSnU4SGgNAo8teAm6mDKc/gjOEyaDKIJAAd99BStuISkG5j1VwE9yFn2NBT
i7SnJzVV3MgVUE4xzeKkuRhL51wPFJ+zCZ+q+pOJkPcsM9G5+LtRnKIDcPlPUaJI
i30aLX/yhtX7BfPegyIYSAx2lpePqbUwCpk5VZQYNmFGQG5s7GgzpazFXwGv542Y
VQFc80uDA+bzM+xoXIWnfuPY6xULU2FBdSvDaZ4dDU4y9u9FPIP38/bTmMduE03A
I9QH9/VHJT3bOQUL5vMun/ahGZX3JaheDxd8Fq7wuvVFWmRdQ129oqPgL9KPlsLS
VW1yZ37hIMBsTLA0ls3L6Axl0TSI9a4+eBv4SYxnvznd7Z7LZutKQVPxvwNOr6/3
5K8Q2CGv60im1UGdkfo3oYPkMjE1gHjM+kI2Esct6vQULEP5v6+j1Lq19C098GT7
meOiT7PlWJJqwmnF5Nstwm01ArRIh/EpTyVy0l/b6SECLb0I2vjrS/Ie8yay5Slb
xgYhDEVrgfVc0UEbJEqqz0gsJkBa/USTB0ZZjcOOhGA1RZiMCyMN8Df6XFl6ZuWg
HCH6aczsKKqMqn3q3dTwDqG/emteb8zLVDD+ANnO+LgecfRZ40eE+cYbVVFrijFJ
CZjxIatgZfyOCDyY6C+Xkf09hUF2yKkrdxunc+AFzGx8HOpMVOajiivLHKE3jZ9Q
XNTW/FT7Bi8v1pg/lRRxWFX+iErgJAVO2VVFQ0YiKAKHGNJ7ye9I/Uq1tb+ORt4N
oha4d0dn7bNih8aCLR21BOibE4Y5g5c/6GX9cB/EOB0d5Vx6MvLwnY7JBYOh2vam
rofO5n8hWzQF09i1k7vij+jAwo9H8i6ZgKBfXpc//o2evRPd+FSXjGg2R2QhpAj1
+xM2KmigwPo91NbwEHrVpQlS8+sdI2TR4mLEm6ZAxvYWvKad/oICUpcZVwccVbOA
eMR7D1dT1sFO6Y3G1JL1+ZjQ7hsiBzMHzqAOwBC54xag9ig8q7DqIsFieqzp+qhM
0IF0DJZxj8qS/i98Z57AsWmbJvVB4+P4yICGNf29V+AQSEvdiQMGCiZZFQlaOSVm
RA/opZaIQcrxJc8rKKK4RDZpbI76bVND8FQvL7SXXlCCkBRE+goUh0iGPiMyabev
e51ESQacKhazroOIv+M33aJ2P4JsbnLr9mF1diOiEMxTaT9ohrcj30yQmIwlEzKn
aCvCQB95rDG+NX9bEn7H1T/3WyvSjbvHXOtEaKmGkW/Kh+B2+Ldfym+ouxWdpRYW
641XIM/hKSlQxZ/cXLb9I/H7tLAhj5QkORR4B/++OOY6AUvdqk9TLGKfFyQbJS7u
Hj9rCwldEUX1jpHXWgs9LYJfdJ/ia0j7vPs3MYgOszNOQKtq9eSkaQHmfyjt6mRt
Y0k9qHGZSyZsh2VTNiXM2ftQ85Tr9suIvhafrf3RQajUuhQ763yX1R/mJAHdYECA
QQuT6/q6bhYnQR6rBV2jYSV6g2K4BzqJlvnHqOkA7i0v1YQjueV8JyAc8DTuIRNZ
JXaaC+/ZZZEoxsIB9Wz3ITBGVp2IylevAL7NFR+aTMCEnOBJ3os4RWDfMl80Fo3T
K9EvPuqoPOsiIzUYa7lmBxI/2AOiwqNOfWsfZzO2yoaVnG1E2kUkvJ9MYwZY1Hpm
BMqnhtR3oj0p4H0RxbF/iAd+wT2TEikMiqPvLHwWqFwY8rG1AiSfM7Vm1VUm0n0N
hPk11G8vAssU8oihOxlfVc4mah67zPoxkWnZpFOWHZiKrWqUnF3p1MyoBi7WhRbg
Bbn3ckWCf/Larg4ABFr5F0QfMAWVyhJNPEEqVon45WLxSQwbxTwmSxupTaYCxSpG
Tq7IR2pSGmhN5gCy/4BpuGA/qt38gWk+chmX//H+P3gEgnVtIbw4Oq1wxUp7G6MY
7EbEiWZdprpdJXIkIfLLvB8rKix1xHQtXf4gBitb70Gm9/XX2LwGJ7J8azXCPWNO
0mIVk7rYv58Yel7jpCEQqxCOx3Z8i6glkvuH7huvla50R+PJkbJoxAZGWu3+oJPo
dvbnnYYlI+JK0CMMIU3Hi1E1llhZ3iQvWx0720IdJyu+oUvUpf1Je8LJIK9JwsYU
Sv1XBhFmRWbMCPfFj/TdJashIWXleF9iXoMP9/ZYYaXmZBbd+bCcVepiN8J745FD
GnICyBS+Fz+KD2UI6UG7LVcglwssWjxKjFjaKN8wqOgSulVYDLkC5/xMrj93kHPh
RAX5N8jOydB0+oFL8r1+HLwte92C7OokzwrPSBlTOKxJE6ykd8l09yi5pnTqe4t7
a86iIf+03qNE/ndeB+gQJjVcATs/h4VmtqK6YcYruP0OQ97WALHdf7bTlPvoG+q0
zroZYzXWRXNq7gu0a/Nz0g/eFa7Sxyb5I/1TGNeDh90aMro8158TErwzUNP1Vwgc
fWcxHaRp7I2y1kCW61Bk4OJdXBq61hCytTualAF0fArAENLbKaTm9pB45BIbao+R
uOJS2v1LuvuhoYUCu71qRAPwOVm3nWtACkr9Yf0X8M/pfpai48FRiap4Ml3rCpPA
1ZHC8kcYi0/7zfDaNp4gxi/+jOs3wradfw++X7erHh9622sUg9bRX6BkuwB8ScH5
IZXRK1LLA51suyzgZet2exjDGDrhnFw9ddbEmhnXLUXhx8z+EnfiZHJqYrPwV5zQ
I6/du2Ydjge37EEOjEfSxRzVtQmMuthmx9eSQTLYm5h5AobUM92TMPLgXp827VeX
Kw7p59xmfpDlR6Tspl1h7XlxSU7k6vQoDlaNsAs1FLSWzbLvc2PC0emYkCV2FhNp
gLfrzl4cZg2SQyOi+/Ks9t6bN04H/NkM7+5Bpv+6ubqS5TNinvnN1QSh+1TEsJKP
thr9N2SxajtPSf4yGRiuKgjcYl+OEay8e/FlnDCGE+NKBpJipmR8xKgumsF9PBrL
CZffyhzXpdKEUAkwpaH61QUyGaytnDYnIfsYQ2nmCZ8LL5NWmyALlaQ/ET7IKStT
deKXRI8Qb5qbjV6N0leUati4DIWPE5AeNfjIVoY6cwi+wsw2TQAybmLgauZbKzSB
S2IeqGGLKvu0i3PTg8p51Z0/1e9Ct2ImHDlyOJcDA6ulLluRUybPnhScx/Qut6Hr
AyESFoOvgbfWM67TkbTnpHYj2GWwoo2+SbBJOvYkH1WdyO9M4nvyepO1gQuTM6cB
XOqHhD6s44Hb2ih1z7eBQl4CgjXp/xvWW6TudDQsZJLXy68vPZJuWIzp700ilIU9
7w1m+URdj2KvDsjgsWqkeo1Lmefbj0LeTJBKbiLw8j/b6wCz0+GW40EBK9jm1ZoU
kic7Ea3CQ6/+bR7v9vtONvESB0cTjH3mth+SbO0ilkwTeBrzkcG3hmuNKpXPFgpG
TEUTIHARU+shU9gNyDcTTytHI3LK18Z5V640T0WR/ty8aB1e3a8sm9BNcLDq2RIZ
3SxW5IupJ5cDB3MJ0tK+sL2xcVD/Z5SfusdkXIl7yDyiDopk7SI1dxG6YWPfa/Cm
puXTto3RTwerV+BrxFnL40pr2dxr7fGGZqbzvggPG9vWLAvpIp+mQXsGx8N1f8yC
NRryL/R9zg0513gCK8IKS7RLUA4F39qn4LswxDyRI3WeTho6i/8F3hXred+2Oi7i
1L1sp1H4ZyIjsVPGB+hTMEFjfw/f2iUjmJDI3LBE9hJAvNHz08jqTDjoXJpwT6wm
WHum5o1sIfJxVNZNPm5062doiKtag7iEdYgQHzTg0zxtdp+hGHdbBedWqbRPcK1H
KE40pFkxo1cOp9zlV/zFlaznkli1rqa5BeMbVyBtqA9ouU1oogYhtBXO6nM8t6JB
XjmM8sVytZ86X9S2A1vKMQctmOfVHBPztHEitqO1mL2H/HTx/l7NOlFsFyDQA+iq
BF+I20yI/eCOX2HsOsOU5sR7ixbVE85WU2xkDm1oq2tkw/6X+DGYt5KNgqQuIJCv
Z/IGVQlvIlOu0lcGIWKbHFoIz55eJqY3YI7uX+WUCvsJVCR2tYDMKkgSJgIpjwrq
BpA/Ix+aR2hZdGdTvstN4cNqUBWe7WaLxtB4EJU8C4RvS27mKp72/6bC95hrtAGO
X/aah9Ib3TzfusrqjtISlqrUTTVC2GtnREqITKPSl3zOdl5or7xqXDbk3ofebQYv
hWGqvSWiRpTd0jcDCmykH2CfNk5sCBRPXe9JdXiFMHu6CN4zWfGUsh6RrqQSyDxh
jeHfM/SOEKG2fuF1MT0Jh2eu+7iW6po861YyPVpAxy/9jCIweVxgbw6i+ZMQ/z1B
Ch/+1+yYnpmjtyyYxub1Uw52BBlLudX3juN0ZCeNThx1psKNslcPVJb0YYfjBVJS
/moqq+/XGAOTAeIe4SUFI+C8QfGlD76uIkKs7roUvPUatfYnVkxjClauFsuPztJZ
yWdxmdJRAWARE/V26RTvd5c2to/ejmX0o3fhlIQUA8AQ9MP6H/T4vc14wVFy057W
uu8TROXWF9rw9gRI8XoAwDCsIJP1z7DX4NE8Md21HEokkSQrhK4VQUK0L2jrUItI
zN2BTHJcPClFkBB06stU0oDEw3BQ+Z9R1cTj0Qm06qZwUH0gCkIpdmzkZuc23OFe
Xk4HTnC53ZUfjB3nWVLohFn9Z7B970BthMRzGdjs+jPEWOM5q7RXVCibmbqK5JB7
FDuObAS/yFXYzj9FnKtptBf9/Wg5DUCcbwe0CulHh8us7g6pJ0XzdmII+4ZuAYRB
NDZ/eDk/39vossz0JXKkZpVr7l4sZi7Xx49N9E5licHqPe9RnTHjPe6noT0iXKlg
LJ85GQEkIq1ImSwYQVuPWMmSOpOD/KAsE25qi2B7DxOcuoPr8I552wF4emZhAGWe
AKhbqOzZk1cfAv5qQ6XiY+FS0P4nPRwgD22dOsnHwQNQ5KpYv8AF4XtFZGWkYZiI
5kqtBE00X7Q21Xlb+T48p26OmYC9RVqYXKJM1ETsI8pvhtwMFn9w9LQWK6JtPmlw
/wwe7e3JG2//4RrpvNzAEPqUMmycdIOhGOgOE2ZJ6ovjYGBapGizWa4LBWr6gdIt
9FFYhYcGxQVEmRaOJOMO+tu6pfq4wzy8tN6iHW66vsSGinqC2HxosQ0gIRxJGdNq
vA9k+FDqtPKjje0ZGBtDSqPGdSXw+Xd4g3vYrK+Z1tbYPIQhapotFw0ja8fu+tPI
RSY+uGbBH4H4bgMU8hz5Y7iV7cqpRdoswABH/vaM0NnQNRDaA9A1w99GATFkel33
zbZzkrL2/lrdNH6fteqz+7jXdUHJ4vME6t/e6XU8D6xWGBQjXXXFu+VRZxYpkRnB
w80SfrpvVkRQ9TwwV9/rxMKTljgpbG3x2ou4/+vmDRt4w81s9IzAvpf+tZpQ9D8b
uVgSm8Ou4C9RV3CI+XQc8G7x3iePHworeET7mU7GdXnob6CGK27WpsIzf9j3xPzO
/4+TMZ2L6Bgn5ZPBuIwhvi1neY64thcRcf7khKUDUzR+47AN4nAL6+6yAKfZghc7
QiqJ12dKVkZ/MXejiqKL3x+3kLV1DpZcP3wyRkH9jVKekSkg4NeIeL/GBoTOB3uL
5w9cYkRxYgzCLyy0f2iuKuTpHddtduWn3glL01/gzCESDoAEOaSyFcEpPahHSIRs
hNR4mY52vUdbIcOUzSAKiOMxF4thUukl3yqSpvMH2oK4MeQdUWuT09vQQqDMm4gK
UtTy5aaR79hsCKjQDPE699LQibC7rfPrSa3cpvr7WdLpvtXzQi5V7FQpQ2gMXCcr
fhUUOHYOP6gUfE499aYAGwOyfpp6dd7hviJ9Pksh51Tj+2g/lk036hmJk0TX1qNt
Xn4kL0VhKUakg9rtltjlYYAXV5x2nHn5jnd+nvT0rhURJ7DSlIUYGMo3gaqJ0H19
2LJez2AA8YDS+micQI5xXMP2pLeeO2T2EcpJmGZ7TPz9G9rwe2UubwthcuO7RepH
LEZ5ACHsOgTAL76gBqKcS1cVgVT3lQf/iNQJQtFbX4aeG9bAYV93nDhFdbs7KYul
KyK4PG5XL8EE/KE75lnB65oGThTtVnkhWl/wQ5xJ54ssmh/mLfobeKehyh6XhAnO
YndsKCBp9HdW9w7LikcWRveHtJ1ulkVKw0JHzVD1vpoe3xAAf6eDOd6xpQnOlV3+
gV6Pc6/ouv0ap6mrIHmYb8OIvfmSMww1/nAOh/tqUtNHZyX2mlyvM94AH295EHsa
ks8p3EfUVDqiYvUMov1IYaM4MTJC9Zxjn2J6a7rVeAYICiML1AavgjSypPJDki1e
T/u2XQzsYQ/gEJIvxBxsb/QNs/8uaiyHIyXlZYVarOq2eehrHdmyPifzE8kFNksL
mBpSjd36u8aIo/2gW4YsNIgEX4ptqeMLoP7Q0z+2kRybzXGGHq4ThBvS5cY1o27t
rhK8n9WbpPWRKKqPNzqjAWD19HOudApoWioEcHdzwQ4CyIwRpa6LIRfdtVuKbLoT
2r4djVbbMjJiqO5MZhsWRaorrpSxVHK1qZl8UPy3DXo10Orz5Cq064GtYp6Zc/1G
2Rt5/4lwFcSAbIs3hCO6un9/oDwZID7eD5Xn//TnRkcbz6T58q0AkERse98bC5Q4
xYWwgVjp8xrO6WVAk5NeYoispu8jCQJaSt8ipKGx9Z8gBJ50KiKA39AfMYt/YdIR
0EjpFku8Kurl7kWow8velOTKZxtnOFdr8OAiXbL62jwiFoySPLPh6tDJjuzsVgnL
sGjEkAKCTSb6SOsEeNHrk1PyIt+jOGsmt+I1WvRTS44tLF0e+QiQP/IH8tx5iZHa
5F39PuG3H0r9Q/aqMrmpaz725wL2FjxUtnGW1Z3EaE6WnJUrYvTc/CJeLsF0zWqn
IiKSBTMG+qiMDWlTUNf/XAmLyJ4IU3nbNzE0r5eBPIJ5e21Rdh6g4cvL048bX1Ov
GS8Zuu0FPFHN+VnuJ7jaOaLKAQ1XR61o40g0GrLXqAjoEpzfrLV0UaJ9JGSPbcuq
jgaILbwJ59e4dbw6azI4NtTy3/BgRXJFyz2vLqOFFDsaT/vQghUPkFov/uS0dFxO
p87eU/nYS5d8uhcRSyx9x83+hAY18TtFjJJ9aNWJVZQjSI42npRp30FGGHMOPWMP
CxLvUfWQQ7f91JfqxFLdmJNPyBWwnVy8m8orkqurFfNUGnXaQLgyueRLy+wF4qZP
FMnazREfSb9p6gBrPzkfV/bvf9RF4fU40u+55FTr6jlkiSdTnohRqhUvDsLbhUK4
bFv9jZ698iGLssngPMa7Grl5H8ouy6DhMN/n9OGxkgeyD4TkisECuEDLMjSQcqp+
48DXt3Q9Lwa81yvMrpmGI/NpoaDoRFaWR10Q83wn9oAmrtVPBSprgEhsS+YQyQDK
ftzy/FWNifaZRLNTEUXzHmO0Y1YJEYsFBXlDmp2Fcuzv6xYq5RpT1WPstyM4/xGr
htJcZqzSMqkawlNBUTNOLWaqn5nbtixdjv3T0DFA32IplNNJ5Q66buJo30McekhB
dzn1+qNy2J9Kqg6gglfiGpLwB9g50lpqK6rY4kSIovSFaZTJUMUqIdkglQxb9Haw
gfyAVjwTB+vzoXi+SJ6OcU4g8sajv5FhFiQ1MCS6JiTtkkCLmu8cY0Qqt/BixDWo
jzGEiX7qSWm7zSpwbhOzLdDFtpH4pvCqcalRmz1vqAmkaxjmAZqyquoSj4He5R92
owWKQNFjR609J3siKVI+IZ6gXEVXWI7POUw//sG1Z65g1EmoBaQ7ZTAKleRqCpPz
op0IcPn5CMOysPn2vmQKegLsOE5R87c0AHaJIPAONyGDrnwtoFFdyo4dR4la8n7M
oP0Q/DrEFd4A7OpDtq0YpgP6SXczqvLerAhDTPlsR+D7P8l4voOoY9AEEM7vx2Dq
M2iU16d9woFhQXV9pZfTaLrMlvUu7unRvw7d/YlMku3kYU5FQ97PguZSyZpI7ZSr
+cK0HNoruQdI2WLeATXCX8X/pWIhe6vg+nFjBfR8XStbei47TUBXrGiroEYVozM/
gLlvcMonmqEar98GQq+Qv+/NxnqUsyQ7Y4J/rO+QcN7261OjdTPLSCz1P8nmMoot
KgrotcesuoFg4dKiB63XLKbrKebOcxAvi8WQhbHpqTYMCT0EtPltRxo7VkcCgoRx
NSkPDK1T5Dx20h5RCCayC4Zi9GjRD/mC9+NYV8bLs1OvH+l/MHm+Nq+vLb42x+Mn
yC5zEzH6L5EbsF9bry+mHtL4gRAaXCCJaAgvoMZAyrp6Pmc4M3iED2KI2ecfX+vU
RD6MEd6Pyjs1rkepQMzq+UyzzRJgJYgQsZDKP5MNGMPJC7dlAjvfCmRYqCms4hiK
BnE3CEV4a+ixCWJmLlEx0fy/mzTQMrFuQ+zo/Q6/K79d9blDMPruPgC3MpsdMWNB
3J8nb2lCdoFTDCF6oiudiPChFNOfkh0BMoKAqOfg1cfZo9UMfpAOXZfMg4ilPsFc
9XG+JPWZcbTW7X9CP2MedTzsX8OB0Y206vGF6X6WwDiu0CqfSdTJMSQ6v9sb3kfF
GecNn9xeEzU1EsjhCwx0EIzz/Mrm7dqJ/djfwcBDUOujYFhvjCuZDnmCz+uWxeRL
DM9HE2EcJMmMNDRU2QPYAy8I/Uw5t0yeB/NA1VOlvd+gjcyMgLoKecMngp13ISHQ
RXcPSY+pvBLQkdVer+7ASe4ciKw3qauyoTpntgkWbwdxMoNLj2LGtLC3p1CtKyf/
jTKQV7fS/6MBw1OYTPWqKHbfItazcNvf60uTJJlZH/VBbiZRLzvO5eUv/v/JbyLg
Hndy+0G3fxoetDSHY+thYYJIEq3unYEhRFdI+czaBWlhkVnm0RdLAUH5BTS9yYQy
zhjVmcjyz67kdpW7LpnRXZ+VKo3g5W8dKi2zpl4V8U9Vkaav3qpPnIj6DKE3wf71
kofT7IwNhauErwjJjdnPYG1qdmZnZZ2kbPh0w+Z4qvwBFNZU9JaSM6cRki/FmEMM
dXS5bwWoJI85I0tSPVoknbVQG7nmkKis70g00nW+SN6ebl+MajO2WHrxc1MoP8Yr
sj1CqqDOp/m2XIHOHA1jyXdSWZXJdxJpDTT4FkUsbENQkfTmlnKs26pPPhfqgh0G
r5hUlCfYh84+IJd4wGJxhBYiv3VdSovRWhcY+xF+YWsBAuL5NubBtXWjlaNgAXtM
k63xCGtIZ/3eb070MqdF20ouURd/I8y/AMbXrJ71gji9h97cbjM8rLAbeU04Q7lv
BkDuJsaYK4KLwtVFQfppd1L8IHXd147jboudGC2OuVBPP7L+kRkJObB+tC8EP6wU
Sjv9vLAwY35jadP8p9R3WktusgDi85chx0quQ4p8rpMM4vKjO2g3L0iK0+uKk0Fj
57XxEgKuiWDatbsJiS1EmQmdxu1v5ILFJn+G5BT73hdAjucJt+yo/T9+TfEmGwjZ
iMsXIcJp7NxBM5a4Ijeb260YTKU9zlhnG1WKH97GmyTEciRSlDmXTKza+29NuNGc
iFfUeyb/71QIYr9X64+GzjeTFwHjD8FqeISrsb4mdV2An5stsq+TG7eT07n80pV9
/rar3/jcaxawvGoNl0CF3sHboCnlvMyrujd841zUUirhE52LJ6IDGXBRBJRT0nV3
DBHg5d6Q5kgN9Mzm0TMM1nDefpIiHrd6AAfm/Nvu17BDThiaJMgUIDFoWwbyGhrn
fjilAO76CWn/igLbhDDzTGNzs82FCPlABFdSmBl0atsclUzu+v8gJunt4Uwfu1/t
Tn4QENh0i87AndYAoQwb4JSBRZmzAHfWJeSd+sqancD6uucFsqUbA6otPoekJG6l
Wsd1SGxn+nbaWhlPrUXedlCy0JGi3/BRD6R7/3juU/uZzW425cRdai8Qn8/OPn9Y
B863h2Y//5baAK77XkFueUj1Nlyp/M19A91m5IekxM1/AgG3LI6mZh01wdXKts/v
igiN2iY9UISHVO2A41zKYH1Jmm2QKcPcApXHQdDawZpnyGRtrSmpZPdw0iADYqd/
IxmP/EwOmUXnTZ6ImV8u6Fpg9zKeESEiq7o5PU0XjXUXewFWpW5uiAyktPyJCHil
FGzXbCYG9MltMpEQl9YU+hlwL3UU7tjjFsHU1xBq/8VS2rh2Rme/ui9C6PvG4pQ1
3E9K6TT1CpnDaE7igo5sP5D4bv14p0lxQ1H9NCc7FMUuXo54rWXqhb4eriOtqjoZ
9m6Dtdd4vkqnT74cdq0nZh0H/0zJEV5/Xs0pxD7a/QaryANFBQc6/ghm/M/GJp2r
qE3pH/rt0O8cMfjHkcnCwAVMU/HGD/spwxGnnuen6KylCKsV+d8WqHxxJRRw+QZU
CiWDQsh/N+x1r4vGFEj4KW5sA5TOGMFi9ebeyRZ9FgW88sTj7m9HLUrf7WSusBxm
y1q34Y7SmhVq7z0TTk0HiF0I7s9y57mfwargFlNZItDYD8Pv840I2uqne1iRNqZO
l9/vyY5Ma7wWdK72VSFzc3u1deIhHypaJMrnE76JdjbP43fW5KXzQdGZYb8i1Cm6
FWtO2fcr/Ab6UPesMbIDrsuu4sVAU5SixtEJ3DNyDZRgPOEa5HyREAXHGmgrHQ4N
QyH3qtqir+JzsCJd0bbdDh/5IXGfNvYsB7hMARdw0E9lBYdjVDo/koVdCl41NouG
6MrU2RtVfpxnVmqdYOEtghgLCc0S/J0WJFHCHjKAA3WTMq8FQZpJh1xXzGdIKl0H
HqVwZoGN5rBmqknAsfRNlz90i82sWNc8rt6XPNtgYWw4Sz2R++u+4cfthWPHp6I1
N1Dq5u3RSh7e7KeGQQf7ZOm3KD26+e95B1QdD67VDUHUnI29NDQajbL4OelHRnFD
pMK2xCr7MMbPLPIEcoM2ze7KM8KIW+ex9lecdxjKQX8eNp6X+cgZm4YaVWLPGVey
GzHJBX/pALcAH1GzjZm3mzN02eiIM5dFTQI7zvhez6hGTPTLj/2OAzprhW/GGich
vPFSTTE2j8hd36p5aMrEwn3/vLcV2nxd7m2e5Ai5srEfOT0+71ysjkgI3Un5kazX
9S6+AdDqattfrKJERUDVVqgOGUK1IXTY/HFRlLVUsGsHPuVq9+I/fXhqCqAVlAOj
TjxH8bvY0XHdX9egFX0KJnF8IHB8ssPNjB4YE3RDPp7vGuULr0ZWOsEFCwCqAV3U
p88FRlwY0q/hj9wkGT9fNTOIuU79UuJ4AZdnNrNeQVDSqG4v7zlIoUWT6YjlZ8hD
Y9az0Rno2Hso1GFb6uI2nODI6YmM1cfBGSf6Oxy1CU8pdE9Z+Vn7ZjgladuOt51t
Y9sZuFrl5koOt8IhZK5AQzuzjKrNmB7HbBvqvuHhfH4cvZzZCji3Up9CAsfDRDB3
qGDaWpMvsk83Vk5xE2Ne81orPGSBXxnmcVQKCp4q01YsLNzhhBINQmXg4LDRq+xj
pYlb+RjzK1qWWC3+EL7n0Xwxw+jtBwObGis8eYGHFt8YNu+Zva4gLoutLJA+fDIF
5MyG51Exg3Oc6g5yY8BsTRQnlQ2ykzMDM1c34aUqG6mtJsWNh+Bd2iTivdi67RiS
tnsNsTkODObTWnXLYdsRQGOLxNpP/wCXspRQhfWbBo573gJ0WFiL4hJahk3/WDEo
130jh2LiOBE0XJg13HFbiK2EeFwtChSC/Rt46/sGlf90LEpZDo1qqlTaxXMRZUo6
XH3MIXkLlmKIn+KQc2/aVjiw1SDErweIgYrD9/WIRKlK3AZ1YP7oGQ1RSr7iKLjB
BIs4pITEaOdT/3Z3nY3vNOOngY/x1YNr93BadCdsbR2088lLo+Hwdh5jBFLmG2O8
OuSMS4S6sfuA7SCbh87AjrVKeoJ9uZ0sx/h28GiyHM7EzUIXYGaW9DOiT+2tvg/Q
Q14begl63uwuEtaKLh2FQ/zINfVeqxAoHxNjhvzbGyCWsDnEOUrnLK8AHxs3pUvj
EjyPqu+teC21c5TgBzWZUxb0F6GJeFPNGpK+KuweCdYDGE9x7F4w4XtZa6w7LW9f
HmNgysth+07XBaHGEpqIuQtGIY1rijjqwR2y9250pOCUoLlT+WyWB4RSEQ4F/620
4SNK/KKbKUr70IfWk1ILooxlbvpJ+wiXK1grXDLN20+KHVcmEU1Ymk5DsMPQ83fz
8sPAI4MxofSc9pG8Gk1aE7y1YUdg1GHDeOw6UqwVlgBFPru5zhSz3eh3IcD3pq39
vSH0Vi5yrWP4M20JyLejGcSjq2G3/T8Pz81mNABXtdEckwW/f7mD/qwjw20sCe6y
j+9irbNy+xIpitHG4sBFq3oGfktElCTRR4Ev5FVP3Sn6qYdGgw4DE0j68ZQ7sGi3
7EQynSYbjgsBywqX2/WGwcDGwbIqwbVpX2Y5tktm2esf9iD5t+xkeYfjVIgrEHid
c8kHxtPBM0tzXkBdIVfdx3EsQbX3z13ZwSH+vZziC/bmYejXpLNVBBkh/lq4JHaP
USAa5ZDhA20iLN1NzregFEFBmUnLaI19Ed0VapoktfdmoCCrrGNVKWIotgMDgCvx
v0ncquWnsW5AOvYKTE9uMZRBPqW8/8e7pjtlKluJCKdqvM0soP+UNEyD3xD3iz5a
NLzV/Rfua+pQEqOECTHgz2aMNS7p4ZxVbZbfSqFyAwvCyI00M0Vmj1GVP/kV9Roz
syrm1OqLwCI3sd/Uu9IlLH6vMw1o/ypMkQ8bfNRxQ/mQLKOJ291tO/NYzjFwuHsP
w5o3PgY7P4WOLZmHV/5LS82XLF5aJMhPUtQnQw66FTgw/bZDTewTIftlcUP74B3L
ZfLTNurlz2VaEd7Fu5Fy46+4hImI9PWuxYvUfd2jsHPXO462empsriRJtvjCrm/b
Wd9W7no0n6uNGZaTRtN9J7o32/RbnTmaflURo6yqKysksJJwnY7JyGFepgSa+Y79
DazwaeHftjvOjYvR/SB2TQf6OgtnKcF6/YPysk6q7QeA9nnvKzaj9w+onzv7SjRC
hy+XrAFvUQvN3ZkqwdtWJHWhTABRt2TFzM/a55T9tVQ7+Z05LDReh0Nra6g2Ufqa
1AFhdTJ1doqCPS60IGJBxEGlx7dKF+jIzd+2qQ1L4oJ7E6Ch9bmCJGFHkwNhsTU0
Mdlx1eSB6IUzby4z6/IDEf+wG+6DoO3YvX7W1BvTrgu9rhTYdVA+7TdP0eCsB1wS
AVPHC1Z+cB6CmPMki5DkiyAa0PRRNurDlpnzR7HSolWm0HnqThG9Dwl41gmshurG
tDkyg8L4vGEBza9Tsk7duW6nbbrJcxlPL8VpLh+GSdhlSEImxgzvo60JejdsXaC7
Iufv/2S10tAcWOmtf1WxwrOm8dDWFSgeF1e2NojHDtwzfeIE77uacaOyfaEBNbAo
XsU4s9Fybei+8q45sZRSSQe9ouBVmTeEDJYgnKjYrEeDPaGb1chEWDUKN/ChXp32
3gg9L2Q3k6z3X/g4X2nCC5WjB2N0GbzGCTY+70lu5kIN+86Ez/AzPn2QNa4Y26fd
QqYGfViG0OWrrd21um4ZVTMqcY37/hfiFVr8tE54/aDMRFl7TM2ca+/6XhLT03Zu
RJsb0ZB3TO5xgmpMtHQBDG9bTO76qnkRbGyyF5eihpBSLwThki6eNcMBb1WLIakD
uiU6HaurjZke54gZpOF6lo+JMU8V4Pq6mnEQyTT9XdnU5ATSAWDpqxBrzzlxVuBK
XT5hhIYSBon6WSSMGigse4wIKzvHrb0sc0N5oITPQapMH7RCW2pPFP8dRk6+wWYL
VUVAYa4HYoV0FFMzmOkEr3TnLtGg0uO6BTASrigzBJknGMUSisG2MINkul/i4V1W
uf6zUtNIhmSQe2KnaudHPb8qm0DZkddLC0rmsXixjgr9yWPLDMi81xb04ok+Y5xL
SWg0wHU+4CrwvwKJBO40098AI1OJ0OnSUJDb2G2HpvPpXmvLGlABxTf/OLGheKUU
XAcTA32CTXoJkkufZ4roOxPS8rLXdEweIp4i26kXsvVFJ2hOYzDGWOKm6+wnyTiO
sW9NS9dbcn5//aJ2iNADgsYXNOs3fdsTi4/jILhwicmOqgcND8pQ6qyBWUWc3dGd
EXzdiX0o5O1DBueMPXp5jdhC4BDuo7TTL/vq3BOIaSyN+NY9NcipeQ22RuxTtXM7
VW9dw6g7pvA4N5c/eGM6IhIzKH+5GyiTu/AWjJpMRwDYUdRgol9hb9xQOje44aRG
s5BUeDsDH70ZZU2p2UYpQ73hzkp1F+JzvSubDIRLQyi9IoWu9sR64/F2KisEil3K
pkpYJexIEckdSAJSAqHM5240RBfDNOEe80mcUOTnpbv1dQbYWZA60+eLerXhArYu
Y/ohPkpskw9G45oMvg3FCdA/1dFWzMYdmRHITsjtQCLEyJDiXbaj0AJldiz0CYAE
H0Soc0lh05N5okWIyWjp5AqerMPCuktzWlPMDdidpKSBtRUBIGjrt6gaIS0d/P34
77z2CsB3S+eOAAf2Ia2wfcP6iVFJq/LcB5bVnp95r+V8tUu4smT0zaqB8YrRxLdu
gWZDem7O5hk3fkn5rhr4eWOybaScfhMkMreUFlJpbnpLvp/FkLp/Ol+Xt4tg1HkH
HRBjqchfqQXs4hhhTen77OCkVZuKASkEOqPmvxOHqy0AgZPVC7LkgiagWQUB3P8C
XoDiDECEQUYXJVT+NyY74JKHpo4ASO5Dpta2yQFzuhXfO64rtKoSo9PKx1ufEnFb
hsLzSxy00Y9rNyTE9kxy8omFnPAYdAStghDw3A/LmwxtN8uOe0S/ateeierE0uNR
ciL1LM59AlV0j9RlZ4n9tVG3aNUy5577wF85N/cIF4fLiFvn2zN2lmhUALr2os7Z
CFm1eSXDkKDoVvCULJ4tgmBcNACS+z2miCqMufXwQihroiWCCl6rbo/DQ1lnLXtr
8b5W86ZVqpjTzCXsUS4rnRMSDcVH1fHdFt4EI1hBFMYLVuiAJfX2B2EemFqdXLkF
6TUTscc5XXCTY8SvszGt4zcXJyBx9ojIL8FxB46WOqeN/3lFhSQ6eQGKJnq8h9cO
lBRz0IBZRvygqsjX/0z/5YVyaxsH+3kZ7wnzQG5i7fDKdJ53esHHaobHB0C0hPkU
CwmPM0EtG26tJaoY2PiqZerfAGZW3CqAMCVktvlBJEaVK1EXtKI+yzOJQP0UXVX1
6pTBtqrvHWGfX8VqgN4E/jyl5OsvGW4R2mzQ0FGLV+66L0XOXD0O623us5uQGhdV
1ydthQYncLbGbbrjs0wqs5LB83sYaz1/Br/GjKGtP3ov4aA+RwAxJvkfqdgUVMCG
eKrqZjnrJlpK/a2B8LNPPyWRejsy6u+VDUetX6Azv3+o8WzwicEkMvZEnnPBqmK8
mDhyIJWgN5q9hzyVtFQ8qVLaOLtnHSGuywMS83AhXBNXvwQE8g4qoPZAUE0sFrFE
qVFucimmPw0u+jMh8rUDcBdHUPQNjGPINu/TE+fX/khsJNJoymo+J3xQWWDANXpi
RZ81G1mZULM+OQHMbxiTwpbVW+ByowFMOiO1jLPxmpurVdF5IJhwuo0izzcZ9XJT
kiX4PXU5dNPKu9mWxXeSQP9LjOw1vCPjJvMUqxGLSuDx0JN8sxWvT6BdgQIZl01r
iKTBbB9kRnndeu69SqFsrSrJcN4fAinTqVATMubCD3T4dmBNx3jCvZ8FFsWT41vN
TMcDAtl7CJvgimGszdt9nr+01xEZje+PELYpGMrpXypiIJGI8GRmpQMK9LGOPIBj
XrhheHqBVqqBqO8vK7JY2ZwYpFnU022PzJgHPcFuYtXF8YIrsPDV+qx9q1Gu/WbA
xbQyoicZHCkl4EdWwwWiCs6swPEWpPA44mp+ypXkc0PCjeB8kdb3eCMta1P4G2kW
Jm92ieN9TjA4pkASRml+ao+pev1qnHFqMbQvwedq4y7VrHDzlaAzuZpmr+7CM1oH
lo6TKF8QPJTI/oa3rTzhUERVxfXr8xhvzxT3jzlCIhwm6CMxjJz4pMRZ56DZ4vvB
9cLFReQ7ujSZ7FjW0gel1CTf5VT9yOy7FwMLnmF6grdWea1erY0r1EoFLO4aAX6c
p89bkcTz8z8/gW44GMeaemeJIpIUHekx3b6CsSTN9ez+BVol20YhX4xz1DvsbZS1
p/l2ixj5RCot6xq4bMnu8XQUHpjr0sISUof7ija6CS0st6OswMHv84NfGFbFVZ5E
O9Z5Mf8cX5Iis7zVHfgim5Q9zNjC7cL3CVKVfW2z1zHnyi1WMGTHPak6xMArVeHc
J0iKhwk2kTUeF7RvGgvsT3JZWm/jyBO6wovjMePBVwduKNxn1bOsQtNC/VR9kqSp
BW0DDJkX4OwT7ao/fXaCPhvYKMm378p7BujkEJJhq3Zgr7+cXKNy5C4f1orts6Am
C9EFbvmS/wAFsFdtQc+IN/yPrFGSUTmjLv2MJZf+EMecodols9jBmoKaNcGKd/Ls
mnNSP6ySMx9BeG34hay9fWq90ipR9tUlwjp12dZFFizPo3jhBGhsGxePnCtUAQiE
UzK3U7VktiBv+LskIGCBQfEliH4tznAMkOkjoVbhLQgYykUziVeyoTZETHUmxdve
V+Riyl6aE0KE/fE4gDH4M8wV3ialzFDIKel0btlMU1fAh59b0sHNeQn4JztPphn8
I+LZwYYMe4vxWwy9dpd8INVeTbCgUzkxsuaU4vvtoFy9XAu81ccodek1+waBe9J1
eeCWV319ahOTZLiZhEVrioBqRvjCSI9TysY7Td6xKZzF4pWn8Or4rj3uxbtsbNhR
NkidmVHgOMCQ85jlKFJZBeYByhREFnDmUDj5nRSj9bA9spwuK5PBw7VHLfrvHgqs
CXYq3F7wih362MzuYIwMu0PmG0uqQO4OSDToRxyeJNfShdkyayXJBkk3fwNEevM3
l8ggCWeagvfr+pVQNEp8shQDNpmcPO3jlvtoMjMDUIEvOoNvLkSPhx6evV6H/Iu9
JcqVVzC9JeGV8+zARKqYLKiz5N1Kq8mgq2pIXkrqkTNn/xM99ZbjO4yWg+4Z5UjT
kYbQ26jWl+9XQ07nm7An26kHtT7YQpabZ8B4psgryfONHFKTuIQjLRPhDG/P8JFD
2wUjwoR+mxJx0z0lIL3+fmzbKPicRsiotMf1MswiUEyBrS6sCaBczVKfuFXavuN4
Fazm4s/afLIEMWvxlsGQxAHYX5uzUuhagCmRqrBFg5ofYuyS/h1xDmX0paRJgXBZ
w909i4qkPu0e20qowFozunSHMfxkkmWHdcAGyktvo0tdE7msb1VASoUn9B2F0EAw
EP0DxdGepD5wKQBjrn2BJZd13/Dixm02IUfwjFujGf7OSnvEKbQnVplw1XZLobpR
c/bDtFX8vWs4n1oyU2LZ9PuGdZPLwkVY0KGS2V25zedwI238fr+czt71Us3thEVj
gee6bat4pGM4JitYPrXNc7rIMOqC9+Dvz8JmlwxlAfkX6vXukCweafucSdGA4NOP
1Urae0YK6go4/fbKKsKCQ6Fn9YofeeHkOu8r+ycDV5E5i+jpXmxUe5GaLx/Uzzd1
S13lUKw+wBeiTI4uhXgmmKvJ3s9IFPvdsUpUdwoSd2HSWfucyGXHvPcCiY5dJ4XD
P0bP73f73VbuNBYrazUpsiYVY3lfe2F23i1u4tb+vxYLS8oarF1pKztSfiJ7ojs5
7/aQR4/KRQw057Rzpw6SmSNMV/dL1XRKbd+BJgMZsyrSbfD+JOcywdxnob5jWrnj
3zoLPSYkIFWdaL6fIexCMZRXU3z6uOkfxm+9ucMingmLf70qC0gek34RHGMi3XJ2
EDtMcsVJ9eEb2oQyu2zgafMPJpW+3bs+dq6KBbz+siIRxsd3svBSOyqsarD/gvbX
iEZDFMRGvesNx3tT2EOb26hfvzAJXShNSwmLUUv2fN3BBshOpXuzi1itUf1wt8eP
aqxY7RgGp93qfUIxMDJN1hKBtynlDXWcbpWsiUaqAp0eatPgixf4hyshzI4/H2Ht
jlieUhf0LfxJ1HxsOl9DzIg3FQIeHPoue4fqFGpYgRfTwQxY5+lAUjbUX+dkaKgd
tgKPla3denzUJRYPb2hwtLluf7g0fbZqPr9u+3eWpLEZi1g6qZpacugbJ0TZrhFd
iXaYTdT8udJKANdA9ZFNO1lVNgwa8u97puspJWjkHdEz/h0QxJwOx2Xdl2KK1LC3
Dvlb9l05h/pbGjZTDLeLv3kd+S9LmH6Nggr0oHvNJDtGiUnA0N1Lok1VKNrWc9SM
r3KVCymtM6FtTg8R/V+gVwZ/pY395O63dmBEotn4Hqc0CK2iml4oFexlSDyPDUFe
Wt+nIYuRPbMjHpc1U1dMgGOl8ryUY3fSwCPjOfJlXSAS5XK0FCOR1jV6jSswyPC8
DHqjJ+WOBhxrYowjdkyxbCbwva5JLoaBOrShWFgOwK1QxCU7W0o4FoVpyxfAHtBO
E5zi5uBCGrtgIh9Yf9kwRFwgNw3qzACS02KSNWbzfsxrPPe8hHf9wZk70MGmZRXU
TYZFUc84NEXpFNHlj87ZW6Jy1uEaslm/Xnd25yiNwNNonjaYleCci1p91eBuvM89
8KHDzgQ6SdOb09QFX3+SwRHyGNxLvDST7txNFvxktR9GzSlWfGx24NL1Bpymgpy6
znFxRXhWdIoZfDErlr5tkFrQuzekGIgoH+q8WUXA+TxFCa3s3jlRalMaaXj9JRe3
7fwCBPHxmD1z1o4rJreB4bUTZW4CSkN5t509mT72BHKKfaNhcmIP+Kxy1sMev9S6
DnlmRq2f3v5nnX+HBUwaVjy2sEsSGFLtYlKMuPGJFi/qsSpTimqNKQ+wPny5bYWL
5hXzL23C5FE8YelzHiCT85TA/7OohgndO2rJYlovtAyhhI6kXiM6wEj8X435Usta
Q74jRMQNqUiB0Cjwm5tFm6eANgjR/2snj5omSGw4cSarH+xIm+SumWm4uYEI0o0L
EaPMM7yV53tU6NAocExC6V8Dj2AgmmSwhwsPrj+7CyzU1HVHqmxFRukQorzfcnnK
I1CWhMIryC9whvVTMhxZJcIcJZZ9wCDYzmQKyW2WJIJr9esR92bt/5FhJRVJ/aQ5
EXs4FSjyprD18M4IYyARx2oAWFx2PBc9Cr+ltaZ8yVyxBzUEIl9V8Qe8KGry18QQ
sxLO8q/zsDxrMh+bs0AsCdd43tzDEbChKDn1ByGhmM2TFIbhZDPf9LCh/bHQKwX1
nSEHL1E2Qw2q/7layXg/AJKPF81DJh9dZlDW/+lEw3OVFBbszMzi+LeWlsBv3XhK
CGUjmIR64iEtCNNioH4OvB5FrkQ0dPg3hV3efBYZf4l6DKjAQBM+na9RDqN8+GIW
GuQAA9fuBEtyUQ6SwpwEPSA29SPH8wBHmcK5lNJePf8LKu5WAec4hGQQxIt9uOfl
sfYfKHCzjFE31/yV0oeVeYTKA6+RZUBoKP+2sJVV0MJic9zSmcBrMPO2/uGjUl3w
ZBOrqtRA1vXwS5su2gFlxDYzBobluRlnvGtjGGcM7cgHOxKGolKu1LKzcphKGXBj
XUQUd33qpR1VEQhbrj35gUnhLg/2faHoL1oDvUK76Uq7KSg7+TImZduSsSGfwF/X
0VCDixisYuQWCjZZyFzjiNGCX0vA+uDhU8tWoYXEqr+sOGjxrufgB7uuVS2t/ic5
tkxinYmIUADLJ0U8RZQAZpIikh7d5gGUu/pdx/nfn361o6QhnL7iySNKdGGxA9KH
jBo8tN13s4TF4Pj6B2lOeXuSig95IIXCa2qiBRzMWZoTfu5tyylZ9ZnQFkDMKHZh
7ELF9k9TrA4vewJmTdx91/9oWbzV1RKKYiCnM0sL468hcxMWZP4IKpcU+lmc4+3j
eUNOqAJ0odFOsoZ7eMERtL0TDbmXWENLFOUOSFQuZRU7QEGDOFWkFOnApZXKtKEP
KX0tbitAHLYdHV4e2dIjLicGfcenyEQHpFDAKAAKeMj0a3ZiExm+bIihOzTPrJjo
jR7t7vITVFrA170FuxpZC/USoXeu9cqA47tI8g283uxkrFC9x8zqR7nZDurjQ4q+
WaU5K7RazW1stZptsxzR9yLLFfl3wXUanUd2kUanO638EkMYWVkWZgnpK16I4pH/
ANfjkt40C8NFoRiDvQHDybhPu32aZ5bQGoqx3cnitbtlwWkPxF8e+hJ0qsDwRgxt
q+bkbZ56IGMUFDKRhAVBHLHf1pCXYv9dc0qzAkBGoQ6LiJKQWLBmZvTQDFcqyRDv
Nj63mCfqUjgle8DBhIlx8F894nvClm+ADT5RKUf9JOnP7tdeLw4Hez2hvatqnpD6
kCCYf8d2dHjsXiiGp6KXJ0bT1GODAf3wng4fD5BgWYpjAZ0K5/FDicXggKc7zK/0
xluErrgABlVu+Qa5xd0DzEBeOnKLHJAHVzAaNfSj4oHF5d8ZeJfyHEOjQKCpgHCG
C5bjEeQluCmXMFdb5Wtwllc/U4Ichp0VUNLMGAVGjfq1eGcEap9WjOKyaBx7ipWS
EHohhOKPWmV0ok9001ypCw9eC7gFv1Rnz0HBKsuDmmBZSY8z2GIAS19Fjhzp4tSu
4k0fUWUrJro+MZdosY0sHJNyoUnOPXnh+Qe0VbeU6xW5/Vg/HK2Y86a4WKLnEMFf
7au0+GfKC8R2V2rY5uQ9YzvwiKr+f6NxeME+KzcZt8bV4xqEzKWcwnjlvtE670my
6DIIGML4HGNKXf/RIx03aXIHSFaBCw+yzeLY/E9YHiz2Lsja7hnPbB4G2ru57NvE
gjInTvgpsJjQxC2fJ5q2ioOBlY8ddj9mouIhh+zN8fzHkwNe/ob/hJ0sWr39f8cQ
/10EcJJN3+YAL8W0WnGdsxpG2QbGG3Ehq7DJxuf2aQDYQ/7gZPnTccrlPz3vxfHP
08MKmJSFmomBuBYtx27OwqXKrkag9e3kHzTWVPrdUxlq5BUzP4tien9iDwrE4OSw
U5nTH/m+sYWS51tdX/9AMQZaL9sdTagxI2deeFWdbWW2sPp8VuSRLXQXOPP+voez
hjAGiFAuOx0gDdSaE3ajwPFfEHivgxn+Vr1E4PfHuJ26GLonztK/QyCcfZyeTm/p
OiNW3LYef4UlJKZpgMxMHU4ca8Tg1p071Osh6b3kSLVF8L6Q6bDwsXbYyCo/wrTK
vvwneBwT8XeZB+nBz6lUF/v0Zl5IvcySKM9rN1u0nBFO0Uk0VyJJODGOGfYArc44
MCJmBFyAYs9pzS4mFITAPA7vcknPxysUj3+XcJgw+2b96jNu2+gIChIb0qGl3qjR
jX2wK15zcfGxShqEjwsvnuTZt1N1yIpnbE6Nq+Vu5Q0I33U3IsvaO7HFgcgX7H6V
nXVz8/uROQbkYlxE+wlGapFwxuV8PAzCAb+k+BtQl3uUdL8t2nSmVUgv5PNOWpX6
zcm6D4PSOdDjofs788h3IGILpjdvZD8zaQAuYfimDNzUaXMHdgYVLqw1DpalJkGU
ndvIeKzjgKySANVKMBVwwA6LM3oTf9pJlZvrKpu9Xcru9cU/Ucsc1EoFUXIXcEQ9
M49ZexD2DL9tS/AVzysnwZCfiMmlFrSex7zIzX6sLGDkPojlJ5PFXGLgJ6WmdGXd
wMXocWc+RkC3QH5Whe43K9H99TxzHLqENhidrIpaVnYKmQfCpH8l6+zw/eaFeeA5
VZQAHuLVe/RH6SZWT0EGsdYKPGzkuEiHQVaVGBJ4TfapAF2O9cG0dXaKyHiNe6PY
hfixPQ9BJzXmjlcQ4KvmTmUXmlBXBjP3QB6cEzeFw+zvNq3awG4HrN41WNJssUIC
GDHaiLakaKyEeYd9G+frdTLib69BXd4hRl+Hc9iUiJ6ucY9oRxmxRUKRPIvN5IEQ
1fzxRViDABIUYUhR+UM9cXQ+gw6UCTuhnEtVpSPeSHnO3orvBgDk6H7XOEaJcTq+
Mh7ec4etqKOeIwDcIZ5mtSa5P2xOwJyYXsqdXeuD0MHDbMDuhkeot/rD7PvNrmQr
CAqv0mD7zSjEZLdjW9VN9v0HTZ6R7tzsXSpE59msvQNbtG3wb2E5xelxXApoaKQy
FQ8LblkHoEAuXxYew626leX8dzm+Hupmk+QhAhEMQy+vMPR/soJ9Jvblx555sHdq
hT3YF04EtETi++cfwm8OF/ycbb4IvRfM/zNNh+thLc/BGb7RSvmXTukzSHz8BSVq
3IrRuRXtnUSg21ZpxWcqIy9iloEpmYOyN9TrWA7UeYIPNssFzg0zFBzR2iFL8Aay
QSTTgY3pMcADi/myR/6K5JN4bF00G0Rfkrxcl4ISkUM1bVgLk1lqzE3E5nPx8QFc
H1zu149Liqhs11IQjWu+qEUy42x9E5iGYiBz+pItDJPVdnnsjDhUTPmjzMiGGkUY
RzKeQ3+Uk5ECH+lnsDQrF4L6w2f2XWnKBCw5O9VeQxkwlJwWcp6mTxqppSaqORIQ
9Xj/mSELYBww+1Z8wYS6i/0c9Io32ngIWUV/9zdn3i7sV102AYJmf6EIQvZv/u44
3/4VI3v156b77Vc791m8Ajz6WRh7mExdwmPQHFi1vlvIptovmZLj416Cby6MN0yh
YQ7YxaGIYHLG2NYhKlrjamdtQw+P8hxHHHBAzJw0aJ5rQwj/hnCaEsDPG1mUu9dz
mgshYqU0sGQzJlYbTVhgNtVVDJpvt0au+cvr9vDdBLfpfJ3PMYtaz018QXUgiZi7
NAe6T7o3PZ3WE7TLiOA0tLM5wNZt3XWtV4DzNK8WedRVIko7zdtIdTPs+evUjEeF
fqLaOfFQ+BNZUcEyx2tdwlXWyWz7983qFPMX12lMBokyBS/25wqzYcDmf9AyqBbt
MyELVxBZS8XCCbbq3TanKekDsFvR5VZJmNDhp4FVMuvlgqTErNRS8EKE3ds8x7at
Mfj2cS+OMhhGceDhtWquUqx77cyFnvyckGtivyn9HQbL7orhe/pTvJ+C+cIlLcIh
glMaUCwmnBWhlMYGh7im2+1x0AWsjDPjpfrFe/geOduWPHUGdmGvvp3ZedWHK32W
l5AEix0MEOg8MRQqyC74qI3NIx9OcXWzdj3yicB0yPMYfDtlPx01Mz5ClDNaXbrV
T+mEfkzR8YLVHLqvEUpfy8AxGvdW7ieAK2tEWjCODlky7df6qCI2QrnFqKBoQpNM
DHelhajNnRShOKSOYM854VNwLxQnuMP1DR4UFpQzTrekSvjvAzSMF4/6QkBdsyLv
GXyf9Izb35S/rSlXhIi5DdiDClU70o5rqcUT8T3i02WILpJH7BJ8FOPq3v1FkzZX
UZDEDQI8Q7dViammTE0y/SZqhwBdCZtrBVsSMwNRMZ740AWn3DYUNZZc4/eny2he
Bq3yodabAleksjrqxNyvjXpgVdDAIEB081YkU/ce4aYM403h6+IcMKTdZakyfWPE
iHXu6dfIeFPh9oSNDylxBmUc632qSVSd1VS74iNjGKHLBCOoNgIMfEP+CC9dGtEM
SsQBVekGEsN4S7vJ3666IpuKpwjvNDGQovzkTFnmvzxFDSjpgDz9HTl1K/V7/f+2
VHZQ7uuyPAM9/gvyzibKITizHdl16Xr7CbrrX8m0WtRczfRBN+mJ1vWJEnzQrNtk
cyveZLqruTfQF+/BwCbmkxsYmEKb9a7Qzshlezmnh0uqBTJGFtnTeI7c2eZO6Q4d
jQgvSXzY6JPT+b9EHBlN3yETE57vk+LJI9xfbLU/5KHRM6v1TG0uV1tAFOOEeGB0
7WgLnN5yKf/9nTomNCvVsZpqAoKAyNrMDVMcl/bbakYYM2lS1kJD8FwBIrtgfA/D
1V4dgpDpltaw4Cswapw7SsqNWrMyXxVTJuP5Urb1FCMBIbopzhXWxGObjSiOrEMy
eDu5dW1UZcVO5FxTguSc3XkttsNb11uHKPxZIPlw9Nbl9PwXi/bYEU0agahQfXGr
MxHfielfUKZ6dgy2mMX/LpygJiwY1qvKJGLfPEh/gj18KIHhzWV0UeWBinMWncCF
oyU73Gq6poPzKheHC9xWUJHc66a1nuVFt6kRhBvPlHRMOj1PbDZysV58WXVDJYra
Oo0NX7tMd9zYuMTVTAAx02JoUhYFbTyEeujktzG0K6y3zTYdXWPxVQ3S0jGK4xuu
0MuP3m53U0pD+h0eeiz0hHxTU52XF5boJ3g4gj+/vYdRtRLQ3pXpy7xZPL/gWhfu
AAbidk2xFOIj9F8Du+tnxNvC1Zrz2ua+Rve78pvSbeGeU972+1EpeJYTA1e6XBYH
6HrdF2uWWKhGMVT6+E67wTe6Etle8HV7oz9yc/LdPJKsRi/zh7TXkcyhD6EzYvNy
FfhnW/Iq/q3nZe/xEKXoyU5A+KD2jX+ZmUiKBhBw/91InWmhWRpQyBX4SYsPdSNP
gnsdSrd/MKgBW/1RXEeD0FF/8kwsyBxpZ6zCdae1woURkUJltXnMkNkcFD6KAL7T
iTyiK5epIej/XOvMv/kfSSdDrTrL2jbh1hNrVdaSrqDMr/YF8sRR88N7l6GqHGdI
5SLqoTDxa3NR6P+v28K7bwpqUFPIkK7WZwIY8EXy/olbPAjOUIzVwY/GGfGdfa7y
FqxIuTzXA1vhJR0eiQDibpOergSkUszr6VQH1T6EmIDRsMk+5z+OCLTx7ib0/z5j
q3CnJzx2ZPEsKIdRbFc0cOLPK0ms9WXmQJxhDaY5V/a2p1EifMDhkv9sg3tFqtUC
MEwG9fizpwR9cqJ6yluSocrOehBw/+0uOQ7oRXRMVbYhdqEKtX+1Iui46uI4AOGL
pRTZ31ieD0pz975ao/h/nqYtRKLvWc+CsX3BI4j37fbakrWCBMjy9hsyU7bI2rnu
lLTBfAPx/U0yMqCbn3pJysn2DLH2l7xn9pfwhkI/n0Pl9/FQccaHleSitJmTpRvs
T8VHNXuvsm3Xbhtjgqq7lHo/Ud4r5PW5Rhpnw4t6+Bzu3DZRzjZw49kFFFmyybc2
nMVKszF2ELMM7Ul3HDCvgJHejHnwHvoB2K7+7AzNLA+xf6C0/Q+gVlUMyeGXXX7X
Yd4970zY7tTzA0QhNFeL1V/bo+2sak34Xt85zuj0Fj3wOs5VJeavHpt9W5OR4Xjz
JsMlivknVLdrMbwhupXHCAqb/eMlgTNfdiL9ESfhJX9CzydLELU6LPJ/YvGNMFlD
ScCeAWzFLp3Wf/TXi2PTwG5CGU/rCN8Ao+R3dK+cBk4kFzIW1Gq6S2IVCnxjk+tV
fWXUyCDWrV6dK3OzKqcnr5IpI8AWkxdi3mHPO1yoqHmXRxOBZ+gFgMZPxkH+BGMt
j3blgeBnA/5FDih+B2T5/Eh2d58o3XID+udb4g+yIHce/i3fGsz5RMoVfeNlrCNS
QyxIVFh5i08L7hBZeXLL2hy2DRCvZ5X1RcQDJlFqzcFKbfGZ9I7uENbGtAMweled
upyqnVAjDdo3Iax0sS5afJSJp7pdlTTYzPbzjnwR3e8y4Rk32hUxNWVZtwsaP0BS
TBWxYXyss168NA2FF8EIIirqEVrQeatdHZy0ketxS7hGFtnTc8kZ8goyFuWMhYHW
iVZJ7zk4oShyPL8Fj3BOX0p0fo9pmqHDHzOsEIKLaAvo3GcTXYDZLXHlfLrm43Az
HFGkac/oKKwkqiRDCobDnib9wgMgqgf4dBGhp8hafDyLISfB6hhPJaLwnPW2+6ZJ
+MOkx3qQJpGB+svjW6VExsy/kk+EeZ7Mipvc3Hqya+Po+35o1mwiZUK4KjFc5Eed
h4OBDFrT3spaWoxTdeA93idqBHgfIl3hLEqOuRCu+9FRU80fsjuHb96rPSWJkx/i
H3l7ePGiQSiS0X040OO50a7yMhx9V2oMGNwtSfS6kmUAYN4h5gsJsPHxOWzoHkuu
v4LGt0d7QiLfPuU2X2ZNp+FleGdzKfjqQbd5FxK+NMjjCQwV32Kt7YfHOC9dnjwg
VRtwSRVSbGupF78HWH/3x9NgRMxssqVQskSr+2bA11ubGvgVgbEpe/IcWYQCrcPx
bNp5eious3KkrxAEndBirWwI25+exW3lVbQg1YyR7e+pqgZmEAMuXzTFYbwmbSR5
yzTqRP3A/r0AU6nIbN2uuDr/gYTSJYvLRiaAfU1U5gj7QZVbY4zYV+V4RrkSmac/
g1bxv5UtO6hVdUBfyS7f1GRYvwh7f1i+ICQA6aHVS0UXHFOs8SxxX+Vuz6JrkwEv
Yc+ZHLJ8v1y5wS3gQTxeURsa0Jg3kyibep3CoCzqcW/ayK0DBEHpDtnV3YTjiK0P
HXTY4dDeBeDwU5RtRdni/PzTw3mc4c/+np05hG+T44HHziGiI4PBFJIrARNoFeJa
/t04IIH9W4TT3fgPsTDijA8yzw9d1Mf7IpZMe4jnTl0ipvz2TILh0nebCAL9Ct7a
SAXQ+z04SNKgj4Mgsxalh4D/eybDga58kimIIzHTG7WMsMDQwealtZtaTTl1dDvs
c8ca/s+4KwBJH5aTITc/7D+gEvJe5ThaoVblEys61ZiP6Np+RbpVzRh/oMd+/xXH
5SpdNqQyN4z26mSsAaIMLP3K8wb4fOhSWG8rEy+nWimJXlnETpWP7Y/galSRT5Or
EzOW4eFwXrAjIIgbEKW9XPEfCLtt7ppaxaxYjL8cmMhpYusOfUrAw479BYGKTbYk
w1pfAcCftdCm11UET8JoZasXWaESBTDruW3lPD38LN5GjU0C7GMmsOGo6WkzMP6M
bWmkxcYWqHSjh9wYTh0itMPmnBMIOrDZvr+EFzYCzUgqZmn1Fdec8Ugkav0Gb7cH
6+Xt1DeTuuZXNQ7wRWkzdjM92EZVR3cIqAEm1coOhUJMao7gRO0QmVXs3CLKwMBF
XVUO2dNPJhuXRpgguRD3/9YPJKQKOEDEFVuIg46OIaOfYySFIYs7bwzkM6wLk9un
D/07dP5fmKHFpw+bII5+rJZe/a5gzO8/nYbUDBOrKKAZy4BwDHyFnEkXAhB8uY+u
6PmVcuLBgc/61jnrSbOj1Nxqx/XJnA+gSes+IB3Dy6sbDslzxfdPeqYfnerrnnJg
uuoqHQsklQJ/uXy769Xa5pbN7u/QHUX8jlQ8yrcHRS+2A3Su/Ye3PZBfoMCUNH3F
J+bzhfko1244Nkth8j3Vw8bZj5aEoHKWQcjEnVRa5faBR/E9LyrvYCdSx1woBpdV
RwoqwjTdapCBbOVHTuLpR8lKP4hUU7GxuYuGBqpFIzLSNbGYD2Jy9NrSn4baLsYs
pGMChK2GmLF+XOXeArtbdHx4jUYk/NRgSkwEr49nDiOpuo1vyF90kvaL3TAkUTG/
rxuMN+MXsZQ1G/X7XUBAWYqpv+ORy6ROUFTOOTZ0wFMl8LFH+je9KCEYTuyZxGzC
+PjHtc5d44yJFeL6JkrW6+diMPOGDlVSWjpr7x6jm5K9gKRSBmsQVaGNDMZJZiQi
Px6/XWuQAmz/1artkw4vHMzSPuX8V1KufCOcAKCXgRYlXRqe3zm3XLj/rkX+Pmb5
fGTgMzkj2VtNmbHWdpnoft8lqFx10s5kMNrwWYwF6Q174uAgd9kJhU0vU0uDCsT6
vM+IP6NloZm89kn4fhV6LQ57OH5S2Je4IYDhkRtph2RiQbgWsid8Uw2iwC6Z6t0q
alFke3I6DbrvJGJYxYY5luRLPb8oOekTWYcbQKGsrQkLrHSKpbCGggPfhkAX3MHS
uMdnsC07XKzuHaQHNsIioxz24AFzThZlSqbB6rH87wdicV1ukcacg+iLGLHp6Bu7
YjsB66hUGPjXNscAAJq4bAT5uezZlvcW7iKwvpG6NKJmpbTl6CXmuF1H0OLZuK+f
ZKOM+7Wks+ajm3xYx6CVNzaHXTwOWMBx9xqWsKu/gkvoinuKZF13nxYn2NAC0T52
O6LdkYmlFfAkg8/gBNmoc6Nkvnkby7UiB1ziPMVgWuj2iZpfBQi04KcgZpm5WrTM
rNd35RQRAfoeqce89196k/RUtni0ON4hgdnEXfcjX9tvTBvvmLpCsZxNIyR0DLTS
KAYKF/wuWi4AdTcZOmN2PMtwq/CQcN7JT7hwletgaWTC+6QlfDjoTaQjhUpgVDu4
/4/aB/9oodQrWcGythwVLFQqA0tZbGzcvqxRXtGRIbd5DwXn1XK7GAjZX27quUuw
yb0lVdyu+SF7hYbQbgGzGjDWg8O844SqdZ+k+zEW0TzxoXyhCLi6RQwBFrXt2S9m
3mfM3QamWfzPPxvW4jNaOR/jKCfbpjCeNfNJSEv94OJNLj7Y9oRxF53n5iZDbPgW
036K2ttiys5bKl5hqmJfieBmkyOAKDEw8Qs++XTgTr+/qn1smGec4vHGEu/++s5E
8fCkZrREiioW4+7W3PkcFs03zymnrqL9JicSe0c2E+MMRe5yOklGPAOyWbhkV42g
OuOxmCcqDjrYiWVAKv5od9CayTe4MWS4dKO4l/4fJsYxOayTkBBTgaCDA5iYvIZx
rUTdvcGnN/zbKbmozYWFs7yHIHI9xfXNNIEVVa8ZIhLzKJ7Pfzl5xmBMBYry6rxz
Zr784YwZDSo9VWsjVtiVJdjXRa1lOKfREx+XcwwRnGCVbpJ0c1gbumw5Nuw9TgmG
gQKKlfch5gaplr1ByahkuRsCRhEZzUqSXXuayk4VosvOeeJEVVjQlZdc81kgAho4
5rhlnLnSbDakrdgigcJJwHM7kljLbiwaG7+NrBbEvp0JURBhZ25H1jd5eyzohN5r
DAKMxi6ESYzYvlhNvCZi4bW4VU7K28gmBxqmZT1c0Yj27MagiatLBQyYoG7iB2/O
CZoMXccYaJBokwvwmIVwJDK38ZXVqhneZOs2X9TskBz1omj4LrV8EVcuhANDlgZ7
HmQndy/v6b6XOL9fP7X2KsYakp7CoWcLTmakZ6VhEgH8mltmmbgz68fgn9xmMs1S
28kdE0n+ta65teo+gMhdPUKBKYE5d9lRBfVoEJbXTrx6ayHifLLopwrgW3aTDGW1
WVX+qIeOAC1tBoOjLB0RibHaAyuHiqgHo81YdkkfWiIfSXSpsezibR5+a7PmZ87i
Dy2rcTLObp8jSYkjuhw0vsYOF9tyefqS3Ih0r3PajMu11SrGKvREI8Czl3gHed0S
20TFUJUfsZg2i8bu6lxqz5yamLFbnYGjmRZMeX79QqQk1B63DFd5xkba/BuXL9B2
i7XjgIfakNNkszbyHs7N8QTFuWixoTtcnkEuWWuYPTZnpYMm8Hdm0vOSjcBphYaI
/V0UnV775OXGK8N9VqX4UU2MDCO+I0elCp5s5/dCpa1KsZ0opWsfQbHvcBrxbLt7
j3bUf5kB9hI2ILz2AEbQ7mTQ+FZP5V9GxjOvaKt8F5bXHK4tsDysGr1HCub0Xqg2
Pj8dExW9mHXrEAr9MeohJtUUzbBvLYxzkamIPB0Vf3f+lQrdHfhLY2B5DeF1UZT7
SoIBhy00znixpT6wkTa6owGLU93srS/K0vPZEsPUzmw+vrS1HgMsNBT4x5sbQbsm
3lx8NyaxeU6N/KNWuicMt3NEYl4z4pFonlRrauyn36nPpDk7xzJNRU7yqftEjJDJ
/YVbwnGjQPOHT0Iz62MyH/KoV9085yWZyi3WFPbqdKIgR/SJsA/8lMLcoX6tRBj9
gBJUOf7HcBKoWu6/NQW2gk1+tuel/CiysqGCC+uhwOICwBPrqTl1NmXBQhM/d9ZO
FRl5QamCzBDCfnkLhLQ9BXi/V5ckHcCas4bD5dDpO+oIUZltsquAv8xzTyUrTGWe
WphIa4NPVsLl+HlGft0mRXZclvPvozxlXHruw6A46n97Zd5UlTKEphYZRXflVyf5
z2V8xHMzQ7eq8/KUee6PMm7FyH4GNR4MlWNSOovv/VU7VLQx4cAfFJJ09IkFsjP9
K98pByLNwO9BhYQ/KMNkjX3o8BdkZECHpbf3Q3YKloMj/jz+0mixye+sU/L//YW8
amFvJx9zWpKClmyehErmTakUDNBghBpXmpvG24djyWlryeBNuR54ebJtV6BJSIfV
tKbLOJvVa6W/RBdlyicOEcekhpaQ1Ec4PXePWmpS58kVcaanax7XBB5L9iTOdalR
Nfg4/THgFyGLD/nVXKHmTCxYcOPw4vLS4RnIOI6JvFc8MclAG5OTQuTgNW23+0Oa
cezH8wjzPC+Y0MvARu2Hv4VJle7gQ7g6VcVxFEtrI++CuKMSXEWr1QcTYP952hBf
kPmG/SyndDmU/I9OtyCf6/HA2sG4pxlhLmQ+uZSU1K6UqVlR5EIT0TdXybL+1CHY
NVEslXxq34YnQ18+CS/GpJ6Q2gZijZFSr4wpHOji0njWMkTrHJ49Ap2t2LCYEtTv
CNxJw0VeE5Aam/YYubfFIF5BcWeO+WZfwKzh3j1t0zomys6o7e1b0q5c9A6CLof9
/FfElKbybG4q2LIIyaBUjQh3I+qKOtklZDXJ+vlBVQnsvnlYtRlmq8RuxncbDTJB
V17QkIsBCDnNvk7HEMpDCT3wWsfAnmMlTofQuvNl8lp8xEDR3j8sEfMIfxQ0Qw7C
taYxd96sSymnf078lbFSoByl1VFr72xUIA3rTXWz0dDh/oe/QtQdc0ZmZhG4VKhL
oC4AwqDFWubs4Fu0LiZ6a2LpX+9tmNamAz6Yfs0ngA6dC0juqeWDP2t6mVv2MZsN
z3R1GHTI35gxyXO4tMJ72DSgcmtl8l0oa913aDb9IlQIg8dL9uA6eFbXVsnR0Hfk
ozYLTkPoXLRJzyOfjeSMjFvN54Vlp+8bKNqmt0IxZRvJ81xrcHn1EuIpq/mrM/ob
hYkENsmjJbRc34BGzRo2hL5Qj1uT3CHXzwfBWHXr2AKNtoJzhOEubH7bUL9P9ENi
seObMh8eJxWJDQMO5BFoxtv2u39QdEyLNBU2kBdOO/GzCLjdWRfLQTlOmK1Gnbw2
53eYWdogiFSKij1cxU68zlIq4uZ339KD/soXHuWr5to4Ze2dfg/ldZxsvmDAesvS
4FXp4YY0GZxTBIZvAme8D47VkAAk7ClWtNFnl+nwzqYCr7/iGGph9fcZcluCUqtn
H4zXbxyGSjArrlvU2xItdYxbGGhO6RTAfzBBJsZEXT6nrvxMRx5rL+DtZ8V+akzg
SxBmu/8DFGeMbkARGJ0lG6eZG4DbpkbShj708vZwGMBimYnO4RLfID6Txj4V7jUz
kvyMu5WD1jRt3OgZXyChkMW2KRu4wHi8f0iJiTyuciQIcr/8g9y35HCGzpfAAcVp
LlUEDlP4zFUDTsLdfrhVktG1aoI7SeYqMpZafS2S8LOOoJwnO+Cev5R+RLwuP/ep
ow/bPk3CXUi65QvIERf47p44KlEfclwNUllklWvf7pAYT/tkVTJ7s+HILMTH0Eb7
uIfs4W9S3MRsZyYTzrZm3v9uUKV66irePyxXuvsWpZCGfLL6d4DDKEKhcqidVcPt
BGpnZyWjBza52mvtYimrp8VLCMe5KbBs439TexCQpcAw3vQ1SW+4o8DcHFhXUS55
qI6DAAmBNgGFZ/zm941PyFgH+pVtarj1m9pD7zUp4vP7Df/oxI7Rb+h/4iln3JX/
g2Yi2WWx74gH9PGxHugI+cdqrwk74apFwGC9M9BrY0Pa9N5ze8kMcDiBfDkyejY/
1KhS/c0XpgUu7b+Bh9CR9BPugqEqugy5etL3zLMFR+8CF49zLaCIUddVe8NobdQp
xxgYo5+nNzzXjMMo8xrEandG+uNtp+dc1Nrd8T4LV8yrGZQ5B+IuGFSli4N+Oc28
3ZXrwr18VjUPaCvIz+UI2f+oM+eKptOMleoOoZ9UBt6+s1rwnPy57UroNI+uA9ox
pq9gPQFc7y4x6xSJ9SEWscM/TCQor1MZn1+kdWPpkTc35MwFYbXdbwOl4AZ34LMg
cUICTp64ROO5EiIkMuCC5dbqbMsN8O3TYCJKN73oPWiQtOwlGYgKrPG/cDk6+yOx
O6qzpCY+RSQrulkUweE/g4g2xq/zSVqHUnLYbCnkg3E6ILhpibfVC8S3UPwJ4rUJ
Rus39E6JSsLSKHxsz/ZSK7iEQZ/ggIZaJDKLl/fEHQ38W3hb1l4rBQiTabGJHc46
MmhmrrlDbZHBgxSCUzbCWX81RJRd++tyR9GjRfn3GZRJ64Q3UlBmyHdlfTFamqsl
5liakNNOBLhaeKCEo5yA6tiAkZLNvDTBoMmyLkXJdaKVGkbJnsxesn/fO/oeCvZM
kA5eKVrp1jmMWl5N0+OVKLyU+QEE7Jj4VBbtoGhS2iulHIN7QVQRA0f1Zuh3E54W
m1/ayHGw0L4Du49idJv6lUIS8gPaQm8KyIzQ0BoyfmAIPkDZNYkqnMlFcmDC6ruL
nVxJE+T5QEOPWBuUQE+DP4LbHIMuCFxokoseNeEDmq2R37BN7FlQh020rQ9WgpOQ
GEGNRjslTtHFh59/HVu9MxSeeQnYfpPpXOXltQGzoU0IiUDNUVEht2A9Pu9woD5d
AasuILOr5galA7JyRP/j98MRyuTuKsu2Gu3rRlCz9LwaU6uoBCrA5RKHqHzdGf6+
Kj8BEiggQxZOvtED7izolsIrzQj4cW5SOpEzq9+EVbEMK3j/c5GnEkuY9cliFFYu
iAkdI+DPPrlooGQSuKryO28HHk9iWsMZjJXmYHucWDzgxs0sehwytR8rbFqaTU27
QU+5zeYVOxIv9FvR8CyeUjRXhJW3qMbagvL7dzN0tO6empR/ZPoOveBu3ShfspD3
JMgaZV8V8bYORzDCxi+T9jyXfL+95RRLKgsBiAfRc6o8Sivee9mESHJ3fhc1txl0
t02oAVIeMmSM6ce0/e6FCv4aUUPknn8t3BanVYB3Oqrob1QgDG9FrSCwVbNIwauI
8233CjaEIKd8gea1V1vtLV0zinbC/jH+CSAWTKJXZ8KF25e4ElxR39O+r6psMko6
YQynKWgJsUk8QFAAfesLh5HfOY8EyJ6cIaVs6O142vl7LGH0rIUgrF7Kb5hZaoO3
zrbIICMo5IyBJwQwmU2TFxtjSrHRZ56uLAEYQj/4RAVeC/2dWIutdoBgl8fjB1ZE
2qitQnjKAlKfdoeQ4ix3eL/YptvifY04smZrolqnM+I2RsMwTRlin/8UPQcuMdsc
4IInCBoGF/+h3ZM2UV6ObDShdTcwSfgWKbuudjy5pRO6VO0WQ4BSVuYCpyTFz11V
G2zfqPr4xQTgA6ANfA8yoMWemQiFEz5jd9hocdnATN7ku10UCao1jGokcAboFvzj
PS+YXz+toxA4tXBFk7f+LJEmmX5kqnLFFVvECGCs56Ez7IVl8FqpNimT5azyWcqr
7N1l6v6k/WqLvAo4G5ZOlhOG9yeQCLoHsN+2LZKNSESX6h8Edmj1m6D4W+NLT0nH
HAxEV1uB2cpd9Xk7KF2PZ82mwrQqVIey+pMeC4frYisUqQiIbrRfp4Q7mGiYXKZG
w5K2SEw6/Lsc4BGHO1fwrcOjp6ulywzPAP8J3bMMybNBPLir0UDSzD26AuKF3WAn
eUVodIqeo+AkKOm1vg4DG7F/2FL7Kpk/kQF10G91av3lKB4kCwFWU//Xn1RRuawQ
8ACYxgL8Zl/Ce1rvoIaoIOQ+IpdUzPZDyL8k1NNLulplEr0sCRsSf5BATIuJWY7O
zYH/KLqJbG4bnAq6aqptgV58/QJvahmMm0BMkMD23v2PP2fNSsLAltHslza/Ri2Z
RNCa+tpON1bsLzyaBvH2GCR82ao5YeVASHpKh/7HVoBRFjHJ1vNHwmznCDDyvHF6
Wsl+SvHLOBL0d+3t0xAE0lehuglEqPSBn4Ptjg74KhvLzrkcBRYnIr9/7VYJPpJe
7o9h2VCg8kR8c6BV8OZHmt7qqEuaYdAv+MQtVToSm4qXHMspSF2K1ym7HFkN26Nj
U2F6dS5H5EgTfWSUmim5sNh72oTJOovQSOUnyF+NyLcQ1dXO5hhXHIno9fSmUk32
pOgrCXFmci27MUHKmTWDLItxpzdxhqSXFuqJcX/TCluO37hKWdtOEBq/uuL1HzE8
PyugFDLmBPEo1/dkj+gfAjEaAlf6uJOqznoecDWFDxa6mBLL56oms9y9u4gWjPyZ
+gtTlnm0z8i6fxdGqXBRH60wM8nXEXdMDKBFtYVPRnfsjvAm/x/qi09rd6teAHHs
c7PgtMLB+TT0CgJGBN7vlBPF289Bmfy8yZWMQRdywEK1gRwmeaxJt9DBopu3QZGm
xQiW81x6yxbgzZeYvJbFn15iycIni2colqcJLPghjgP85qCfB30r247UlbH0RNa2
OGuyC/M/kOPikgGgM5wSGhxvLe9WVcyGQtJ0+1+GpSFjgk5IvwNTpDjF7L8avIVK
2hRpACMv0kP5irndgOpGLlEgANNJJpflcxDFhrX2T+2UATX2CFazTDUGnH+xNa9q
eS/VFwUb9dAYyQ2nbaTWq8wLHO/973tyXr18YMF3ggrYANfFol2OIBJZCc95pypr
23+tXYIV9GNHtYhGthIHeTrBnyKzHBA2OMf32JPdQM+0f3JykaDMaX7lABbfPiFk
KmvWFIoV+/z4szAdTdY6PeMKRKB8GWK2NI7UkDl32JY14RdvR1+n9v3DPvvSbRWz
uVfznKM7HSEsAFP+4my7h9I+MX4My657DPoZXUDXjFQSc4vQFFcRjnYIL0djfAUp
SpEpAZdFKiFD/H0ZxZ+sfIuwwinA3aWMpJrAqeB4MONFXhjVqYmxcQ6xD+XigCtc
BhuRLniLnV5uEiAQeW8CgwFimedVXyyvxx04XszuPyhIu9jD5XRV3jjFYF0S/key
lyyxKcDLQb8Zn/zJGyxuQBHgS4fBhNnfVu4ssUVUr4LWlxuX/cHpiD1eXAXf8E4c
rNwfcG7U0P0cIYxQj44VRAbxyM3bgyMiG5HKFE0g7sk9M8ja3YdNNlA2MUos9VKM
O+TJ00XhmFFO63nTGBj8rcAqKygjFihDuYkI0AN1oO4Pb2c2yjtWfwAUOxKVPxSV
ZvaGpMqFjUrXL5ycRH/Nc3RiRu7hWGiXL37nl30omxOM5vJdJZaUE8I07Dp+FZaW
3b2+BTy18g9SZc/e8qOmViobIiC6xjaDrDnKdG/YMd8v3zGUhRM4aN06neoumAmg
kbkY9FOM/4ynGYqRlB0VSAcIDfAMtHcEtLI/oJ6zgV8iT/S9GOEdtp9jv9W4v6r4
x8HP7OmpX4xc3sR+gGuKyzGFFBVnSkAJb0Er894uUhnjAhrkWOVY0FNiMAfTmkLI
CT5wwuehzq/gjgtFw0NGZtYG3ZSvFwtFMAYRHBPTWQ1e4ifyGtCKs3RH3LNGb9pf
5jnJXx4F9AF++ZXsyIuPDnqiW6ZT0/OwrDz0+xjVQUIHOubsUtCGPWxey1PrKb+B
VY0TVYapc1sKvRJEb2T4kob1w7gQM69ZNZWDx57OtqnNyatNae/cQwmIwo0uDYCy
Gx+ZN+at6Ak/nZhTIL4+bm16e0N1QuMH0CNDOhDuLMLxx8Ds/XA2qTjaD7YkDlDy
Plj6cw1YFu+BAMRjsFIJX/bOBdZt1915JpubfHLrMJoRRgBBgdoeePWqc+GjEa+X
y3dYDxdxh0Ucx4my0jqVJSu/pfHNZIXd3k47daFCEGDdjMCyNUsy9HWgPRo8esIP
EfeMQSrOq7S+L8mZ9YT2zWG0ZGIx1ux92Bm7bVtDRYmdOtkKAtpv0qGECuCFBam0
KGCGMOCmbIguP/HgVDe1HTm5sjwMoo1UOCNCvquM73MvdnKg/DLdNjrNkT+lVnpM
MAydVel0OsPFFfYiW6DUFipc22krFWK9/AiuvtXmT5vMVEemtXYJjpo7QXOGKGo0
9QqVbY3QoEz+AxPzcEKtGIhretpnUrb2cwW8cB92fAhC2VkCcWGXuTg+O0bNjdAN
TqFeprZSmUvG8baKbuBR9hw7f/RhJtSwelEgXwFS0UeEzV38mxANyUQPDKn330Bx
BbuyMM6+5w9zOPw2/L/n2+D5XO0EX+D3I5DjQqhTVg0GLc4l/RhS6sLBuuRqyYA5
6ONkK3j1aVYrNIEYBEUgShEPADrc/pJyiMHr4swm05iKpmpKnQJH0+75IL+fPDU7
3VV8PEykYs/pdl7A69UKkIYf/zekIu1nB2XD3w/uWVavKku3jPcd+R7N1jGFgqjJ
Xl0EKc6yShJtDBYVI2ybGt9aEw7I8gkfs0b8MpXSNERZWJj7D6Rryr7sC9J66IrI
s8uiMrcQr8YhcgoCjgbzerHW6NhUXCne/5tMzv9YBxq+reB5qmWjtvERqrt0VbR5
W6U/ujtnl3meFxWoo33ik1H3xjwNEHefNVGQxEEuD+pARfdfLPSMF6AkZFXE2Ftd
vBa/FLTqmtyNz1Xz8KPny7aY3kXdIJQXMfr3sKvA9ICAK/9+L1ecvIUCG6kyyq/t
iwLpaZGSvh+olR1VBUkcI6dtFRIgoOPqVqe8G4zt7eayQjLgXDS5KPgKAsWEXBqs
W9Fu/fr1j0vrpU38/elNablFs2tIEKyvAvjUQc6T2kTVNEaF6UqbR3gt6xCVxv34
WRCrTbAiuP7zEgOSEO8UfRXi53xlR8luklq9s2rHCCxfbYQK0MmA1SJS6cOgtNQ9
Bx2WKvpwWO7zQKLAMD1n+cnAtsg+ioyWyfrSmOYjSq+mniZB45SVp2UM8DZoQ8ca
zD2/BpDnJ7aUfSQIQAlmHgPNaN0zUEvUrF7xx/vSJx+Ri7LjiwdMUjGWEbz7vCse
JOQiQfMawlMcp2ZmOFl5tYfZw3juPaFwwSihMRXNP/SW3SxWUIQszYqvNvXCyfKY
FhYJfqkuUWrqO7nEbGNdZYLts9WLyG4nlt7n3LppLW8aWXWXAU3BxxGI/K3x6LoV
GvgUq/mywGKYCcbXCU4GoXeaim2Suc7KhtkVgbycICXfRDwA6juXOCRa5FdGt6zB
8u2l4CVLlciz+ro8yp3K7YyBGp6c6ue7hozbO/1aAtwzp9Nw5QKc4PjJYSp3TbV1
NW7r6gg275w2B8iz2OeGjc6/+bjn75Sih8Bl6k6eou6ftYAv3Vv+cJVlTT0BwUjU
9wTq7VLit+/xB+5bsyS3BxvLjKik28fV+PeY9j4C1bv2059Uwj2MCo+o8NfbU0+I
VokSulQLFTnvI+9Hd3gy5Dv76QxD5sCsTSwKJVIlXXNxYNz6nvAcizC+xYpj1ufX
PfrHWw9Wrrgc8mVP2NEWg+H/rzr1nVXdogkMy7vVbiZS5rswj3UyJBG6yHB64D8C
7BKk7o7VIeHolGbHUvntgqan2iVl1LUNFywXCQLXtpeJC1Yz1AC0hxyl+w4Vhrou
qAoQPSl7eVCLNgBHW2/9VPDDLM8FnCSxKvSDgWL4CdIiTZ5kpSpi5Ftfp59+3T8t
2wRtSEdBUobKv7vNXdrHsazSR4b9OSpGizk5XWycZ2zl38loaw2oXUhVehI2kayv
ABpz2x0xWjNUGAv9R0QYA/fAm3C3zqv5XlfO8anM5/gaFMpxTotW8zf3yFH70ndF
qn+3XVb+ntVLqBOjaV+q1Rym20eBscYnVeL3squaUfLWlccburkDswyndmyXuth1
euRw7Cy9zV5NsPXi0JLat5EOu6qXmSU1Yn9cZtJapctuPFuaJ9WvgrkG6SjqFRAf
iuOtzrm15hfAzphwTPBhFibPMGaa7vSk2dc+iQHqJZ+flIjmxye/46zmYx/7Mtwq
XR0en5fQs3XUBVWKLHraFYrO0o9PgENyMnPmU2pqk6MbCMwE7k7DGPXBASoLjBd3
2C0s4YaRssHiUCenpk3YLGtmeOzWwSFVvL5nQxWU2FYCeeBp49AcjSdVFHGFuJFG
B6/v5nhUgCQwJi3eHx6M9bckkETEgttmjXVpkVY2+KtDbXiF143gs3Hls3Loue+Q
UFOEJLVfn7jNGQfywXtdiRsuuvI9/qjCFGZCbnVsvjc77ZcXev/lTSRdqxWPl9XK
0GzRyEqp8289A8szxIzgvaUe+3bQhLlpi+GshGvptF11AmoETK9xphZSAVu04G1G
7JiyATGaarmsXqxDspn26hcWj8B4pFf8LjI4zfyWk8H8ABhKgwGquLtPXXQ1LpVo
dXqska3VaNcujjGn13hgMfREJTPi+5rM+xfTh5ii0IwgFpUumpacFEHWG7qNB5lj
386FZt88scicIHRrP2O/rQDuSf7pekfFHogbs//i9LVyoXjaKIQGv6Lh/PtmB37x
NvFSogq15+vfvNK16MG9LWGcLy5LIf4vCiSJnm48GVoaAq+g46CByOxeVsq8ligW
CTmeMa6jY+2ErJyg9DwHmH82C+Rhte31PwRUnr9jS4lhIFcY9kLs+nIu215xvgXN
E5JFwmmJ4AHbwEzwdWdWeRy4LNGEkQDQVUY+4fZ4Cnx/nLudHrxPJJJq6JFHKINz
B5dq9vpE6m/cSMhZ3MlWy/TyXOAfmxVZA4tyfUYAOnxGMWCdYZrCEiU1FdqE81UT
/uhZF+zqZq7TDtBQe5L1j2FuKKZz0HspYGTaoiqAm2AsC+5YBGv4XAQAy/G3ZN+i
VQDhMSVSxsGKV6Ngz7s6hr+NvzV7Z1Y5Qqrb05pjzVVHYfxNPxGo18L2brnNfrvm
nrUK9IPsu9BuQvRSxNiPueQZ+kqJBh2zJh4EJX4LLNKH0LEabbS2I+KCukgjK8Ax
lMsoJMErKmNjDkF7l2C9C6Zgy+hdEWMnpqq38ZmsyHhadElDXXMTz5dXZ/YEr8nm
GXm8FoMawHWcuZH270AspVqZcA2q5XOlZEGeOp0VqG/b1VWRfy0f74nTv3pxv1QR
Mi2i9adsKYlAeUFssPrBe1vjxwcwYkR/f9zpchlakW4JOWYQhs5cZ9M8LI+fiiHh
N9U9iu1qDzkCiiKZy3bmRbcBcKO+eWKtFBhmM3B/ZdElWMHcxSXLmZ+TcLehF/6f
hrpdwEuG9BMCCBWGPh8ghn4KD+BDhIf+0nv1lma6WjE1rDtPZqQbw8jzRucaf4Y1
Rihu2A4wFnY4oLVq5D0tTGGw4G67C9i4bcyo+nBSDOQvIYs170X5qSV6TDV0uBvJ
ZwDdH/N7nspEeKlN+IBtu9Y9LwOmQ7/nzy+yjB93Oa9+HmGgmtouXr7SsfBLRE4g
iGdKMEqEHnr3bwF2Xn3W9WzFtlAGEeq/GiS1pEDlWVpxJKa3PsgYNlg4b2E8tYbC
a20ljzA0qP+W0ewp0/IJLorXlsN+GrebqK9oy37z8PtlJfpq1VfIlZnjRbF4GSbS
wy5AacaXzE6aTMDaxu9NqmkD/gcBBuk1UI+s5ff4qnkJAn8AGwpuiHKW7dzpcLcx
DxiDo8k3dURz10fAAQb4nFu6l81T54ywjjCAZYOWTKqS/XPVpRpMp+3Dn5snKpFt
wFgLmamRVPCb8PwgoGlqLakx4T0zBH4nj+cah0/A7L1S4vKT3eB0ymM904y39wW0
J8tgDtZnomoew8vFktkOgeMBsrxZqcgq5rO2fWXlFwjqKdVjZQuij4JbZr3zBJY8
299xoGPtMjwbsCKaIswcKnjHwBKpaJB1j2ZdL851XgKf8K0mYrHI5HFdpJ8+kyHU
cmyPJ9SMHU5Qh8k1lHyhKf4qKbFRpF4PKEj119fZ2aCD+jSe3jHW05J/n0gLskfb
axzFQ9G3erp94Chtwp60iLRmsMBfLTlcT8rTYpbWa7ld6I9sJ+23H/OmJHl8ukNX
qx7FI3ntHiIgdj4lRRlaDOIpnDbpFpf6X+QkksZH/8mU5lwSFGi43o4WcjDr2mAb
3kQ8ct6v28RmWEpQGeXc4rsMspP74IaepDNeG2KPkt6vWwd2kpOy0dZHB6rWy9Sv
eXVNtu7irjfHk+Jsa0S5B0Ipc+YLBVDHt7qbxip01aQWofU1uZYMlg/by63pPoMH
uoogYc1bPF5qtT4E9K7OWO8VIZ4sDUOsznGqHddi2Fdu3Mn5hWatOn7G/kBX4a+P
oc2Vm9qlKDo5wY2UGcE5g5ZlEXxbamTXz+p4dMhcMeGB+OZLa06k0vtsWPpJ2e9Q
3hNSJwq/+HvtTOtQ4ZfINnDZxZcddHz1i2xTKZIP0wZ9fVNYR5vWg056G4Nxn+Jg
To0jOToAqXsPiYOJoNo9oLyYotTBCZrZBeTDsqhFY3hgUoLV8hjcHliHC4R+9bCU
/qJ4+ksiAZOa4tT6oU9JKAkX+5NxYN44O3WnhXX8ssEICz2biyszZlRn2YhXa01B
i48KMGXVwfbCc5ISO6qfUTsx1BgexDSCYBHXsEVdpNNJT8lMsQ30K+Wpg2taONYs
RgGZTymxO6hAN6piL4nOqyDbx7hd4G2R7465nZr0sng5wsuqOwzt850JTPgGLz9K
vfTFvzafoHiIiIc71BRrZYwbTzYG4hBW5vjekMEYakCDQHP04pydZTKjx54fPegn
deWFuZek4WMl3RIRfey3pUQx29XOUiYKxbl+N/jnxJXGKvicdgxAOV/s+1A6ICsP
GYo8DDXoJ16tW0qt1UAneJfjzri1j+k7IOG6DFtKN90/HfxMnWnCLrima/IzVYUb
aP+Lt9nxaDU8wkXY50ppsasfyTT9zw/D2WxczOoxRXSLmqz/v+WZ6r36t87AoiDt
49En2IGSja6DK4AocbwEi/ktq9HU05WUkb44fRo+wuLNgE0qSXiG7t5avud/pb5M
TA7px/FLt3kE0+iXQVz7rknHALLzFZ3sflz457yk2TYkKpv/Ui7EcHZV68vzVYT2
TfiXqVfTd2lGIbqRDjCEmXpoUSrbNt7psOp80fGO/+kc24AI1t8m8IYG9ziwr7gc
80WXYy1R3I90q2grdZ4SSDMtrAZ3gr7rbqvr57p6wFiXvcaFQXGfkrz4iLQHcp4y
xh6DmsXB+T1H0Fo990jyhesmqKzBGVxWRAR5MZanManHx9Ppbec04/dZPa950w1o
/tGkUmILhKooKO4+Vc+WRe+nPLeX4CtFa7lC8eE6wrBkfBkoySjSvciEJKsZzaef
6ztcOmSxIjF07sigFYZgd7BdlSorligHHyVRSrHzvrnosvuZLo4r5r6OCtTx96VQ
aL9UlgdaXY5hki4riO/95T6c9pvvwqMaX4NBpeir/He51i/FIJ4RCEKThHLP/yQn
MHu9+zmfE9XrIyMkG3W4XrHmjjC9iBfU3QfocfoTu3MRLzpSoW355COeIFpTb4Su
MPOvoEcZrF0aL8NiE8dGfgP6fGTuFMhi4IIBwd82yOY92dNH69CXA7sxfarNVBgx
yF+lUMcCpHFZdQok36TbXGdrfp3aJkryfaTi1alfaZdHTH0LpRQwNWNW1Tz4fs6Z
sHo0PGkjrVY98Ebt1iKJmEnU7Nxjcr95AeBddyGbjRiNkudatZd28SN4hqQIQbqA
eVUVNTSCyCKMffw1WLOoqgIKppQEKzJldL1azt9fftO0t4L2Iw8sOtszwwoE+7fE
9S4tzA/PeX87AIDQWeVPJxdg3Ldl41HbWEg//pym75kjC1lvAuLYwT1njm5wtkvl
vrFRl+TOYlnmqaFiqEw5VMr8U15LqMlwgc1veG+2caYXvFMD2T8n0/zCmsJw/XdT
cxkGGFgsXqqeEJ7DxM2RXEDGzCdbwZf7M4g+eChIrAqqJbJHyRFKiz4mkFqoPnDV
GWbAwioCdWLXhnJmz3ZaNaMCDpAcIWECYDfXpiAhB72L0uPNTLU+tcxugxmfMbtV
vAeCeGGsb/EppABwVDutVmSLsyc+Yk9rJ2jRY2CONfTSL02415J5KN7uESAQsdfR
Xukpr1xz58yWM0ag2quBuTl1Sd23lLc4kSO+m/CQK1Rn898psHXLnvdv0bN/B9h8
GMfFRIQInhe4bPFoSvtM0YuTsjBkk2ugC0QvZiZ7o/ictH9QS/hZCOJek7esovns
27AQNsf1RHiEGSmk52dXWbVWQuao+eZ63FtiSQhEeCXmifBrqwxeitMrsOF6Obs8
i8/AfH8QllD6XopUpdW5YH/qqv1KIoki7SY2aG+LcQVx7zeceuOhmkvEZV0loTbK
VTNRne73KtC567v85rtRC9AkPIz07pbnubPClXClfwsUNt0AVJMfUm9K1e3wwQyd
Rs48e+B92f6bxwAyfVKW7wLGjq+ZY49jJtiZf3ukWs68sBIm7pHBBQMwohDWsE6I
a+Qxdy/IO3+zb/MacoA/aalNVGuy6hMpZKhzXuaTyChN6cVlWqo34LEuL7ijRZ+l
W+Ku985aDkBkV0pnlnXjaw7gY7Za3pAQ7u5/9KTJH5MG0KFW1rnNogwYQxl281MD
3mV1GGpFwbYHT4KfgvneOfhgRkhv6cnlDzg4jSaFRry5qfdMRGM8auRJB1WqQQCp
E7pygOPSpmGgOS9L1hpfS7LxeVy1sFNXF6nqnC+6xTsuHnjfd5b43ZOPcGc6G6r7
OlrZ8Kh6Iv/ZAL3JcF1P27JxCzKt3tWjWwZqAUT6a0gxgfxnLg37VAcoOnowNsCO
mbttiemkodkpRkS7hk1p/j+LJLQWvckxBLaTyY6LbkOtPsAAhFBsKhhVDjFJiIbi
Ps5DeSP6B35bKnKVxXNpqeU2wu3+EeqZQRxe0OmE4MLDN8N08IOjamBWdVEFXwJ9
VHwwlagybrfbDwvaqp+h9PqhzYCBwJkZUj+O7abn49gqNxdY5+TBHCB27VzRFnxs
eaQm8r2W95tbHFjv798UtSa2b6rviy5vTd+CZ6FoNkud5od5l7xwVo5UCbXHF/Y8
iFw4iXWSOnPWKj/SRDbPiB6Nhvvm2EvxxQWuQ9D6y8E5TJN4AYt0UTr6AhziYJja
EsBvqFQ7XNTXqnVTIgLc5F2tnrBwsELniWQ1O4ktW+iqIHpPTcwS9/5m3jp2EqmW
KbzvNYheqPNtej4NNNY3SmGlmxKBvyMhwsZUdiOz+WoZXT+A6lJz6o6evnxGat0F
CumLGK7i+AWLqnY1bn6tkyATk2rVRLuRO7H1UcxUeeMmYv5eK/Pjy7dw4ADcKtVE
lX19eJ57IGPd95xY3WV4pvQU+4HYme/bXkCiOY9Thbms7pZKOLw0f0Ep9dHhvDWF
tp5A7/sQ/9uyq/L1BPz/LGfHkAIcp7NOVFiboB1Ht90gfUmPV3o6zDZa1Dpm0uSm
wZrpUu2ZJUz7Z6uDdTSV3Da6hrjBaEnoQgvyh75DH+89M6agGsotUDyG977lf5cS
CZr1TFoHTgDqMoS8Tm/M4lu968TbE5VJU/8riqe1FK4qLaesNGU0jGQWTbXgbL5e
WD0KxYHfl/z4JMAdhtdBggY44lNUaMlZCJZrQwcPmryQNjvJU8//XCNIsEIqXw7Z
scYw2+3zhdEFJZ/owwdAydCGPIDx/0/iKS2+tly8CWYT73fVIzxx91TFONKX3T+/
clRyT37EfwgvAyAO+E1LboGEfnyH7EbrKVrStSHDrwLvQXL/a2KiNpQd4iEhlNWK
ZaKAFXqbzGHwYx3hq7ZjaQDWJWU421q4LRrMtHcFy4/Fw8PQJ/GVsKtsabpn/gha
o/h0ZEYVGNH+YTVm74IdU7fQDHQ8eE8jMRNnNuUpYEGpbshXq/umdXM0uZT2ITKs
0gMM3BuPoxy/RBYeDhYrQY1juH7T0aZVtZLt7lfPCoQLauetaEUDFEkS1vFh3DBM
jT4t9EpnOFQxpLhDUrl8+sQPvxPb2ruhjDdFZoOX4xKuUNaED82SAK/KMKYQretX
PbIiu3y/Sycr1zbkEBJTeT5vLa/9g/ipNhLuEdG0ZyjHRufu8XHaqbFza58pZH3U
E7PkA2Twap1Tc2WZhZ57mHQnA/Eijfxy4K4uDIr9Has9zmjNQv48jfjouloX/26J
kTtoU31Kwme6GhcWqPKdoNcD4PofiRGH3YqyYmy64SRywCx8mTFuUS8sjrzD+V2B
76KGFasKcgXUvCvNfTycPoPiwZZQFE4FEdzcgsYLqF0L/Ft1SC99oWrF8sxhHPNa
wKldhRNdU4oSUei+G0k6oCB2qyK4DKA64uIjvT4cIYkQc+N+n6A7fWADHqzvRIjs
Ow0Xw4/7RCDQUyY7qGI7nIzbFVIqBtmX8NlgBBBpeS7Ugf2yccaoqkPGbNxpsE7b
b7AGLcSN/2Y8lHWP+WJN77gNYF5aq+4u0RVLsm7WZDmIU4TjfcagNSOkXOy7CMaw
RG8t+sbRkd4h/ar5Dv/cUqiZao6jFDyHu4yEXFTE8oBI4xnBpaRCt1AJ2iMsHeDt
M/iXx77zOySOTUdgZn9NXtZmw1WMauDAPRXQqLkq+ePs+VI9upGn+ZXs1f1+oanj
ndrcZysMSJgbXDgUQa3wMVhZGIAXbATR2nhcyOVxavc7neVwT719eha+5shkW9A5
7wBALTNVK+FBZO21x5fbHyg5QNxfzljVnldZ7pNwmzYTW6qdYegC+X7P+vYk55cb
3cDkwDGn+jia++p/OQRlbeiWezaK4rskV4X8nmc20PLuOM/AimNvGYkIh66qif2a
YCJLJlJcmAELds8EXtG7gs9wPMRHeA0K8bafofdVSvLoyfQVHpLdm1n5ksjK9oKP
gJBsw8qbU64Ne0A9X4P+OUE1UxLhuHjXAydfwCgyUbvdeJ/azk27v2M374ocIWn1
yeGy71hUtyr9GVHh1Z1JPYG66kcwN16qAw4mny77TQ1LMYQqIXawjfrlbJq3eLQW
OfmYx0oeHvCxA3wPlWTEQpSCcW7xkBslgUldeDIJwMr9inv9y2B5veE9yTPCBKBm
2thFunp/OrGet2N3I4f9cvfbZNVnb7f6RNikIpJDTK9yxJsSFFAfo1llyTeZ7EWl
SA84x8bM3DqezfT6tL/2AsM/dgWybyke0owm89YY/7XmKWVA5KbFG+o1iXu19i0T
e5ggSJNq4yLnqHyQXmYLw0lextzFJlr/ZOojToTGUg3isWwnO+XwV/3kKp+XTx/A
JMfMW3RNBGj4x4vNexkRLOFLJYbScjr49C+FAesycEnohvH+qL1sidQFaoZ4Edbt
IqfZ6t1hMR0p5VP6v4IzgYthFpSEbslOmdc+7N/qkl5X+KnJ2EPy83FledXZSXFH
9LdYDxhhYrYZS8Yb9OKeymGYHEXQ6wh+lxoEmdh0CkOa2MNu0ZGRes5jccO1AqNk
H63OhQ/8iZVyrqYxYfyKw51kHM0G5aNtBHPoyjg5VbjSFqnAKfRHpnPFFHBDKZyJ
haC+cXruu1mwFL/0CoNs73ZpUe72QFcpvk/dz9j3f1DI0lVwYStkPK7MLJBu3p9I
LtRWtDuVvz/pzl67pdblwcu81RaZHtr+s/si7Yl5GMVDUPY1souLNwxg2EEHL+u5
WNXj4ZX91lRYVUJkwb/IvFHqKzsA9TJ4FmNQfy+hwB2sKcp1t6DD/d5R1xJ6QgFn
yg6hcLZIMuvqNq7TbiuE/dNKyxe5Oh2s5C7wZ/UFi8iLdt5w1o7OW39GLqfEOpXO
o7WcnxZ3qk70tnmM0mMVyjwDjHDUm+GgT3jeWfyybxRN9OaNmTj5+f6XWASY12bR
6fl9sLljoc31gdSfoUUEzhY5Rayzn99QkeYb1qtRFHrNnyt/1VLzlZvSjKv0HBCO
I1fVpkoD7y6BkShccxIUWXch1E4kU3E1A0ol6OSdr5HWlkMaFhw2DV4Et10raxv1
6+R0X1/7d+nmUv20y5s5CyuXDcJaqP0iozEENSz3Phr5q9Dv/9eXj/52UEzLJpTL
nqzJA8jBEMmxdC2+KAGtrpgevLlxj7QmmR2hd9khCOkkSksVkgpumHC0zwgrfyQf
j8CR1KbBRIIwFiub/iKfx7HbHiDEJV5Ey/u76fbswu8WvTxfW1sPa0Btf39vrXWU
Y5XtyCnMDrZH2AnUl11C13ziZg15IbmNprS8IRfJAb0ABEQcj3wqzlnYi5Plrc23
lbA/y2tsd14ibNgq0PR3whnkw6KJyV2ZXNmkQYovpZZj+GPF9+R0+V+vLFscP3Yj
koigAXNG+Ywe6UP0LLDfzAqVcVVy651DmzhN48eTB6Ak6h/2lWQ5RYQGcBpCr8W7
1SGqCcRrIDV6povQWAAibFpPYV+vXNXW75VtLJ+SI9fSz7q8iU+PewszTWbprR+/
sEW+9pZ7ULfdDHIXDllSjDpCwiwW/fVTC/KFi2ro3dljY2Ky3m+klFfLO0CNYMKc
jq+9xU7HsNYJVMHlomHDNKHYISoMarNNLTq6r7FXd+SRZmqkeNk8WbDqVExPz96H
3Zc68giBbm3a25pFQB6ZJ+Y1pa9cLFeyMPpUY9DniQEII+lhdFMBePcldxVWtMNC
q5161jAVlET+l4fy8akaxXKJiDx5HpcsIKLmNa59PVqLPYHOYl1P/ZnjMKJc1/ZU
1zWDOjnfnwQBSrN/IQM9ZD4JUyAvIpJFYk5cEhMteq2YpgjZhwZPIxr6PWNnWzin
wqTa3dJnR/KiTziifL+uexpdPNqpJRyqu8OA+XrhqPX6PdR3iyi94qyDpnPGwyn9
6CU7umKp8FNG1PfbDCF43w+1PUD7pF6vpmRfupZeFk8+cTK0yr7+Ix9i2C9KZ5Al
6/2Bz5a3MLDktYdUpXeX9lpip4wYRjASXjFVsz0XxMIYdGYytLayPHdL16+Jh1yz
0/cZvCjVMjuunfoOFVjM5h+0bX0AY/RB+HR7d5rHDaHhHhZnwn2j0v7wgWwlAOHf
DIL3DWflmWDnUIxv76V+V8i9crngah219K4ukUbY1N8E6rMgSE0c8zeL5/+9/aaP
ldELWIAWz6DdPPaoQydKdS9Bu89kVBT9wbBhkMvvGD88C+P8LQAJCpBuu0N3qV+Q
KJpKUlhNEAgoMAlq2X2DyeFIk/Qi28qlvrxMCNj3eQit68rhGXLj7hFSX3StlU/y
DLY0J5b9RF9KHdPRgUjZYTp41NyVH7jeBlVIt7BPA92OOSA5UmUTN7yHvyS5cDj2
CAaTwy/39BRYEcboK3BuPhkQlgui2IzizyldgNlBlrdiI+VuHMSnTl3WoHqDTVcq
EI6XA0mP/Ge72Kk1o3VhwaEM87OLGZ5GMNgJKXg6+SI5ljqmPnCmg40lGY3pKZIL
NKGxoa0kV43MpqFYdM34KZRYNeaUVxV1Uodz2tbyxAUaiV+TcPVcvqBwmRVh/9Ui
PHaCaGjGpwMqwcyQLRu6SvnNKFIYlwYAENl47+vCX2wqiuftWsdZDF+lWdetff3q
xpildfENO0XiUBBgzjRByj1epCH3mB669zkySxsSr4rFkhZjL+Wn3n/bwbjX1rSk
LZnOUKCv779xw1YUFU8lw+HfdqyMzpZBK1SRWap+1a22hBpHOZ2mCWIrfwA1MjJY
1AcrUYuiYXPj5PK9L5a60a6K/h3XeOMFEcHitZNp3GyVbL92jbSg+Q+MmD5NWzcM
EGR4gVyzq09VqNg7AhGFFFRVKkb5XKG2/JMoBiFicuDHXQd5MDuC/tIgkeeRgxxk
O9QWdAhKY3uIeEWV3hfJ+y+pIS7WvCiTp+UPfAaqj/mByB+kKnkEvlHpe8kLOs+v
Kih8lgsetDHASN0jCET1Q8XVdkMBap1oInExzPPjrDtLgJAC1CJMr4vx2OYPY4qO
4OjDBGqoeDZrgU9B8+JWmLdErtw0w4GCxgdmffE7nQ6hqnGt9aSLBgJtX64DviWW
TpsudSwYCBw21WPpYDzmqVOCOpc+1Qhd8mYgIegKgAteI3AnMUeFi9zlPkDVNzUY
RaH0ugdehHtNpVS5UMEAXsQLP+NATTBCurxL0mVnIV2oG3HMbuNvoMOMJulNSb2M
meemKpiTWoFPM4S2zlydNG4E1eZXoqYq35AwYcmFoka/Ex77lkfYFIeThVeHYyOz
abO+ehd3wAQ1YJ/Bg+9/QcS1RD4Fh8aoan89oviXaTVFQ5XimcoRrOu/lSxJZCjf
rpM0+GDIrX/x1yARhBpBbAZVeB1GdqsQ+uxQBeRSst9CMkStqFLZO5OWDsiEt3fN
ka2jxnw+XuL1mo1pI9Yz8yz1PII+7NN5vhJcF/MDeAOE8bTgSVZG/hye0tKkHnHU
Rio2sC/tB9MUfCgr77lseWaoJTgvNzIfhwqPWVphtImJyeLsuJ573EL1kslbDKfy
FxMuLtuSWwJ839ULz8Hy/tgoc8VqsXiO1lx5EaPWr0R4GGRD+FfQqzbQHbl+Bz3j
uqK0UU0AojjzC7EQ7Mf3x2jr0jwr5rZbdgH7KE/hJKeyTCQiq8BssxCbfmm8tTk9
k/c0J9cFSuDlNu5EmDGWK9aj5BJ4+VBg0b0iG+0xC08U6hkrnl17GXGuJYnsiR4m
maEvkxT5nerOC32M+VoLEUnzI5fanaqZ7uBCIXpkqUz1gbym5WJQ4XNHJrue9EJm
unmqmUEkA4MiIqvadEvBj/wcS87tnWS2+Ag/Y89VLXP8/pGZemOS/rjEUy0b/YeL
Mq5kctytvuG/eDxQ6gEp1SzsE550rQai5lUIJ6uwKhWmpETmA3PYJoKYBHp0pewh
emVC0Gm+9J0iuH0e0gVFFVY41ScystedLVNdFscKTPSGoC7+4GYKTV1+PEEyOfJ7
KOH5mnub/viTdkiSdJxS8nDU+wpQUeWeGhVIPGOrdv0fNH9/JEHrjGEQO+XrGv7Z
TTs7om5+V3Y065800KZf3ie8rqPaER0EGJ6DM5xGcuaJQhx/iiNv3gYpj/H5ZY03
upoUSvcx/HQTCeu+njM1dYLrwPESyo6H26RRqOQb4JMkDX8oC+THryQIwDE/kOvU
irIOFm5zaP0l0wMlqVXZZS+ABE79AoRafOALsceY8qjQemQlUgMrxieOWCtzVLmT
NQQcJOIbSfkkWKJBKyxWT/1XSf6oYtsq12ILVU5HM8J93fsbR6yHUp0L06U4X8hU
m5+nY9JnWB/9lyPNHND1f1afp7Pq2oLVnMbhBZsSr0Thw1LzTAZjpyE3waAZ6D3j
i2lEomjDHnaO72XBAFHa2hk0LuoEQkSROQJgblYxlxpeCOffcviSrHPVZcvSNKyQ
Sv3oNoLiXD8ApuQfHxnpnC+27Tiep4zZ3SkCkUYAGCeeZqw5POT6Wgn8BsixUE9i
HxkBhuGYuX5XiQhE9qNBmz3GQGE30W4R423cp07lT0JgI3LRVCYIao1iyUgDIM0R
VkZP+/FFJCL33Z1jjosW0c6MYdsvgEDbdoPBPrjRbQED9woj3aquEt7ZcU6RRwaU
BoRm5PrqV1eSGcuk9zEHFkVPCaO5vKJ16VOWpVl800Vop54Knr5+/LDbaE5mhqVW
TUMTeeplEqhIsY72E00HThez8WUaCDlK0DEi0tpactGXGhHsJL9cRfzwBd8qL8Hc
mty37hw/ps9KSPsHLD99ncH/kxzXRzBwFpmzrmKi8wBIFKLekQMuUSoj3fWIcLxT
BZaOVtNiRvw9EKaZrNOKvP93kOMhceSZpozE2J5/TiuxIlfY73musKhEXtIOalLE
htHoKM9D83Dqm14EffBfnc+HASzwNUtUKmdWhLw/4UUAyoiZ7mWbTTZ7nRtEMm5Q
F/c7H79jTMaGdKwBauWfwlsEOchxYO2/dLgznX/taeMgIPjftsVjsodjNnTUSu6r
cDOKywkfrBTfAqRIpdUlHUOOD7v/wVjImlIIX7czFXbEHHg985j8hxPascQdcElo
gvNws5yPjhPdJThUhrg4kGfVv4RDpFv8ph9XSn1bYAhIhcLogaBrTxIJPsPM2frU
+Xt6gmkzWh5RKUAQhi5OAjbnyBpPSITZgd9YWVukCrGTfPTAJ0AzAB6I+savtsa+
WKWjPVBfAIsaZgm8tHr2Rk1Cr2vCY/FHaLjggif98OLpeLqPEpEGvNJCZDsR0XH7
gEu3pv8uwixi7fGlnHTxPx8EacsuPxyE7RtAGnN+bx3UHtg6BaNCQ72CujtPqfqS
OYYSoNtmYiMwBYRbU/0dmhXPWK1nz2bPMSZuJUvJ0Aa5JGOeHEFgfYEVkeP8mHdZ
n68N31rBTJSXeFHT+ddRYSp4v0PD3lEBJrH0h648uTAfVQ49o8QMVY9tOFvi94P3
OMqRx5uLCt1nmU1QNn0Hfgp6pbpOJ7TmJHDGijQPFIGDzBI/QQbbz0a2twNBrMpd
1HfnBvlYb1TKXPOHx1/9zos9y9NMJD0UqYidQSzwZu9Q/AvGT8QoQjNFK17mavGc
4P9uN5A/gDn+7xYjTTlJ8JBLTt6wZi8ZOxQfDfVnSL+28OaBHI/wbIaYQgHoQBv/
7NLnXms3tdl+V2wxjDR1Hgpza+Q5B+LQfWjsYIz0x6nehL4qIoyYwW8C316F7aR8
Kvodt1+Pi1RIQgVVzEdXq17NyR7Jcg9Q4qLkn9RkLHxp6SUaKivgvuHyOWXFmW56
7ym6rdwB1GN0gSx67VuXcU4Sy3oIUNFWp4hJtRVhMv46mkhOYeDOvLATA+a0IgBF
gARZzSVMjdYHF25tvqv9ZhqkGyVhgjzgW6ExGa+oLSEPbfnHBisuNan11GS5tLf4
O4if98n0ynQXM8vy70pim8iquC9c7OA2CBRH+7HV+QE55nzBgwR3+qpaed4qX4VV
2DkqmDKl0xtvc7NojgOaddoKAKlaa46bZsvYZbFmqaNcGkcea6ZszqbOon03eC/H
RwZU6isYf107oNlYpOzAKyx7lXxbf6ErPGggU3Lr8JUOEPbKLkhWp84PUZBLmgpb
WpX558jb5nwctzikY4DApV1sAfIjfuScuN8UpkT/aLWH2mJhxUwla2jGIBNwZNEU
fq9PcN71Yi21zhkmXc2nKP95NVvZmVLqNQjh2HHXeacczeKMtOHur5Tigp3ADkAJ
I5QYKhXyeNlJ25xKfZ1mm1Y46V+rz/P1t0m0RSuiAY1sKe2tRM6RtwQispQryAFn
8A70wLxo24dgO6JTNmYuH958OwNFkKGjOMmf8O238PKDMp96nSbgw6dRjoSKAAMw
+Ksrwu69BJ8d0vVlwGRrQNXmRy9ydhNnbksfReC+KscpNZkJxVECf3S1qfLa+eC0
d3CT0ydR4Xof/q1ivezleovwXwVwRIqhhvFZaK0PGCCcQdsszr5966SRhtwdGHy5
1xZJoGZQRhOLqX571jMp7FQs6A30puQYpLf88yY3hhZw2VHtki43TZqTB9Tn3Bdg
ZfMlxg9QVkWyorPhXL09FETP1XSpcLe8GLfTRTXcEpUFkVrsfSovIeA11rDGGpAb
Y9AxQVFdBW1jigTqOZaD9prrPbYjTDZ6PfrC/M6Zk0UKItN2i+PzOyyWYuh+idTw
gIDPj/yaEy9jkB9+xQf1bO4ErturkmpiBWS4Fbz0w9aQspMRJiB+V2Qj5IeHhwfu
af+qBvzVU7wxpIX3KqLSMX2bGGLi8vso0i+lo0NEPxu4jj7jj9rhj4eeIJGvUknV
PMJvb0eNGEMg2rOAaalmeurG5g/IoiMnT9iJ5kbxNkwGvTJtTKcSE+ohl9ePmbah
ZETjwX4uVdJGP5xSq4aB7zYej6SppKzjZDtoEN2jBUyVR34mmotobM8CyvrZtuN/
mTD2L4F/8NMLxwTLs9YMKnWVymTVrREe4WqJghxWkOp6CuhJvuF6SQFKrMkLP1lK
uZa9I2NtZ2vSvMNReaEQa4aaGmy0ik9M4cUvD8PGIj/5cWrbArWgLT+JId1htq65
9W8QmSf1ov8rhF0VfGBynPvEgqjWtiQA3EmPOyk2HcbjIoRFKfMieCzcOOX8zkvR
D2qWc76SJD/u96e7A9dSe6urtN4cbUDyGK1PYjo0sLBIsBs/OOAf7IiTJ0o5Aiao
WCEOrOwJ2IjUdHWocdO6Pe8vj0NCX0BKnjaYJd9KwY4GnnHRlUM8mvd3wdhhbO8q
5cV8tnhG82giVb9j1DeBtTFZ1Xs2jvYvfyfSbZwx4mzqeHdFCHarlSt4/d52xqEW
/cd8qLKXeukwnV8Fol3cQ0L0osmdf9ITbBkUnC2iWRvueA3VaOiFNosfuGY9cae+
Ll+gnFcDJf35hrvjpzck1u6JlQ7xebdAXs4436NAixv6RHCroW/lxNaE44nbtIGR
WqOAQdk4KaF63nEOgjllmxkBWNoDPHgTRTapWowUSC5zppszAwh4oGLSUuoDP7IS
oNPXukp37WZhefHAksYPKnTnzoWCU5FAa2KzIeS2YdVhl7rESFrEURXxOTcFc7Ks
zaDnggPxXfezfkFIYUsgTDFmlJIY8NZvR/29KwOXBVZ8ZP+GKzZR7ieruLKtOgJ0
O/phAtigyFTFRByT613mnHv9CedtgNchEMHWiUt3ZnueTNNu7IdrWgEw9wW3lvey
zIwELUTp4jltAJ0tQ5JAXLUESqlhJm1zH/bTUhmLqr0+ebTEUlqtK3BrmFAgkviH
pchv4YglPrt5kz3yVWWLO/mbDNR38h8Pu2R6GGnBBBdIkvg5NgVkRZ6hCmTDN3GI
hLe2XlLawlbkO/HZ2shpM3JCqzn/hAFjtg2rF/+GbuB2el5jYsiigruOgvkiXZl9
Q7znok6/YRui3PDb1NmEI2XdSy+KuAh6/jgTsfYaNDIm0IcE83/L2Cff56VZobbM
EDTVBioo1gn1AuhgijZaVin/xX1UKEMo+IAQUyg2etq3Gr9jmKjh6W1tlPlYbvn7
H3gMPhPkVa03l+FKRrxrWVophVbCJTSEwzoiRxbNW5TuLcnUF5Ad7Oh5TTKCqrnP
yE//oOkVjBBQEPfG8tbn0f9Th9QUbuE/xkHPjknMvfrDsNUzG2pBA5EqJfLHFvHC
GOgt0x1gsm4YH+iy5gow2WJGE8kPfMixiuM0J0J5LR5eCbhA7uCpnsiFP3AH51lp
Z5K59AULJnJvKLmJttByAsTQZGarFk/ba6Mc5CCgM+TXc3uKNxFv/dm4UNway504
hgF4isL/R8DZrdPFR7se9EkAZU3Db3m1pWstHxJvR6QGZbnSvyWhfZ3PaRBFRixN
nhCnDI1wNxlXFCNhm7eUlPL49CzewOHRlHzUiS3EZnSVlRuEsgSDxun62HqgzoBQ
ySEsg+6xUsWTnmq6pP075N6qhOrGw/NmlUASiBUWnYbIgTkCqMyzShEKIq1xMPf6
inUb6IRJBBU6WV0b6tuMbVX3nZSwiGyiot/cOku/Tt0IX0NbxJJDQ0C5n6Z0csAU
UyNmxh7pviSIMaJgWJKnia58BQrJLvAOTRu7KcSSyEkk1a8fwPBU163lbGl1+R2r
9qrBzmpYWB0HRKtaznc12hVhkL/q69g5aBOENA4IYBephSblOygcEJ19+cnq5YMF
VRsc1MAZlypgzLT32G8+VCYk5lEWFunZ8EQ7wv/ky8IxOWL5fZDL7H+7xpiHjtDY
4zjGOfK05hX4ErScvo7KiptglVmHsVDB/6j0cLa48YS9ZHU3QXL6yCy38OQL0brB
zrWMoPmjkbBYJnvj9CakGgG+ZYYUq7nl3fzzvrwX6fnU2imoS2/s4zK5Sf255Jzh
U2PuFgEJ7nKIMcJY/VqREtqw6BkspABNrxzc3+FP8CnQY8LtrIhCxqCEZpRVFND4
GcOouDhQcnHewLhssNwOF2xls5nWQAhujv9xphiwdJ1I5mMCdZLrRi4fKG0P2Qer
NaFLtBhaD46nOVwobM06yuq+ncHIEcaiamLhdBVNbKX/zoVIDvsKHCItJiRmrvpL
QsejiuItFRbIOJsq7MTBE1YTM9VqTkEQT+rEbe58j0/e7GtKirxjz8Qs63B/YYjw
lMVyyiPc/H1ZiqcmClI77xZCQh+H8AsStRkSuUMJGW4JUmi3Z2eDVRlrkwV49bav
VFvUEMZf85leEfcWp5A9zMlBa+pP5XsP9Hqu1BT1fWKmCfsiNNJN6k4Dry9lbq1Z
IKvG0V/PfiV8b8TTIKSX88Gz3SXALevpeIBKaUBvdMMAnrABIpM+996l/TbeDMJR
grEgsxnrEP6sfpVxWAEPkLM2XL1VmUyo1DvYAKHwgW7YU6vmdmvtv3RoSpT0rRzx
zd9sRWDBO+X6SyXUaTwqQMpDSgPpBAc2iz8lnNRTJtYnXcJWfvtOTbbSJcpsEtKN
zTuGZY2vvPXDZNVBY3a8wBAh1NrP3ODTK2nLyDfUeLf3A5tLBFKbBUCcxXbgp9Se
jn9IPqBqP0exmTztosylGs+bOLqWSTTxT0beS7sEwQkWt7/w6EPM8gebIDlKdK+q
5AhkSZqacy9J9kPK2V3ImsUTysc7+BM1eUORmTP0BZe4MvjUI9m1Y+yoKwZWFA7J
s/nOHmTymekiaXmP/UJJs3h0JumHBQUBAkXEz9/KvC6tOhijJiVq0Keu9uJZcpUf
FxzFe6SieFAi6hxLYusfuvnx/erGb8H8O/fKbR40cLdJ1ygJCTYvL7cE04RmB/1R
iOv2ODK+MnutJuTtlFjkwewnA9s8mb+eMfGpsu8sVJE6OSVFuwjSXfNGvzo72cWs
+AF1fztITNRja2vRO+MfM2pmyuUgovfnzk0wLRESfKFAwkP85mmW/LGSSiZdc70M
1VM/pSLuBAtvYy0WxrS9U91uxUqw+wbqJC/at7oTZ5AoUe/Ys5ojNZUN6RHJhDlY
N3lJ/9SCjqQyavmH7RPrLhv3rSIIfjJOWi5aWy17//asy1UGm6AfiVRC2tO/qpER
2qZc9mFNfBnGDqMFRsW7+AHXM5bHQ9LMBeTuepTbxYxVG3JI3fQFLLnQYg+aUn/v
qtE4U2ZKY69AABzYGmfvzly8ePjNU8bxa9hrJ3BYCwCab2E0T5cRVJIF09D7IdB3
jFKwqwnQJROXW/wZOFJ511PvEZT5c7GjC/Ar1cZolQwBlE8aD4oMESxk70DUIn9E
NrjGsbknEbGofh1805PtrAQM09cfNh9k+oifyVqzaT7owowKsZG3eQkz3FjQLoJu
6/gC2XkbLSzJWqGImRm1si0ui8HtxbTE3oigJmgIMQFc+YCPBwlt2AXVnT1ztv12
KH0YtaG9u1HzxYtBFCBEz19kYwafcZLpcwwFA0pawPcm+mpia2+LFTHs2TxdwY1C
kkwNNVcgcKRKRiyXHRbfax6KugWspWR7CSnK1t05tDCXC/n85Cg+pAoVRMnt51LT
PkaAqKcGi1F6DmGkd0gpdSOXvVphvDnqi0bUd9d2T/GaN55CzEAKnZJMRmg6bwHz
526V6S7Oi1AG3hLrwizgas64JvwwVNRAj8PNmuJSC9jXZrmioKd9YphnByWHeE7x
J48MN93zw+TtNL+CHaO8pe1GO9t233Z8U/6oDbGi1rbNB5WnhKF6oveHwmfmoLXY
P5UBgQpREzLAveub9h1KBWraoDfL9oHms/IG5hghRikFP//5l1XJvv1P4ftkVmJB
gkK/u0zQc/+NgW7Ry5NF8JoqqMSCZ3R0LuFLLEoSStihU8iaoQCP7QJerXX3nNmT
98B56A42UM2Hhgtp9qgQEQBD6MoPBDQ5c+Cwpm5E2bwOBKDxmu37H4+aRm+UEXhh
SDCmJcKMRNfBvyJL3yqgbnBXg8u7Yva60pmd/BlgesAzgHP6fsm1+DhqIbgeIaW0
`pragma protect end_protected
