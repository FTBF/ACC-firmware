// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:58 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nGftrw11JPuzN+NSElt3bixslmsa+QCw92PuosjlF0ClvcTIyMxf92Skeskmb3Wt
NiBruiUauKFgyPPocF/zGJgovO4sHNw+4fjVrz8lnbOZhPUaWhD+SIfSmXateac7
Vml0Hij88+vxCP8TJ1mKlsWg6uOtyoMlQF2a13ufJFY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20976)
+0ZD1h8GwDTwzP+MwINSKmTUu2S1AuqeLADD7oW4kVqreK6v9bbx3G8svJcW4y88
kieQdOQZBEJixZY4j7CteIhI9dAydD1XwqP6njlaia4v8c1jckMnvhOqhiwSH2ds
MkeVBRbwjtbx6anHC4NF+soaYH+1cyH8u+ltAcmnSH8/1R6iV38///7yN3dv5lzD
5YWvjr6UiHI382ySNtDBGizKlMgHH5UY9yFYYF1CuV4CUIzom26WyrnKmrvpBePm
upR4KfuR3U8VC7SIpm0WOPsJoY7jfLYfiCXD5P9nyNSd6/KudoUEauM4EDvt5kip
TkuMIC2YdUHyC2y186zknJ0dovCrZQMDjxPy2AiMWNXHZpFfxwr/06V/oq5nHoAY
N+vLdGvmrllsmVdyfPmBzuxbSSI86SYxuh0JBzVd7E16yG+6psBedYVtuunffkhs
mGCyysOTd6vWthslw2JFdlCZBNyPoT7UD6A2MFF9qc478LlDUDbepjO0bOA5oQNz
mmnJP1Z4f/Mn39/9t+jsKh9Zy4dmvkW561F//5crZW8pWPcDZLwe1E/Kiszg2tK3
Yj/nNFwQkIAoe7BBFOW6P2r+k6TObApMkelTXRo7Ow+o94WhtlTnTWVcLDUJ9vK7
+uhA1/SnxvfQHoYQW5ZGJhNTyNU86QtUL7buDlLX3EDOZ2Dco7AZpN8xaJxatI5b
DYu69/YBAbG1jH687mC1fNwdd9bZ9upsbw7d09GqhXp1BZPt+Qtq3yi3c2+HmqFu
aslvVEBnYtUT+A4CBie2BpRYlokltBu3r+AyQ/qgzmNIKZcnORJzp3jv1WVmmj2x
DpkIPR/1e2NDjhPab9e67ni6pQFShYlbZqE6EFMdUZYqF1nm8/6t7iEdvgy59T3c
BlJhRykY8VerYswpdBYPMhSkuwbsB6sBKqKRiJUaxn2sJDkwMfIp/N0YR4HfCwoo
U/644Cb5a6x5we8HkjQ7LplmYwXGU2gn5oX8czScN5En6NfUypftQTjAudqe0m3W
OTnG3o7bmZ4zCKJaNwNLs1Pt1+wrs+3wSnRmc4rf/GZYFlBrEkivHIAJ6CkLx/me
3QMthkbzrpv9SHrP1SV7o2mLJzoT+n83mN14OrlCFbl9wfCr+DiVt1CNY8sQ8KjW
jauhjGB089NgViottFhQ6+WzQVUqSkLjxXDYMPmDg/w2RxBCOjWiKSkNORGj5n3v
2fX4i46C4Ag564i0yxRohSimY9zR8vg6pmpuWpAhv/w1bm5YkYd/j3Lj1rOlCm8g
07LwgIFMNQSPLcymVQxgUliGYhRISbGHGQ/Vl4puxrklYd5I7uVlG4eQDy/uzBYF
P/98ItAjs1WgLRPjSm80FF/Bai4pLgpkWglK93ntp1JUc9NFA1qge1QM7/MU2lTo
t1AFvaJ+x7tMSvg6KaBYhcnEwJKTJW0Yt3py5aSbbqI1bm5MtGSa014H5PoK4z9E
g4HR2cWGSHL7mVlokkw0hBW/VDg9KL1XnW0SQO8LV8N8pmd2ATGsGHSN0O1akJlL
uM0wMkkj4Ok+4WdJGrxu+VndCuNTAUdsRJf/8XsnNZJ8TUAurn3v6GjQkXaVA28Q
iQZ1elKObdKXvW63N01paMmsnW/gIlXHP/PrfxOppDlsCjBhV2cPYmkVQ/4nRA/s
3CJAO6loLgd+1PO2NZxBUIQXsIijTW0f9yZwbReSnGMhiTr7TgZOgmmN9/9Z6kFe
V2+wfb2YyK3hTnf5/OejqA4jwXfG4hJi4E2uzuSgyVbn9yGpCneRy3X9YIMDV7W/
RTRLVTtZ7n00I4hhCRrCDRIdzLB+7fJPtZIiYvBvgF+lrdhpfMpTqykLzoUqy7/7
ePy4iZNFTNpuX2lDVtNq2EOUr+vZRR+HpCq6pWw1r7hNcXcrta2SyvsPoF6l4ZWA
BbABIz8JSFeAcYYF7VzWqjbxbKkBp9If39wOqyGvUsghtJBtgBm7J7fib/CCb1hF
ruhfAEAW4bHP7u64Y0tiGQGaQq9TagylBq1z6gEbdHA3WejM8+rVcuv1YTcFl1oG
TbxAHIW+NfWT/Z7uxpK6bUUz6OzhIBRyH9yphP/AR0RvDS2m9oC3H+xWvdki5P+J
84MOx0s9qwdobVpncs2uV9Pba0MkJO7CBhJi72EmmR+TeXKq1IY3rmmv22I/9+d1
YFUTomAsVla6Agx5GPr/PPfRF3oETUCKCvmLw11GmHJZR3YDscbPly0J/9L25Han
Fc6BjGrGBMPZutOOf3OAi1yThapzukKipR2eVvD6vuDOEAFFZt3WzKxEOZjibplh
uwu+XBIO2fOiMf42WhaTeOo1hlqTo8BA3cqNYxdd81hkmHSE6rx+gqqJduxKePrF
PhyQx3HoGMqP5+nZbi8MJ60o42aWyFKjeE24S+ElIm0xzrVTsSe+L1rnpSWN7rcC
OlpxE3BtNOktmKpCC5h8UPzw12lDsGGFHImH2YUSgVQd35QhQldIOQVT3S+3o0uy
OzU3teNgtQgphYLUMDEepOVeTiAq2jkNnoIYBKEwMpOfMgq3hvgxjKF0I8hcsprk
RTXWT/kFYNSu5nxZwFPMHa5JcfvO8JYa0geE5JZc3Xuxbx/p3Fd6hwBDL8bFMNKj
3Dohl5kh8EMdriGFyObmHjTxKF441TqhNn0My8Yy5cN3gFz/vJO3AoeAV7fskUGu
ELLoW+tHXnVV1EZx6N2jYg5E6qj2cLXqZm4xGaCvQztXluosPCnjqjly02zqW8BG
YwJcREs2Prk/WUODL7CBp8Rs5rBaJn9hto5X77PPZrPloU1WnL2JGhYloNnd0pOi
WuDlYTi1p0pxBLJT3K572SbtbliygQdOiFPSW3ggr+khVTtBV8P7QrKIgJ4WypHP
KzgoGsxyhxLF9PIr8WZJQ6jWnXVcO99fRg5yWrac96n19VqtL9hRft2weeiqeMy6
KmtQ1kHVlceG+xyvjF8t5uGqJbeVK+t+80AAjkkqEsqhUfwxDya3XTp+kwyY7Uyc
PkCLB15m7fjU/EzAup5pPux80HKeXBd9Gzxjm0jlhKvSprtnH4j/HRi+xnDbGe7g
zNHgdGOnz+6V0V3fIWY3/yH64BGmJF+rjYLFnKwO2pcFVFtwsXosqchoSqP2KeUX
+Pmquwgjn1L0zG+Zm0jQw54IeJj5Xp+cI7loIcYhb2qAWzQHacIar6IL1wqvQ7It
J/9o5CaAhh3DmU8087SfNda8FLgfiUmytGdYsiZdsd33Z4MOoKkGBJVbjJdF+8Od
nKAZIr1OxfRyb/icKc5hVVQcbNzDdcAfF1tJU1Q+9evGbxMdl7zdcDS5Rk6CXhM6
twtqIiGvSM5U3NkZAvJNoqrbJL5r/U79kiv+Q7FE4CDKCkeOjIAPev1QWpc3t1QF
7kaRNPRyPBkmZA/d0UTED1lhSyNtkzmKyuYP99mRWBB5e1oNCLEfT+TgQegE37T2
0X554q6UZkApJrUodFOgH7OcP/hPfAJRI9o8LIEZ6j9YXXCueSzqsRd3RQ2REF5N
kkKEJ9wkUceJt+6mqVHM2utRNFwnxKJ0aWGIkcRaunbMHo0fju3Nb031PC6cHoFz
8MI5TkSViJGRtGJ6sPbz4U+06IsAoc0f6CmX5feRet1rP7TZcCrwQz+bzVR6AYB/
Sm0WgnNcOnmArLsHp9gSq6h7BZmMk6wHNkM7yKvnxGSfcMSPVLmW3i3bx7nXUFjx
T36SUqfDGyONypVXdNH5F8NrwGHprZLnqReAxpTlPlgQnMEeRQwWk0kKgHBWAXFW
6HcJpgJfWafDIX4NusTBGYPBknFkPZh/W8hPz+Gb9GywW3p3SlIuQ/tETGmp+Spx
ULp5EY26Gs+hYBZ7zqR0LMuNcEFcBCDWx3smaDjroAB9e9osRQrC/8EfJFPVv4fd
gu9l+PCeK/2rHHsu1e1C2eyvBy/L80miVx2t3IqaliAB1+6mYrcytG2WuX05gHwd
IF69K8QmIHdcYiCV8rKXvQWMJHNAMBJjCaoWZ9+P0G6WpCcGk6zW6x2tiYmMoeh3
Cm5ZPUhLrqhbz07fs7EM0AxDZksjqmCL9HfhLBIBDIWkq1gLu91bPrj5LfXW1P8v
bAIDuNfAiZakrBZ/OqZotu5ZAmKqO/XEIybuOdxpW91+w7h8uX5Kd7ecj4EprTv1
jJEaxIFZaPVa9PNoWL8Duml7CkfKDY6plbHvdi1eQXGsu9CxU7YidU2gKwHbaXqS
uw7G7kqW3ePCRWN3ghROdGeVGNjx8l4K591xYshIWgfjvoi2xyHh8M5r9Uj3FYkD
dzWNsg4vZAysvLgDsIT218geP7iDo0BIgIsTpjZP+81WfvtqiT1TVVT3bxv9cPzL
6C6jqYO/E3zumrlhgQhnnA+L0I3PCLzyWrRSE2K3YL3cB9ELLo/vmGYeTINPtZRa
tFAV6a2OSGTF3w7S5nMp6BMy7N0wP7iwMZ10kva42t6rPsfRsveyXG42LxA8ngcp
ksxh7PxrtReEpJs/WQ8yeUwabBc0f839Zwr6Qkie/8jVVzIR5vvjQkqgP1gXC4uI
SjM5Qy8i11ml4lagSnqciinKlFq/UQvB1rcEZ50qDD6hKFj56Yh4CD2Cao8tNYos
eEpt/PnF01gyncz0ZvulKnB2Vu2A8fIVM0JqmDKrKMaa6mVJhR/xdZC+pt9lSqwP
mt1+YzYmFsbND5oOtQ+dDheeGhUTZParFezMq4EcRjOMvlnZ+VqRk3wznTGpgazn
i7Nel3dmKODPg1niwj4lDFU+rveSABT0MEKEInd2cHJ/XeWirNuniWdKQhbf5qn9
5Yn0uY03xdY5tj/eRWEfv0aN6PAV1zazKTHYEJP7YXKxSKsZFKsksYSjd1XCivdg
ce0Kg1BkoN3PQIR7G49ECc1aaFIEp8Eox2xcjzZDLz/YvlhR1JCJDR/ecSAhOr6l
U9/G4BTzo+X4A81IvVz6qwZJIUcid7ewm6XSlZUvC5ITFAqotxgWCZcDt0zmA1zS
8AgvKKy52s3c3KbSx59aZ2P/HTBvR5ujv7Xkug4jI1GDE6oLX4PjyUhfpkTDbB6S
xJvHxVaF//+sYXlVqprvydx+CfSfNL6709pgaH02DPNn0Iw8RQ6q5UiKDpHgUb7u
bR/ZeK2bm6rQsysKnSDmEhbV7mzDAZ1LthNzfbBVQIGUSqdAp564p1mtukBw5/RM
wUga/M/9Bk3U2zOcoJjBeagJcXM89C6lFwsCnMVuIcVPrdcLHYi0KFrzl27H5Ydp
5TRcZrLXkLluK4SdMTxjbttRWSoeRDBI3JdsweaSJy9LQMZD/e+7aoHuuQRCWBME
13Mvydwyu4vlScGPC8s8Sz2y8s6YA+0a/sqS1/3bHcD9VyqzLHsb/vlr6DtSKa6o
TdfoCRELOiImsNeiZ5ykUTLzq29iYhbxzUkqqXlDTTH8w47yHKMRiYI+LNzSPxgP
+2Hy53UEfhKKpkgx9uFFFPVdMaN1sHse5T3Yj223iPPIAxOb0LgdmFJIHBWriMvb
m2aN3UTZ9nk0otVdtvbXYVaS+4aJSTzwYyiT6qKxaK0acfueeYGKjnuJsRZwBEci
rhOu7jSwQrNRHIHB7S+eqKusmIMzDD0j6D54LmB/LfnD9kt/64mVbNkC9v4jetJU
AK9rlw2BaWTnNYq7f2ae2cKzsvTpu+h1DQIGxo1BTj21NupTpvsnNmmyQShVhO+n
S+F7HwYgH3QU4lrQiflZW8LOUsU0lW0FE9uKcUsfZvurMt28RwX6ZDocnjS7jZEy
XqPjAwcM5tlCOUph4Zukix3Zi/HHwEVF/VFiZQI5QKaBn7B1BzSs5pw8Ve4uMMsj
VbNgsENG6/zkEF22RUfDQwAZDkZZg8V8BsVplSYLGkaGPiz+MreIc2XwFD+2stoi
Nei+AKZ4uhrXVAptf4r8IENbOuEj0yh/udxjUeU4Ie/fAZd8Mu3f+FjDP6c+B06d
caIME49cRA509yFzATLfFfG448oYml/hDASC3cQnURfZ8MeSTIt6dHojyDNcTmEh
8y2ZYTH5GG2+yJvy0A/N+yp+d8RGxyEAtemmoH+6XZ8+9L7wAkPEaxUyL3QRoYAU
ydZx3NxiCU3Qlu/c8F/bDIBX6LSbw4QIwrj8uwUFJY0bP5rXMXMuNnMiqf6+trQR
I1xBOcFJ8E3Y4DDFZaZ24Bfu4tIGNoWn3ovzKflQAZrny9ooMeSl+Z89oSyoFj5b
e0YhZv+do9S1+KnQ/IQgTNoPi2eSuLQgFcw8DIp8/9Zz4e3bq0J4XKQQfrgNsaL1
1EnuH4WwjqLSqASZroEC8fgQDRVRVfJWxoTIhYch05SWzg7q+n8sn/2TSwVf/zGN
B/o3m58Pt1Eib3K2uK3BfCGW6X2xkWQGyHuT+a1faR3h57nh5xtoNKXmoEL/IuAL
EBp0untpmfYcFjQrvqGG/i/7M3iirtcLybuKlKnfZoLUG+q9YUIQ2rppvlceWIck
0yo1SabfTmOK9cPj1OFSTah6tbdMCv04+DbhVpgNnlvvy0WlR5QwdKnebELfljQ8
9KUwBbbWNTvGy1aVCuxIxnL6xkVeTnRg6nuJqUflJlhgNYTLGM4pvFiU6ORoTPSb
mJWO6QpdSOXac3Si18u1vPinU6gvA+v717UMIECyKzHOdg4Uvx9MoWET1+uYhS23
1t2eBfm24UwpXLChhCWlm9uWTN8A7qKqvckGsVX9qwfznbqrgGnmZ2gpkJCvDkhr
d1P7Bs9PMWIyHaOVntO6UL8Ud/KULS867vcFyWwHTT/HkFoI3dOlhNRNjMgQvPIs
SNTPphSCmG1OQTY/RfVZq5HOX4InO/wHXDlM5RlmNbshxWZl8VPO0MsV/TOqueT6
MeO4msNpW4TuK39ZALLQgMzmaBUU6Gk1KT7gmfgX9vh+QDXLBFIIXShQAccdl8g0
IqXnbkC9Sc24yLVnveO/Ne1cmaKiFJSxNBDaH3QBAY+KJQ9V29/R3nKOboZ6v2T+
nRDcQMrNSY+R8gdk+JX/gXwUQ7SIIoOnakUSJFXl/w4QSe+L6n/ZDoMbXhC0GmHU
0pj4rKLKmJm3KUW2xDEDnwCVarJc1twpknyU3nu3fMt/3IOUlcgzRAp17FpOxyNe
R4+GvIXLego5dJKZ3AcJE0KVZMrbpZ7CTsoFLhpOZSfaMl07/yjsr9SETDkXRyxu
p722GRCmR45z6qPU3OgSZgicgXNJXDM2Nw1DhFH0uNfO0BuAnMsDk6Zm9jV2NEGU
OV5iES19M5nTVjQ+nSHkBUi2456J07ucRxW/M+/u4S2oBegzyyc04ewkrScOfsyZ
FzQWUOhKFlAZWlxOViO/Kpm8BReEPG3erYiHLa4NirtgmqRBdcBSGmZAyGZ/w9sS
ehf6izxa84RXTMRGNPkbwY8ic86c5m0XqLQeMgAWXDFZtP6XOeGuKjacrWHjJBNs
eb81k5s6kYBevzrKfiNjFsFGt1U+r2qeMi8T+WWGDNFjhd5BI+1u31rHu4nGLW/d
9ccNTQAdLB8eY6wIBDvRBjeC1fXpxh9Jg5ZGNJEEpbu0qU5+XAUNSdsJ4O43ybF7
EvIi+/maJ6gSPU4+ne6e+q9KRwRZufIld+Ow1l0eCOHyXND0SNx/1YWaOzb8IanU
I3iegiYeQWJrCcmWPYBvzO+efo8Q0L9P3ogsUMbaZ4FGH7wa5WWDOr8cilYZmb95
FVEPSMuzgF+KmHBEyNDY/2KY5Wy/jwTZS6pCApnC5MIDHupLY8wGKKL1+qvhe09h
I55upFQUHZ+dApaKxN4rwBEcILhj5Hhgz3uiWNY9AG1RvDkj3l3l88ZCGzh3jWrB
PxH9QdwTDRWkDJOSRp+JpbvUZWrnvvfgZiuw6hItzviPnm7qRofC5wprBege+cfX
iS38qtorubtt/Hl1drsU0HDqa724K7XIJdvZbEpTOx+gH9vg4qCfbcgwDbqx/Hpj
IHoBe6/dhtElc50uCMGacLPbas4cXYQcv7HruLO5xKZPESg7AeWFJMsAPfjUK6hu
06AOJj6+OTYEujoIiUQaxKUmuQb3hxSOIWjtqV2RyIY0rzwi6rPm/170xI1HxsV3
a6p7Rn5+SiNcUhO2yDPyfdZeeDrwSOOvnvsDWZksvESYFQntbpz+FwU71VarLJJX
opz1EpQlLo1ZgysHz98KKPxYouchUN7smKtu8hpeECpOPh6Y0a2YntQvsDGaxTjF
lB/C13WWsqzSneRDD/LRgDASgTXwyDfN+79kFSuH7yqc0ILfZqZ6b9nu+kVKHqpv
p4j1JdNY9Pfvqe5HMihDV1723BBsX6FcjjmmbvGpn1Jc+In+uwSU0IHB2gXKtteq
FJgjNMQS07ZuTAn4n7sMsrACSWyNIw7tiPZkssLujlKMESKLtDOVtkEWjiu+gLjx
I6V7ktEMvbAKzCL8Mvr2Luf8aMsJE9cB5kRXAuy32MXV0z7nknjmuAQA8g15Tet2
RJx91JSBMKOYxFOJcsX1lJIFhtMFdu58HM7GliODI64Eg9Qv1/hxa1rjZJ2BAW39
dLds/dYto30T5mFD3kbDGgo+jv+1u8nXRyKkBi38Ep7H5pDE/tsjEhUaqYM26t2Z
C9SjrnE/bflNk6hLradG8QNrHgGE/+KCdTEt0FtdMsIw01k600YYeUHi0c/Ws2kV
RsCDfUVeLbTeSK2oWTjyNUDj9w6+L6gGSkUVa33oaq3RbQNl3YDutavHXXOEVIro
+xTjs0jpwbjAjGAIOFsk4iHxfElkb0E3FFlHW31ZVQDTMrNitw5MubpKODKeykbg
ypprVcYPF5AfxgwbmCaZVM66m/5pAYKC06NSKKq7kEqZYlGKuITkS8BoZnaAVHx3
Lz++6st6/h8UHWS/b4uUUTEIm+AFgISysV5mW0ftANVwnL9m84dbh/UbxNBr1OHL
HsXHgPSS7akMsUjrreSVVy+wFYbiaD61PgWnHOnxGBpR1QTA/8BAOXP/GBz6d3IC
vzSVz6RQZAHqcf6yQ2dPKDZVufxEcbdkWY+tiBUcVVdSYDxU1a2kDL5Ilcd2z5cD
uj1mFy8+aTKzsCA7uQcCWboB3JO1fzkVktDARXa6AuVoOtDR2j0+YLKsOC0LKaPi
mvj92f1zae+1w4y1Ww2mYdDwHY/Ig8n55m7QIUQA1hOizV9mEi8TY4cNOvA5g6ik
nsinIWQVXfj3KNpMhOhd0KSTB6FeCp5Dctc/kTGi7cEAHlxYAbmkNpyq7bAKvjxd
IZEag3D+3aqZKAfl48X+nremtILmnm/A2DDf4hbBJWVMSl/G8PAjavGxRAkrD8GI
88gDVIird4ywJ7wX3Z5Qi+q92A6xdG9Hd2DChFl917sAHaIZqlPiqsoz/ssnyaJN
Yt+EHtp/EYNiea79szMCydcvV67T3azOPN1aiib8Ikp+EojAGDfOks1xgygXyaKN
H35hClnPLHrWIOjwqQT0p9Zo8slMZGkVOj90qzcEDr6wrQNY0LBwJp6OXaw1y3oh
YVBnxt2jN/PxK06LoldQNYsUaL9lSRgZX9llmN1Z8suE1GnL5R59XSxeimu1n3xQ
tDLQ10Rej8WqcR68HYPlt4kzcIyaAEPaJJwxenHZ3FUsojysJ+MhkO7l95RCeL2e
ifmDUaA1ZrqFdWAkTHmNASekt4mSVzanGcL5iyTQrYNh+SmligmZsxdhHkWSt1IK
TR7yf/vVARX4fipx5ZY1/PbGuNu9gqXRpebhQkKjed+7B3ViyXaoJFMwK1u2Z5Az
0dGQYHSNXWD6zFrWRLhk1xxaoums02vlGRDD5yL17qD2RAvTEYZnaWOTEqGPEo+v
tQToSl0LarXUV8R/gHlMCQvEB5eRKopMqReK2G9TkQduqfJDepMcJ/SIqaEt3plK
c/ttVTim4BscR6hORcS2zbSL5X7GZwtWSwfNhWUw+1DeqTVmNSiOSe9qAFR+p16z
C7NlCNz/WW5dFx5QQS8Ll9KUJEAWDP7cdqe8YusGotNyaduYoaHOGFv8T3xspDmm
xRLh7PF6kZiE4czUiPXiBu2Hf/X08y0mmtnc/6HU6JxohPXZNy0bcPavvs40yTkB
0+QvBXtwhpOdgYBG65FKI0bzKux0YpeC9NJ79kuEbt+HVr5diLeFBAeDrCZ2gj8O
KddzKCgJ69i7fSIL2Et0JuNYEDrADCHqg741rG83qJqFPFKA6+cT5B8/MdoDC/oY
AVRv+k0repWIke1xjc95go1Bxnr3N3uxpWCms4mFfsm1yEgXdxEwpZSwu5YL1mNK
5GbfwMyttgTOLCjhJ62ox9vwtPa3TRx4nDizSLWs8ogvXDL24Yas/ujGA2966ojZ
hc677rI9dOBnR4m6wAhJJENodm71pKydAiaG4ysfDxXiZ9b8Xiyo1+MuIHValZeW
/ut6UdwT8iMCVUa6mh7OkMD7crpEF6GqbEmO9KD9kpNphv/wMln0L+yNaABeXVDe
YA7wj4MDIGMjf8y0pprsb2LOhUuJsjCz7ICpamQGz6bqT+ZRLxKOne8crWaw9kwi
vq1ao37AW5U7ijfeCaR+NDVkm5BX6ldhkxcp9Tu8INVhiBs9LlKx/3xcHr46XzpL
Qeruuq8NJkDIJ3E+PUyeXjkrVY/w8KROH0/PHR/H6Dm81WkA4DrPiJjsLinjOo+E
inlbi/dLXYvuTEyc1hmCCITrZSndnbHT1kS30mZAPY7TlTvU5AAltNRhm2bZAArx
2tFWo+ZgJs2qRcIxWbB5uaskfE6+oCEqNlJtv3Y0LQIHLincUrDGR+Mgf9QkR0W2
gmfx6JuZg77YLuoxRtrQRVRMoXgYZCQ2eL5sd08cMxr1i9RAL/ZsDYvgSrG8iIUU
Lc+YuIJPfaOryZVSE3lm2byDytbJVGEthxxZWTJE65uMP3r3B0VednTPCIcs7+X3
T1L3tsyhQYU1nEKEcMKj2oaxYQpdRxaNm0geDUbTAW/e0dnn/qUlrwDGAfpOJMs8
zd43In2oCdnonz8GXTqkEW1c1seS0RDdpRZ9l5+6YT7dnqSaKZ1+LcNkWP2aQX4w
Aw2vcBQYklXBY086Zuy0mQWyZIiC6WhzuGctHS9lEHXQy3m2erooCRawbmTWXvYz
i/RvR1APqmYXcFwiQZgFtmhpuwao8NKytJHuRmEp2KI+V6CakPJ7b+YiQzh7ZZ1L
JnmWeU2ohK8j85dUMXpdcOS/nMwfBiq5DwgaumAgmNJWXUrwIZznhAizrZq/UwSw
Ue+fHTwz+CBBp21BN9N7FaW9LvLoE1ZYO1umBCoNkT9x/gF+F8H34Z5NrNMSWZ3D
kYcszKQ7iPPc8UQrW1koa2D246ZtVg5jvqIyzYEFukWjMbdnWi/gjOzcxHoyORZw
Xa6fSwtSL2nWU56JYq5yCGIK0nzHNCXWfJuPSsFlhAP77cvyLZ/AOc2J93+9xqPY
6BAEZLsmajiynN1HHhFtcvfncrTjvsyQG7Z2tQ6MEhFKs/nFOttrO1icOTohx+l9
m+R9GNt+p1TEx+iaKfgJ7iK7nmpMa35m+wp3ObfXv95RJB5XOOlpGPCDU7O7tGjo
mVd6yVk2BzdNiWPlEjGHS6GXKQ7gfkm0pVQ+3Hs1Al6FhFrEXLjb4TupDp1DXiVM
PA1CdINrrYNYI5kWxWhJlzxSAgvVV+ZY6ZKDy4VdfUErV8YtvnkQJLJi0u4q8el9
+CF/njHGykZ+WmXOzc8Sn0r5KxPUQlm4vOTTgEyaqQkrpxxwAZXB2LwNRLhwXVDO
zpwtBlGRmCT53y8DViJYL8ooOYEqI2rWIpHSzMcJ0QaNgN8Bi2Yl2VxvBqb2Wm3S
odsNdsenSe3coZshRvenQ+jySwvmCNwnCy/RTL3x0btQbQUCLf9vhPE4xSx+hKxh
lIj0OVvTV7NFOgdvbwSClMebfvFhQkHpsvWt3QeZL5dEd7y8pntnQAm+/dZdewCS
SKdCa524Mm2EzBUUNqMrfibJWk8APiLmgnFQlr1a8Wl2ZUfbCaiEeG8Du1tthSc8
Lma16TbwlycRbN6L8DQV/ByVJM8MV7kZsmIgPsHSK2wiSBRZxH2xiqKFCAjugfUp
0LXPCJmlqIQTq+qzTyQwHk/3BwVLsAV7kyyB8KIJEwTu2gROpV3felsJtLIYVOIZ
FjO/BCBrit5yMjnVMoRo236JRjCNTt7OL5yrkX7WigYf2A1Ic/vGtq7zhGN51FaC
ZdwX7kLv5Y040q9WsVQ1xW8UiR63wurMCbTMAEIb3ytIDqumP0IQl5D1Gstq/8aN
FQskxfzcbcZEwhqS5wFABw1TC8H5Yza4ZqsG1q9VHCwkRTS3ah+ziNFx9H2k9iYL
KpbNQN1jAyJ3sWNcl8T83z4MhbUMjjNlOK9gv8QwtWyq2RV6dCw/4USyyMxybzw/
Z+VIePeLZIcDKxZ81U0w4GSDIMSNwW62h0to18stDzhEbrjD9Y9d0Dxtx22S3KkU
Hqt4o83yFrDbZOsv+kdKSh12byMYhtrwmuZ0Bw9aRTb8lbLPdcCTy2tonoE74fIL
mhspk85Gu+nrHVZY4vn93QgUBsmeMK4WSyTG3gcKHxWoMTOjc0JkMGa18wY8SjME
HQdqOTz1WAOmW3TghnkW89F6Fuvnw9B6lt6JwvEO9ncBu7Jp5xECrX5KJgwF4LPE
E7NknEJdKio1lyO7hmN/Kx+NW2rtw/AUb2x3Frsc/cRMBwYliU3AbtjVCORDjsQK
SWdlXaqDKlJ13YyQV0lkPr76lABU8sCvg9TUqVhs5vyf9T4eXDUGG1c7btPsr8BC
nhV+wnAI0wTrBZptSeALulGs6+Uc0RltRqlvis7I4FtWgnfi61fp1hw60jmzSaI5
gpzodwIr/xa1CyVS6ss6yspeQTD9+5XgB6UyQbfUNyjRKO09B03x+QBoVsR6ozJQ
8DUAmqHvZaRP7IoFf2S9HuO8cMzBndQCWtzLHviyGMqLJgGIT3aexXX75IexzshB
sivvU8RIrzsENc3EIgms4EhLsFiupHXZZkVEXyGRaeAdN+/TLiON+U1Gq+QRyBzc
y+p+fkg+Enbv1t86Msb1CaYw4d1Atu/3C+KUcEiKFsbz9XSH7iO7goTmCgfyLi17
LdACxqDfIM2F4QGKT10PaEHX0HhGdmaXethlIGTTtWsCAPeS7/xEXOyGfosCx9OR
8Qwh/uCSErySpbooMuo080k9w90F4uDD8si2KVjexGatkYNEEoisUiqTYKSI85WL
rSF0jO6orKys+nL4dm4DEyJkVqXYcBAGB9JPNG6GmPfCbIVh6OTjuVAJPoYYOYwt
C6obGIZvS+KarILmsZarYKoRChaVvQjyFJhZyxQ0XCwYl/sWYqkmV14Cc9DDLMn1
vckk0qgelYmAO0/d+GVreN67Hg/7mNiJbs31XDeWoKShr2HaWhAyLIX5oLufyW/X
fBF0Rp5UkAAH2J5Jw/GcZdxcSBuhn8sLgVV+w9i80JQ64DLPtSz39tCjimrdew1u
3g7CiMAWtIvdDZtcgjZlc1RZ9tRscyscW2SwTko8EGj7irv2CB2JDpqnvvlo2wrP
H9Pii+4uRZrIlK0MaLkwHO9+egNcZ6yIulOfvS2WDyRoGuvvJeUHnWPzPbeGqWn9
fGS5efJiuDvNvLW5nPPgoTOsoAwFSnbvMXuSbSOahG+L5vW+/KhEs6hWb7Z9v5c9
hkTJz/uKS2vWvJIcFV7O82i4ZfZYidlnPXovRsQFJ0lGMhxo7USjEaIsP7UO0jpK
GYDZPFDh+t/RU4SwgiA96J3r4yzY0XoJnBjsh6grunyP6Z+aE3c8xmWf9hJWxwpr
27utI3Qv/KE3oSKGIC86swweKpZgvc31/EOD+z/20HjUN9qZhr9OEm3hX3NwRPef
CsSDJ0KDug9pKo58SuoEhLIeoaOarVUddpZKmWlv0xP2cMOWC5sgWg0HymOZ8hO/
PfzntTlYDhNpejWmtea2oHxJP9NhMcIDcOFG82n+BQS3uEUpmQvYKxNYUD5oAF3K
ffmAXoQbLjGjh5AT0j2ldXzd5TOSRwKM+/9aZsVd1oFyTUNBR7W00LbCIbJapBta
wXpXiWjCZtdxLRHKDSiAVT1ouqTndldhrzeny98KAJPAFxW4lJ113ydN+c5VqN89
gOGANoU35MEKtNu3vxhnLqHPHYsnD8TjetorlHJLqCJgVA76gmTIlizLBFVn/vGl
zqCQLNuFFUgxDlst+2OBtRNk5kQcbMWsQFaEwhfuktdbZJoVnGDu4Eht8A0YW+oD
HgtkYiDYXOH+dAZzNA+km/OJgj+AW8mX16J6Q4+cgirGTXLnO3u2Nt3yXMM5Zol2
kudFrLgTItubofOjjhRhxdaelTNmXq4vniTBr/RjFEkaMUkXDGk6rPtK+69FBhnk
oOcgFWwSp9xsrRQ4OHN+DMTIX2Dd1n7uFHq1WPjLMAIPVWJikHtFRGlar9RV7GZf
XV62VVgk0AQEMjd3zdVodQNTbY/wlSG4BY+D+n+vfOFkiL2U0aWgPgXEl6egYLF6
q9gzoj1rHeBWOYxwdC9WlEYmM9jAARNCz5/w73tRcNsdCCGIPfKYeN3nH8x809k6
xZSC5Es+gjcpdNWeU5FjCe64c3NlENT4FfR2BnGjidLPxF4yzRNcgtFTU4Awj29C
GYQuKmVY9MozyTet2836WVahRrnevWtPYdGBRFKF9a31lYSt5oTaJUuNcWpHYn49
9rpLWjf5OTyYwNNliwDUK1VDXQLNzZe/ZjaXAamtgMoh5BAblVGeuiCcihHWO37P
YWCTgUy+O3teSRwFnEhfsTeIWwQNUZj86bcavLXVKfife7DVL9KU8q3rYOROj7Vc
mdeFedcg39NJRxKPabXTU+GiV1se7E2kcv9wOGNzpjkf63a1UQMq12IprZwg1h7u
KyUP/9PDewYo3mg/0P2/B6y7ZSnIy5Cj3KUL39D2xXVs5HQRMi7T0uGENvfFHHQn
o5cNIHG12wYtLCdvqJy3o0R+KpdGfCNRGjWHapbmJck1i8OeoddOaylWaaE7pNw8
sSjxtLBxiLmh8fgxR7eUEWIxJdAe4UKJYmNxdN5L6vZLLMXuOutGh52phqRTPHEB
tZPNnj7SkDyjMwOPkDJzvZQbzOVbAUh2/a9G5mCL4MUszpgmUsnr9hif7h//TZtr
11boq0ZLejx7r6tO+bKbyuF7TukyFxLzakkKe1Pj4vmJKGmBcSTnrOeo1UOgGNys
9kKivTj4ysTRr29U4QZtF3br714J9amYW0T5P0M2SBAbaEYZYhAUMC2VveR5brJK
ygj0IYriUacgZm7QCCzV0EuKfUb9UO/TSZ9uX7BtbC3y6Eu2IxXP1sZkxZ5DrRe5
E5nkdFz41l18LyvOPyRfZ1aIk1SxykO6x+5fYibeuanrwTLkAif0GQ/ujyu9WtCC
JrcaZQF10iNFRGd8iWyg2C6fG80420GC5n7/0q7cBCGHAs9XugPDd6wl72pIJlch
eeEln01yR1JYRxAXX+KiZtj5T0qma5WV+z4XYjgU/UtEDBChhJJqtF5WNeEqQhU/
OgmhHxEymmxM4FPYbLhcjsGMlSfb2Lot+vIME5Wz1i1mf14WaRJMN/Q76g0Ma/SY
7ld4qcpQqM5Y/31i6kuOhkxAZziefqydQyBayukKdHFl5ElHybd+dIWY8gVVFEEo
Y/lF1mfF634x3WJMGj0LQ73yhVDE1pblK8408DTkWthQs9OOKuaoAdQUp0xtjg0n
ZUYTvqJ5FNEx7KW4L0GtmPjExtxy+1uO2UCJ7egJUl/jZUgIpyBMq19J+0/dltwl
Wrrj+pUFaKkv2rsVSCSRFovru+0ALOSFEF0BopMKtggg1sXx90yxrQ9EnDX2leIV
KzMygv3cLsHNeq7n5Ng/BPlL2BDXajUPa8nGMXKgZyt5DsoAmp1YHcZaNkh7fkO1
jSzaLHs2yzbY3UIanzpuzi81OzerlpLtAOepsaIiATBCAe60bJlVTnrprsLTA7wR
uwaMc14w2IPtVa1gTQQi/QfUvNhHzRh09K+EjPdsedRs6yfNfhaRntVTX9pjUJjR
vrrnXokEBdSw9lVT590y28orl8xGrjeaSQyiB3VUv9mqxDnHYAfnQpEmbu0fMxCN
GxrIktHzmGMoZDUh0dd/ThewB3IxWqmmhraEeZCXKq267zCrzG187gzCbNwPqbF7
BbLpEH8+9058nRSgBUWUuDWP+KxagPE/TcaWVASz6og+HCub2d8GkOE3KbFbYUoP
q8uxGJzBaiobybKExYPztDcEUHZFWxc5l9rR3L0NRieTCCYlG2P404tfHPLwJnyR
YuYD3oK5by7yxhsJs0kOHDfqWhs9W7JX7Ee8BspBsP3uykaeNzZOatKL9u5R9W1t
HzTY+HkV8OKP2MQCcx0WkavuKcI5WPS2Uk9SoqxT1DWiTDnq1oLcpTmlzXxinQr+
j9gBnKnPI4/RcLJDkv37Q1e7LXaVbOVTlZXs8XD8RaaVpGKVNPpiV+OO22o4Ny9v
qSNc8PtQfFEYG4yDQKSOtUgZMmKqU0kmr21ER7Pm3wiJz7qww/a4sN4AnkDsbEPb
Eca4qs2lcdjq1UD0DNQk8rEy6Ux1whcMqsr9KtafBD5mZ5bSDJOtz/G2LGniafu2
dlVdM9u5Nk5+QS8SSl768uf6QIA3tST7uv39oJ8j8wWq+9Pjo+ozn70JZQi3LJLd
xDhpYUx57EKRlK7xTFxt2GkP+OCIbVGK55GWdpFimyVckQkzemgUEfoXrfu2887+
mobBYMl/hwRK7xtpnEbMxmrwG1nAJedaxpVsFpUQXC1K5hGugDLArzq+4jjrdDGe
mBcF7xR/dXLAl/u2FuUngbHOgzv/v6/ahJCSrkqIzZOyhHsAORbsvvcqjKR2SpUC
8TwAmTiJ+0kG9qZJn0F8olo1dmEHOi+0UHZk8ONr5jGegDbfS30eM9qqiSKGSkxS
gxTMgMC24UqQbSfS3q6YlFLGldzYeSatwLQu/To7Pl52yln/IIpGiuAgLnttA+vd
dslbYMyzKOx/7H0EDMuSw72u9HyhaajGn+BL9oedlKDOLcg+nZ9xCPGFzrQJhWDU
Kva9+BeiXM0EBYOIIsP0X3UFWuyGJ2aNNssU6sjc2THgWBODsEsuX3xEomhDhT18
4Qs/Y4raH4LY0i/E7vbSLlxXLuBK+BTz6HLRdAR1+ILvMKcYL6BERSIM9wf1rAYE
DdOMmVbMR1WdoKZJFFTD4GNSPLDwZicVGcZPZ5yk3Z0JnAMB7//vRSqvKXv3b3I6
HXyoIpDSZ8kKMGEnPCNEUKe1y2FzzX8AdHsztwkH2/Im1wNmVlAff2Nksfw6eRqG
UVJKLxwtJHxOHYNZzDNxUnxYzInuEpmv72HfUcwIMF2HZVaGX2z4fv8CLZoreUqi
Peg9SvEuTEZNfXVF6R+FbSyjiKoRkCPWK90vAGPHBeafCWWnUyoxDvHugwVyVdR6
MT8hOELmxqK8/fdlc38rG7ozJwYBUjLD376yCZF3xaa70SR2fDc/p9p6JUq3XEns
7q9EBP+jcHYAMlZmwRmkb2QNUv0Jfj7C2GcDpZbisPvcwFrzhBpQQjisFuRb+S7J
Pzy0Ec82ubCmgdIS7vPawYruDQlv74qwcawyrGjH6hh3lSaMYaNDNQ2L/gG+X9BX
//ubcEquw05nb2g2i6nOKWT+WLHUFol/rQlkpAuvZYUE4OfP4rjW6W/Eot7BQNMs
cEhOfaniwH2MDaNOP0Cu4HmguI8YhIbLoIipwkLBSP7NSGfhYHz5n1EcwR8/W/XZ
Q/xZbvTU/HNP0BzmgkO/2QJZi8g+q+XUwjrKGAeT1epE90o2Fr4RUoPXXkniiupq
p0yiNdGoygLcYwfbGDsMnedEkuoLQ/9QIozaHbCIWKrlA2ijekdn/vVDBzEkTwTK
OsS/896sZvq3mOrquzRf6VDM6z/TRVJnP8X5bkJMT/gwJlNiM0MTbC0yidWXBJSD
Pzf1IwcHOTnn2xS95nM0cNOw6hA1KH9zMWT+6TbO3guvuEzIKhubfF03MwlEXt0C
m5/SJCxCvxbJXSLAMpKVRdn5JoNizGlBA7lfXejKpksFvUfXQ4sOJ09a0LFydV2D
WEF9/x9WR8CJWhNtxWq0hyQ4Rgs0Ro86ZQRmTFGrVNAtilkPRQ0QU693oKyllx7n
Et2V7i9+W2TFvU63r1TY/O/cZhaOQ7ljEc8NT6j8qDklF1UMOf7h0V2y338a8myA
o4PaOSiS8hJFfovfJek7Rjpx1UnuqlR+iF0i4UOzIQN9VOHwQTYlhqe9gYzBuJ/p
k0zcIE/gPQvWp+RkMviy4oWVfhzuslgAtI/1jq4wGYy+1JTGQ889YryqZ3SehH/X
QdbxfSg4CSyrPlm0Taybp5Le0dbUImTmeYXg68LNP+gRhgJNYNfjYf/LSQ4sWZ26
RrJQRqgzMcR7kJPmJjaMQzQFYHJvyX+ckMgBtJdAic8Mn9KEwxsRiFI84RmksVy7
t8BsHgB8ILmRROZDbF1oy359+wfgUXkpwk2Etu23s9HtFQRaLTFzgVW2IYG7L9GK
blaLi41ElgltMwPkVF2bPQN9vhUidxrvnbvtEy3Te1IudOzN9w0RipmJl6EQpaRh
I5o11Y/QoY/8PtChzJeUmq68TDHzLeKdgwdnLHJlMgNoBoI+oOLAmF+vt3wRM5z2
T4YbS7CiqgN1sCpxYmxqsB4GI+wrsw5euWYGtfwXy2Gc05SO7v0mXXlEJqrLnYY5
zX2ZQjBOD7Xh93532TAH1f8bPzfy66gfQlRmR/jBSsf6MnVJIUnKnveNkF12/nHv
iFFOOZR78/vsUhLN81Q49cey9IOvee72x7gPA2ddlkHpBtddYAAII4s+DpasQwk9
KfImv2wsyQQ3IhD4LZ+RexIjNM24I5kSXQe+vJOiRmqbdMYFnNLzMbI9Dpr7T1rM
4Q3vfYcZDrzFA7+vnNVlk72hOR+L6lqKSzjdEEulMhZz6YYDL7p1ycKDriaL2HaM
pgMRFUCDyzsV7ItSNE2Ysn+nwyyzt4Agjfup3hUQUyyc0d4o24GUmJO8/GmWajqW
6ip0xXNcxP8U1aRszGlgcTg/tnZa+1ZFxw5xPbsdJxPDNOn7W/lZ8fxRdNrFDGsn
GP3UUcgFym+1n6TH8YzbAEu4K5tFWg+R22eT36BQjcASDPI6F/bje9CNHkAgN6+j
DTKVLnKwch8KRGHO+ExVaMIo/m5hRoL4oueY38YVQjbBI+9VEZ8RGd3P0zwJ59gT
GnJWe+PirkymhUNOjVzXWhs0084m8YEmtDURsn0vFAC4CxhE+mlsXNslx0KxVOKj
YFc1kmuMl4kq8tWlT8/iZl5r63/i27WVeRAxXRdzm6dnNbu4f+uYm4HVyXQyRNHY
oSQB4BtHG9wST3RfQZUl6hktau6CoeWENycDjQFaJJbSZRBqFnPIUJ/o2Hte0Pm2
wsm/uS9siEjG1QP3O8UhuGGVRSvJqbiIw9Vo0KSIu9Gavb1NvDZTm0FcElXrbm6s
vmN1uKR7wCY0HHJcHy1O0otoK/WQ1LEOe2ssBkpUIh+xY4VatRMrd66FUq5Chmfl
tr/K35ZJ4Y1QhYrwyLnIYPb1t4rwDCErW0zPoeGv2ahQ3KdOQFE6W+OQbMg8xyQh
PUXL+mvYvI4bx9IkyxAbMPX/iA6cj7OE/sBypWo7mO7UqdMy4LYzsd6mjy6qx3YS
pHCa7XFLh9US+gYe5DudV4jnsLwhvQ1W+cUcgE1G1rC9qx8AtSkx6UAJwyRmQNtB
KGb+MnfgB8ptFQ4pxonQHdbcG4ulOtFb62NoJiphDI+vQzHgU3SB7LFOJXXH66pm
YL2iNCcGk5rGOmrMsqqUhDvadWzEYB7OCZHEAaRJTE7D96GceE7/n/Bzu+qKdd/m
kf2j9IVf3OfgNcLzz/yHHSVZy/AnBeIY8t2kidxtDiTR1j2UYb6eSeBx2iUG6xE2
W+qV8ZZxZy4k6ryLd7lqe5SXoMIY2czJPN7MuaGTJKNsqBBJN+KUlkUNzfryq4CA
8LwRfjlz5JP3VkgAeGKu4GVDMpbD+hcknqjlFT6xA5KcxnR+2FbZ/ywjzBCVBmWD
V7ZmXI2zFH8oubiy/xUW98N4nQF+6ZK2wFGfzEo46YICR+pX2rQR9e5RFs2mescC
5V805LLGwRNQQnM69wzO5eSGOGqhVILppMbbaiR3SubctezkqMWMpewm8sK3pIvQ
1p1dqnv2S1rBADxyIJsFzd9lOq9TDrL4HTpklL7KmMOZxbk9CqU8UjlpWQZ3EwiS
8VLKRlCuLZJKGBRWxqmqTSUZ4RMeUISOF9s1zXF4mCcaNBEvshSC6z+ZqCQM8Y5m
QcDSck4xd+u9/5nvQhsm2Ln5tZHn0NkFfnVrZVtiz0hpoTgg5VLF5yUnicd+Qdjp
tGbzaxBxyrBOLK2ur51Wof50Au3G0HL8ivq/XOwv30fDTL3wjW89hnOrisVQuWE5
tQ+hIc5+RoQconF9BP8h0Tm+X2xKwItzEQEndiXUq9tJV7R4p+fXrbAvJ3NElBpg
bIPPFHNrNOdPw7yUH32PX2GGFuIvkg1XPyY7a1FaKkBSGUkA7zpzr9hOVriXhMw/
0NPTrBHx+YXwJ5zlaeS8hZT3POYTAF827RoA2q2sFj3dcHmNcSYjKUSoprlmE0pr
R0dAS4HZ0OWO3KdX1c1m5QEU/3srg/az4Wkv03agpiqmeW//7chyhpoQpinWqqi5
tF/PEWqpB6QeiH2iNZURkcnGGVHJtSfLrs1myin/xOA07NQWrN6MszeF1UHmPJ5S
hteDaji7ped4nAzeE11x80RxFbFrOwwbD67IKSTa5YNbPcqAITjWI6xFVr72Rw2V
JS+BBgytVJEZj0Jxcx9FV3GamMlAtG+7mWppuqtgaSkjbc1FIihqvVHnEYZcajkf
1P81U/5xAuxmb6CvJrDjY7iKbamR+Dr7bddEamnBPydQR6ju5xeXv22ihSeJ5SoX
DS49DdrNs11FgTWwIGzg4ORhmEaMx1R1+EPwW1DRInt/q+/LRrWPUQ6XcXbwiybP
z/obN8efHw2LUdVz9YckJ4g7Xo0JKDHQ9BVk/OoxgnrbngLYor/5LCgzsOHO6RMc
xBrqnVLwBvDgwGJSTpox5DqpFM+KqZLPuuvOtKFZ2evm91/w6Pg0nMgtM/5gSM2T
m8TsJRrmSMATyOfo4cy3OM7B8PwyRP08lNmTBodQUoEPzRahlTr5P9lvmSgHfpLo
aNtIMP2nGiuLNSotAD7a6txYemsMdk7MTeJ+gxx4UjAytvSwxI2sNsLSCn0kC9c1
haVZOjMfKam4SDGgDdSLCKQ74YQmQ70DftJSi5KzUhwMhU+oRVDfmKJa/ZZjI1E4
r4QMoMCZBOGsyLj0BvAwvicAD9ekdnI1uuk4W2hxs6xeD5nVE1srSKIBQfjYUsQ0
gA9ja1r7ca5FSNm91Wu+snnOiCFDjlkjP2FasqOpPwdbQ2UOm0QZGIJMblHRPWBH
Bf+OLqRLtA2nxkxhrOh8T0/qA36Isq3FCvpN8AMz6XvOiHesY/t2AwZyVwnVPWur
3v6XOOWdx0lmHF9r6r4eUsPof3ixslGLNgo83Ww2cC1S+VhQKGkQCaHu4WRc5yew
QY1YPId+hRpRJauGW8O0aZJn2WuTG3MZSEHNuWBVuWKWE5h6CyuKhyoPQaTR0Gow
g3pMCfefMN1btdCa32CQyAXEEHSrGM0b6cgNad8+pVtIBGzJWXwsfdHXrhcRV5t7
/2yZ0fhUMkpUHklBwO/bVLmcanU8/iO1wFR5RIHjVxx/w+C5XqnVB4W+diel4eSo
z5a+QXkqvTjnNld1RMgXHkFEEsmVogWOO1xoHnHdnfMlZuA3sbZjB/5rnH5+6iDm
q9n9660RIG5gkvd3mR94ypbXQiC6wXyabCuSroqGCVPG+f4z45pYulX+La8/MMOW
Cjz45Hkd7a6c6LWUG+LILDlwASByr0zAlzzDRvM5xWVYIuG4aLWyemXFb0JGSDOp
3+Mz1u6LD4P5QQdeD9wiOEGNefWlaMNzy/O8yCoIBABjkQwFy9hy6g7l3dnQEUse
/66LJMrL2fnVnTZToWf8dP9jEVNhpKGPGCVNj60wXfuQtNBVLIoA7u8hFYYdFCV7
frYsAFguKknLZcg9vSGxFTVwl6MwUI1Kq7L0UACGkITCHSUeRawZay3TjFKGNzq0
h2zFJi6FUOuiPREZDF3cOBxOgZiV2U07xx2+2n8GXpSTLaBAldIgZjz5tdTf3EpH
92uxcD/oMrT91Km82NiXIAVpCeVf6uTwVplw2Y04KPAkEdrSxGot3PuPftkyn6ca
j/Pj+nWcWRE+9ssM4+ekf47msoYHIBothGcqOJbzUfVQcOGi6RC5lnEnOvPMQHTN
7IxwCgAOeJm8IKXpHMxTPbnXpjGE0KW2F3Bx5/ZKk7+V8AbpyiWyYTugc59MjNd8
gsb15wnGX1YtlYPtOBHSXBaPSyH4VQ9LtDcf2ZakM5t9qZBMktMCrpZTuLAExA38
xuoUdYb9vKNuXCh1oynjQBB2D/RWXzHJ5ArX+lp9w3kYvVfeL+KDG/2v/e+TJjsa
68NJ2ze2jsV7suk7NZ1iNHhafAK7JlGcymFE07AMAMbl+DPiyLupgyEETU0Ax+Dd
7EIZ+aVAvJUsgcq/PyhiQy1pkZ/RhxU15mDBjLDFQPgEuj9hUTKRCocpwF4+IFwW
SM8VmGfYjT3jCqlEdMDqed9GM6ABJftMNkNFVLSzdBwzjabRCZBIvlaCj8MV5nTL
cxXE6OAiNpabQwSJjkQxfWqH+psJkustovtCftH8Q1vO2Z42/+MLcaj0JQwqbvEQ
aY0RpDU1in8Qyl+KYds0faCPj6msKUl5gr4Wz1GVypxsvKicYCs0VRNndeOxsKer
ggYS+HkAuAv9QLITu/VAV6iCLey/YdPaFy6d5AEOi54rAbWWr7C/ff/DzbA7FssV
iD4Z66+kTKCNsAwws/KOfPZ4uaer4xdzaAZxjXyGTICaSNalw+ah1ckHephJALMD
trv/o7lzrImcn4Ckiv/ZleMLevWcn8BU7yOoAW5EosTfuZPzqRQQ0wFuYRzY1Ed3
HFn/XsaQgrXg+wf/d1u+Az4p1jcuBBV6dqs/yl156/3yYBdTGqUSBbdrAdCbul7f
/EXJhpsdDCgwwIfvx8EJ0q6ScM3BLXqooiulaQwPuDY79LKuJhjqBrfRJt1I+VE+
wSXJpwW2DvrsGyiA5aLuoW5Sj5+ZD5ZBLD7kk3DH3HZg6ghxwSshUSO5EufJuhDX
qF4a/BGuuivxIoWZwxvpG/AnVm5rAN47ySOmMP6xa3KuOZIv76ajNly8c94sOscZ
Rhy8OoiuF3XBmET6dvrOSuS/cKNizZjL4MGBenSxUz/oyM+5SvrHL61L0hAUeHIg
3jLybccIw4Jm5Pr4Xqb7ZiahLbCL8nxThjTiuBKxnsgpBTZl04vEiPFb/CTP2dM3
A+GpkJSaCthk8WF/vTpkmhOSN/b6rV70ebHuszARSOaashdFL+yDWBPGM9sSvTNG
grWzYkaXlF7/vMEVd2G7JU9HpgadWndOOWie5T9QR7hQFzCv0jHP0UN3JmhrM64k
Be5RN/msFi3YQgmwrheT3Pb4l8DUpDEWxt47RiwP6nmper7bXdVV3ca2L4TwimCo
0PQL+P6OqxJCZvhowU2wuYFg9l77XH6L/BaVGqg8OBeywFTkJGgrjWFutNcxk7wh
hiI9mapTZoKf2zJ+HenuGERE5ia6xHIe5YfmyiAntynU2xAsjyJdLaB1mEknd9ri
UkHLXS+yOSGYRgXOnxQXnM08LcyHP7vXvu/6ChjP/fdecmWMbFoEsgT1qw3TLUmJ
g3B1iQSt1DUeaOp3yJ+CyoETrV31UBAffTxicqDd3exV6WK0yweFEUm0TWGlNpZY
YdWdgPGly3YUy19AmT0tLCBb4Us1BWBAOx4q8Rv7d6PK2PosraFZEjQmZbk8qG7d
Dbkza0ocm0UtJfIVEmfSfCU8RAuNmdzqoqyrAirrIYM+b2J7N9Fmy5txVUNS9gXY
WFcuf7PJzOyKwIZ4BygUsPtuzptJY1W4Vupo+Ycrnec4DPwBkLW5n2Yr0zReUjcw
q/1U+UhVf149CqAnGNOyKYbJaMz2sU0G/4NyRkAWCRoJPMb7dkevoAxYpVl93mxL
CpWPA6854dK8KmG6HSoP3+rZH9l4CA0mEJKdVoRsh23Z1RCnWlZVCeB+fTKMfh4/
LSgKfBNpuqKX+/5UyB6jZmCN2Cn/ouoJSR0RT0ISzwP/MO6aTqPDn3eXzWoRIpRs
xTNNtvrNZ3KUmXw8jxZLfCIKaorPgHvuZTeJzuDwQhyRKu+DX9itl5HwNTdqcQA4
deOAShgAe0EmqukrFuJK0bMXkqhxH93uw7bNS1CZjTxf5jKomyqd9oYwXCUIxwnd
W9xbLfeOsU0hd7QPp2fzH52SRxJVkLLpA+K9cLDcfrM2bbVjiGUulCd0TaDr0i9M
XcZK/RA64NSEHkFYafm6wxOANV/3nNuaTGh/H3ClLOZvIWJU+SzGNZVB0qNdKgGe
auztNzm+woRIc6NicbhiXk62gKL+j0TdDPhucAcz5md3jUM8j3hnvX6fsjbs4yIF
KkyJa7BJxmUYNbVRQvtw6iGdfU+Sj2q++KD2IZd/OpkyX+1Cb0NC5swKVhZGl8/z
U2UE2oMYeCk7PTwt1hDzZZkwhUO6bKgHHviE2p9K47j+XJJyEq3w4V4fo11EVjVY
RnmfqJElqEQi3MJEYzIK9jsj6me5JJFIzEA6MexeD1IC54sH/rX+12IoZ/I2EnNq
fweKjxKJPiDHzfEojFJ1lw3HMS2ZA72JZxKzFj1MV/Yivy73CwDf5tatDfWGCDQj
z1lvA8rqrBjyRFuZFBvKDioV+OCRL44xI3MKS5wp5tRo/HF4rkRIex3GBOsXrB+z
QFnzn7fMcy/BwJE/fg5pzHNEJ096zQJ9iqPL5QuPTKjK6cPNTYnYa+AFqXmLufsd
PDdA5yz9vP0SAAZysyvq9XvXHZrKk7ipuFOIF42YczeaggQoF3LTy09Tn8PIZpLh
PY9eoDkF6q49daCDXurPdayGjCukG0ZZm8vCEPG/gtmCQ7qdkUst9snvFNAvdOdH
udO4wyzMJv0RN/FG/Yct38EmHcTG4Pozc8EsrmEg0YbMGgWp+arfTseZrQj50/Wt
MtYZV4SovninocxUG8qwtU+XKUlr28i2H1VXqaa1mXoptlNCgbDtX2yoO7zlmqwY
r9V8BxZuGlG9sO474ZEr9nbPtNOqS1qlqDY6iY7uqtfaGpg4oH6FmMhh6b7M+Xog
i25DUy3MsGIgNIegy5Q6nMUDOgK3ryvHIWjFsMR1s0X8ceU4CYI/8+poXVCkFNVn
LSJkyFBmncTKyzXcy+UYPIln16BbnLnCynj4/YAodgPhq85HTl9hSRK+5c1XifvA
ZfZV+9UF4BFXes4IrEzME6a1qpZtoUnzF0YyWB8Zczx8xspDaIGjF4ibIIuA/euS
nFvrsHSG75J0PfIdxqivNZxHqAzIiXuWTemsidh8bcXeaNXLPIuvRDs++tBL1XhK
P24ZUrlsEK6LIJvzTkORQOD5FOWD5Om4Sl9pPMAYc9qrQ6M3+1bXufUPYX28dRcf
VfGtYy2N7BfAf6WUK2mAYk06pF2awInTghRieUX9oYnmy3jrjmNP8Grkokpv535j
sFQGJd4f8vxWyE7NbeS4yrzSxEWBSF0v2Ygq8LZHhX1/cQeRkgVj27GCsoiY5qoZ
ze4Fkw7GX0O4RLg2AypzkQAg8S4g4pjRDViPcxbPTpyy4c4+ML2TARyOyIElPyzn
orduhPPIRdU7mY1pBMuJ2D+bLBsQdo2nzJ6pGVsLDs7lDsoSxOipv7BkBCjNfCR4
rCS3vJAO4mRn7LehNV9Xo8GR7d+0w4+2E9VDRJbxnHgEwoMp4jFNiPkMGjHdJ/jG
7yJo5pPGPgGiai+aJ6WF9klZb4RBMAwk5OrGJ+W6Cn/vmRAI7b0CWcBiVP3p4jx9
qT3SN4FDonOiKU6GLbxL/JCZAFDV9ewHoUln05BNyonkmiqtbbtGHBbaQlZ156vq
4ObxdRPlTrONyEqzWVnPlUp1T5OJ1yyDERgfLKMXbrRrHmBeDDzCRaoJaTMft3RD
XEEcpjA5Q7k5N4XSBScauqrlo8gZgf5jdJuGf8ADZWqLUj441J2hLI1dBMWAwXki
RisrMWgMDFyJat82oAIfASXZqOH1v9MyTxzGRuQ4bTskXRGKWmggKYX6leXbAXH4
oiNp7DWF8UWtzazxuOUaan2rWJmw1wc3op41fGlg4z3uM48YUp0DhKc5Qlmv244v
J6FzU9hNJco6yaIp7bGm7V5hXdl9S9WBbS0R42VNwgXSfO9zzz5VyZTFtDotN4Fq
N3ZTuHn6Ti8nw/ACofF4hbQn50ZUI5Jy6nEjpO1/yf2imOy27PvM34Ee/F7BID48
nSJLYty/HJipoEjdwgIcwqnprgfK44pFPFKx3IDEnVWJi9djdvmjAkQCg+HhIcxQ
xpefOsJYt9f/nyLJeo8FYL5iqcChwSr0DHyG1ARaNY8hVFHjZ1hvmPfRW00ahP8g
UKsMBC0tcw1NYnl69VpoTvwOhOqdlb2znRvPbPAyFwx+4Tyv/wgMMNSK93LzXE5h
hyyWtzfQPCM1bCNkx4r8r4/fV8AtRC2RTt74cL3k8dChHUVFk1cGyEcgeGmodHdL
nhjx9eFOT7EDN/QTC8J2w/E0AfpHaXxILY80P0pM2ocR6yulGjPF1JFRVnT8f9bz
WgT4gygUlc2rAqW1tgyUsa5/yKSJi1fxsqg7vga9fEWiGldWkH+cqDCE1gYAIyoQ
6GD9UGrqWe+LP1TdXZBpvTJCa+SV10w0+rrdVaXF0OwV5k5fCD4mVDk0wh8yiacs
vPj990S2rg7atn+d2EeN5USUOLRMyqQ0kVqj2JXCEeuxSDftwBAWLzh7u5sdP9uk
e9Gsy4EvifB3QJU7md97cMmM/JQ1h3xgOX3BSsnFXTiJLnnq/zr6xRAzDDGBstuN
gYEij39gr/Mh/49S/8Sko9NSeWZ6ZoIOxyCPUAXH1TvbQayTWmXpDzTbwda++U3W
0Ni/CTOElz2Rs12nByhQu1mvphseCLNk4xo2EqX7HqkrJzFl5c37cCwwaPwqNO7m
AzUHS1wfCC7Ze1nUiSkBcRVGxWaE78IBIImgTLLaT5TRGsu+QWvsWvzpqUOpc4wX
JCE7Vib/nA2qwwe4CtGLB+D/wKxaVZjoUekBeWF0RrA1ETgAUHyVaKYT2B/K3ndY
KHHURyNOkI4v35B8/iYdi9N3me7fsrYb5jTVM+7YSEqM7s53WeCXfNmjQJ6GrLMT
BdevGn3rfWm05ol4KW/MhF15w/X8Dj3L//wfDjIuhdZmTeNHocGvb88WxI0A3EXY
JiqgqXiUR3RX1dNwjnlHfguoyI7L1kdoLgTmyVJhVw/IYNarEnwpSldE42bIRWby
ZDuTF8v2uEUYyd8T8mbGNtRZ9Aohf5eVU93zBXyXVjQ2+F6xkuwbQokAnHc+iwPn
5cAuynior4jwTtuN2a+ziF0Q572dPIY+XiVRD7afLNGZhHMq/W7imQkEd3cNwYhN
42k29nZViR1lqbLiMNmO5ecW/OrWZve4ml2e4AHYZGW9i3lsQfptChs8/qqnXPYh
kfnl1GzNhYx0viXB/pDQbWrKYIlDtPOXCowC6SVWLQ56OttGA9AKLwlCgnDoPK80
b8aqBA1f+JCHreP0JUEqJYqJVy88WYQfB6Ai0wzF7cwrg5lUfA7v24VgXaxTJ0gW
LYV65b1qrOar2qjjSDsxB8n3kii2hxiV0xyqu3GP2oBaXiH3XTt5k0nsBUB7dbuy
D9T+RqESBHcj9k023LvkXaokkiLlw1FsnlyiTyXdYHx/kGcsytI3bn5pPfwsy2j0
A8jHef44ZrBZk3xB9y10HRprz/t3OBT94hwMze5nSLHe6MMna/+tGmEkUJW+GFnn
`pragma protect end_protected
