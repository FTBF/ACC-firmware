// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:24 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fGNTo9p9R2j5kWvvRS8cCNfbVY7i0yaN8xngvHEV61dcvFVVKXzpp8Y8ZGOjuF49
jGaGTzRWhj9hu+mDIuQUGoNN4X/PK0b7NfTT+ic3NgtVeEVDmcRQcUtud74zSSGR
R0hzNxbKJLD26mmORHJ4cZ/4DSBRXAwoNcE4YCLN6+c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21904)
GNcu79Z7ZTuoRNdfVxTSp+IsQa8x4az4rf+mWA7tnTAl9Y1sM6V7aQMy6lBKE7qj
dHjfogqL7k1oqbIjy7eRtLkkEBP3xPrGdDR1Y3e9JTh4tL2hygg7YFUrf6kyZ5zF
TQ+w762HU03IgbfQpBuhWNYxIyVMpyZPz3iNXaMuh3NIltnO37zoaNlFSxfH/9Be
W+1aYj+YC17VDJ+mtjReM5ips1amsLQ2ytnP/plsm9pkNWTK3uX1NMvyWsg9Ip10
jyCH3/opz+PqbmP2NLxpk2IT2JFL85uRcdQOWXpOe5iFT56FXsQ3n7Ofo7j6hEhr
ZSbgZlwBa6ZpBCzrtIzifp3754qPhxfImR2OxRoVGsy4BIfBBlXHr3FBuoiTgcKv
Pt9LMK9o+SAHKYrjvkw0gGIzXeAiFLecKPzALcsy0iLPr14js9hds3pCv1UVLmos
c9gAPr8gMeouxRenMXB8SBmUxbpYe7/AJ25ZjMknE1FO/Msiz1WzoN6i4Y3zOh5P
wJlNOAN1oppDATIGwSptG2aN3FTQ7NkDyFeZBBpBBg7N540Klx8O+z2qSMu0cDgR
QE8CYRHv2JhZHGFnZ55e2u37pCndEmzldtzcVWjBzRpl6EaJnBNztd0mjoJ97Sr+
jbzqk47g1tQsN8W9aY/iu+bTOd0q8A3QIoN6hKLZ20uF7NBHCWV836zJRH3ivAB3
GvAEDACP6JTBl9tVAf5Wt26VEOsRlGHz5VINOA94+qoKZeRhXXGRABP5U+bb7ac4
RprP4KKeX5Pde/H9r+vQw+ZeC4s3QmH/0+HtTrgfWhRw+2IfA94ohyyNMj8qj33l
3HT9j1BCVRhkmmUcnr8CnCJuAS8/sPadgw3GeUcI3K9DyHFMirGTsgLtiVhcwJr9
uMhA9KJt6vKgFKoW2P7z73BLbH7nzQYq5GxhSaLhzJqOjp4DAU8Pa6hd2uS+51t6
xY5vRWDpTEBtXMK6cB2XVkqv+m5QIAd8hmYvBqlXznw3u9Zzbjj1WeoF2In5zfma
ZoGnFSW5+McssrvJ0t6/GZcTEk6B9nGxlU+BilKuZajZJhSwqIERr+/pH+QNe5Mw
YkRECkqsxrWsTvpHf5xE7fDch0bjzu1Go879EThLmfPeV+SZFC175SX5+p1+Jks/
td4VvrUAt3SKd2wAfhBoJslMpbWcbWT5MnCzzDujyhCBLvwPrGCBW5zcGhopOX7j
X3NjP0+Pg6s+j/j28plGR5itRc+Upna1JUWjPwJvSYSv5IlwAVbj3Z76SXffR8lG
a7YDDOJA4A8Qbvsa8ZQvUgwTVTPzz3fV63xNDL/Ufil85cxqLg4e9hW3Kulm0fOY
FQsSqezlglw4J04+LBWd02eVqxvL136P85qQbtYl5/+bKBOJ4An4KLHdf7ZvuULI
riwzuCCMSPSBZ65J4vxO9qGH8vlywO/eJxH8Eqqe75bhwYGN7HTWMv0TZTPOFHLM
taoP2C3r+jg+tvGLtPlb+ohFbFTiB8gXF4xrRiZPS1/bVXYeyhn+2HVLHQu7Rn2e
cIBWN8TAwFpDRBunte6xZFDTjXanpwh2et80Yi4GFpQamdOjfZrSKxKJxJdd3Wv1
snen4jfcK6eEF5Erx1XgP7ztrbBpwjTvnBl8N/dnopu+/oyPp7gUxhqLKJ58glrZ
JtWM5ajfTdvph6++UfMct5j+e8qOvybKqRJEgzQ68KcjjZ4Qp1loHX3kfmtLkqJW
cjjTogPfCpr3vSAJLlz6fR10RuG1L7KUdQnar5tSN5Feu8+javltM5kUW7Lc8Ye8
HV5jdObvWuzriGUnsD74gPerE+Bbwr6By93L4ZQT21+74WlGiPc0kvbj5hB6Uc6T
hAlu422sNPTxzwLYB6GPTgd4ygt215uGgrWDR0oyBjGihcp97I91v4vIZgHdqj/M
XpK2FOTrcDVczKJFYwpCFi24Pt8A+PZ/W5JUJSr/EOSdUJMmItPbAEgYsMJNH9AM
mCCGkoBUNX5Ghi4hjoGQsYoBvUky86UnIFa+l5FxnLdY0yLB2N+R9LXlIPE9vRFs
FRv/RLeq6yQ1pK2mh6hpxAW97lLMr9vxa6qfKfjy1X6UOY480/FsR1F+2spp19VP
hlfg/W6Rv41sxX+7V+xB1P4k33vq/UuOShbV952aLDDaq7X2CNc5GyW8sLjuSMIl
4u1Kn0bxRTtLy0vr1QReVjKKBIEqLZC7Rqv5LIrbSpNdo/8o8+FgfigZmLDCEn5I
A4u1+el4F68eeYpaYfuwuI0kd2IM42zUkmNfeH9FetTR8YEY9kD1lBs8HbLdtQCb
+dYea6YhgDuJ7b6axCfXK1OwF514WGlbGtJSV1C/+X6E95beyzDFydlfu+EE15py
e+UJgJi0DQSgMvOQbIARmDw8bFVLd0pWP0IV0yTsVYtzjwhVy5jlj0SGf41huNwL
QDzPMN1wR2UQbNIAKa4PwsbwGdWIzWoUGYzAtR+dLdGhoQiT1HPDieioKZhjK5YO
JAcpzm1wl6MbxX8UVwbiXWw63DL4QfXiKTFhgDNTLA7xSwXocmQscATJawkvISOc
JMYBIKgYH99UKuc4FzaBklXaUmZMkx3qWPqK8xl0rjzPLoSCgQ0hQlK2soewdqhl
B1m7aSPQt+on9Ep3y4z2rlMqRztjZmw7g2tGSZIvlLE3hJ6jX7IaAQK+IEWpVNRy
freQg3CwHlznT7n5ywe2iUYnjehEQIalZsrts0f9MhC3J4/FehMryBQwNlIL8pLj
GcVZV8NjaQ2iejBCRlyziDhF1wkHyvLe/lTePdqgmvlk+S/mkN/z6fEjA36YbRHg
MVb+mtfb/OUhckNNnsuSAaV8RQLKLD9mzWgbQCPSt6Q2mWGJEHLAJ8UAHxw52V42
amkzi6THRAf3PH81z9DVuYLZRxoD30cIcHb/moDYzVuy6YaO8XybDogb/ny67jck
DZvXnjabIlGC+guK6iQkwVFSvBI9Jn1KIZc9057y/PhcBK29vrHBSv2aatLBqy1O
i4mXMj/YU1KVuAdyNpmhxObXaXR1mlAQ7MMLpumAVeM6yMUvPtr9fZ49N+tlzOSi
ILTjtKckJaYz+6O1jAZsAd18ryuRberVvzYBsQdWG50Ppq1lOXeEdBLmU07Ny0OE
Vnp7KObYcUb2oqfxownLkV6ksFm0R65y0Vy8lIKm3Uwk3C5aQb7rvgDgS2zcjZ2T
j07caT8eONqGPSc/Zvo6wM2TAIg38BhkkWm1Lfp9t3LUabSZYJZt+hNTyPcKPdry
P1yqhA4efTele/Hu8uvF2haNBV8TPfIFldk1t4ijfcaFNBqz1+Taby9mFiz0cIbL
+7idkAG7q42wqOI2niYA6fUWQkVsvNkbzIt3DKWy+geLQ7assgRz16ymS/bt6IB5
WUXzjzn00Klzkxzyq5aGrSzTqEP3mEJ4ScoeFrmYIjTACTPF28YqDUjgu0RYSt6g
bxWhqgX/ird0WCC0cFQGI4925d/fi70NXtqfvVYAphMix7O5WXC9AC0XNoNq0Ej5
TAluL/zv7tl4kRUzpf/iIGwbi+4IIBhxP27WSz+v3Il0g836PA3jioxOA4VyvWQ5
ajk4wFIZ6qOwE9B8DwxNZUfhG7Sj4aB98H0vlupKrRfjWh64VHxqTHPIQtDfoMVY
F1KVXrEMM/9TjKiqA/VqVAdL7amPIko+hrIaui0WKD+RZ02BqSabvGV7It3yx/aE
GC1yM1wd0B5fYyH9EqM2Ue4b1tu0svxs0ZQirja3Ln39MHjhkPUwgv4NfLLlTrgT
7R2agN32EDIpd8IgyaF8BOTvfYA1bHWgB0FketE9TuUQszg4orIIFIt+BWvdWQ/z
dcSh7Dd2VlosNVA4syraayR+0VZCR6WBf/vAq3WkVOmqPTgoU59Urdcwp0RodOjF
bClDJBK0VfcL0WPQIsWDhod1DTdWu5aWFNkoc/s5y+V55QBETCQg+4T/KuBw0/LK
j0bkd3C451XLBZWtQDOw5Ap1uEmoSxpwiQZI4kaorYN7j9A9vRedY6QZOKyxbD89
7CMCqfOwa8Nxp4VCNaR5BDq0TlBJF6yBVRpdw81IfRJR2VFsVtTh1QSOlDu3taEf
bPHI7DsfLblQMofFEDyaysEOa5GazfA8/ktVkCN9WjOi75fuanbkdeoBQNpndczQ
YmF17wBl79JdA05/+NwcHX2/nAgqF8oaGPJmooSyhmU0j2YPy2RGLcZdLT4Vt8iT
ynOWAm30V83SEYcsJ4GZuW7BYX3LD7lWeJiLPhDg7Q8487/SF5d+1O1uDm11E3Em
qlYDKJkq92KgrIuS1oLhHnHhaWqARJrCMCLoaUegbvkXKzUvkmv3epEob9yDLXoG
t3nCOX8TRtA34Uolcjar03OpDOYpyiikJEkfASrvNZ5yKHU38Sc45dO/noVvz1f9
ZD0AghWvxZ/HudoPV2PqvCA37jba2OABiE/QhgA890acaLprbpFojpuJZhHNT4TA
GY0vgwAclvARYIyq+kvmxkxWYBMxrplZsJLDZQJop0cZO/1+twhEdRFpdP4bBQ7V
8SYLp2mtO1FfxJsLjzkAf0HPKBIp5SKV0XUaM3ylI2LXB/hve3WD9O77y0Cls9b3
5PwHOb/u2Ze5q4hgqO68fk1HdYRqp6aHsYansoD4eIArHoX2qAz4GM5hPxzq8OO1
1HhbV+J+LSTPhKUNfe3NjtdhiKBdrdsNV8qXhJ/cbt5Dw7T3K1taAvxtwz7YlJ0y
TTCOuE3oQkckba55mHAPbkVCH+FspOzX9tBcQOdeHaJdztOJvSiCR9Sxr6UB60yB
iOi0cx+N76hJ8gjWwMvP3WcBLRidaO2emJl/ey8/s4qheANQ1JWHi7m3x/afXjix
dlcW0k18A/5UipcOfG1jWmLDTAQLuedKUWoE7H2dZ712+QJhnJCsu1dSCFRMVXRY
5I9iHV3HNMxj6u+KwjF4tFdIuk29A+MvmCnSfjYFjqjq4zRFRrx05LpTTrh/y/FK
DgA+BuDFuKUSSruRzq3sijlQ20Mn5KvrraX0HVkRv0o6m0Ki8NiWnbI5mN++/9nF
H3LBvpyHzVyBgmLvWLegECovv5sr9PCTOcie+ofLVf4qbA7zmIYLy/Ne/VgYb2JT
YRWMI9ATjVQ5W3zSUZXqllgmACVvSdWFdIkH9ulzhBJNSc9WHomOW+dNuelWSATc
t5pangIgtxZhyT5ToQdwSHMOLPj5BIytlj0sjN0p3bT2J+Zx98VfXvd0WYm3ATxP
KaiH9wDiF4d8X3H3YtRtMHgDuEXfSUrj70I0YeeTZTKAhBHrF6VAHrXhe1wJ87Dc
fDjluxkgpqx5LBsKvtj11rlAdJwhCKdsLHfgogonD6hIVmVwpAQ+CGAfYvIWxPDX
k7jKXJ1x2hemJ/pwTrBQlH7Lk5boLvwah3AfnLKCBcmWZPTg4YMfb5OVvay+5yyY
vdYu7FsAj1eNuWVoXZxWp/zLUEvgUOoUrVBz3+ttvJ1zJElBOhNNEPEwRMheatlp
BiMzUgJ/f5Y6DUhT83aq6GUfB0sap5fAFQ0Nqbo+fFPH7LqeSdj3lEiKj8IwNe+g
xRZJlofj9vliSUq6nPWCIMh0OUgYDvo1cdZGndqTFTGlgZjO9D9eTCo4XLPgGSWv
+Bv36gekPfUYZ7WzWjrisKpOsf+NMrPKWiuxwfLbc2Vjm5xfCHkVvRqponO55y1a
L7QA66olSoas8PNLvkzHxMboiLYKdzDHSaZX4bQO9iRObtEhb9BDWSOMfKs+rZ5l
oynDyiFnZc9V5Iqo2n3hP3u4eaRZXf3Re4byY2xSe9YqkKcU7pFFtZIVZkHcsxqG
1SAqAZ5Pk3gVRPMyFSgD3K8eakZMyOBbJgGWt0v0FrzcIxjY9PRy+Rwnk5ManX+p
3HmdKBUCJJE7x/9DMVLgabKSjv9xSB/WwZ5c6Fw/ngCChfapIL/QVOhg1Hu5QBYH
RWy+ErR4UIODVYAQdk/Fp8MEbKwI5pto7Mcus/qCtd5IPus9lnRaeUhGJy7f06c5
0bxxLXYjlsfhMO3w/nCUkDFPu7ARRfyLBz3pqIqd/AVH/oQBbMuw0fwS58BBHrO6
nnw7FnZubR66qfbK/ikcXm1pRZ1yL+SzTA9TRp1cEhOSnmjPXhL5lb1rnBU+r41G
rjjnNxbPImAPE4PocLx+qVDvWgOwed32pPdE18ChfD7pN0EyKzn/JAttJ0QZ7mBT
tgE6e7B7VYOppP/GLLgAqKjIJGOGdfx5yQh3Y9Qr2yUSyP86EzwWsqTFLt6wPEUu
nyZspkD/BbjjZCpm9jpYRbPqpSwupB/S2z7hlB+Hs8i4vP0f3ryrrVyKQCflxfoB
npCuup5153OpsWYr8LfZINgJNO2BLUfjpxaTpbLjLqP8kd6zt/dkyhmoWtvFn6Ai
gywOVa++SbEnNx2jZtfwt6Qob8MhddpVVanuZjk/O4TbAF9wjtPArUqf7CRVALCG
aPwdVtfvGpy+UIwB8a5ygOU+XWTWWNfH0znwmt/VrW9mTkNe1KP1jXaQPmACWZd4
nfqDS4pzmOL3KyAfrQBytmkhvyWT9X3NUegvd5i8v4eqcz/nXsLLop9LZAjEBM+7
A98+zsaxXXT5RnIzcS/czzwDEVyCdTCUvGtHIfBaFRSesg3KOxIliFRLS7lh24mQ
BSQLyxfJGBGNornG6AMuvTBSD5JuYW0RDDDZmeEiNhOFCjkVJfHRCOqSHP64pNgC
M4YhxxHnMQnWoWdgIDdkYOaHTaTxiW4ePM08Czxc6F7VYKk4zvDflmJxLYOg5Fxe
8UHJA5dnsqI9G4jSwwzaZ7sDDAbUkWXIKRqq0T6VRxPOSyA7mj7C/DNENSjPvgEk
pjUX/XwgpuWivvAF6jDhmbwgQjIcE/LxUC3QESDz3D53I7hXI14u50ld7rrFcy+1
ybzJCqVWxbXWXtMQqrmGiMAlDQG2aiZj8IuEYODj47R/SlAqnbDD8zawyJzLFW0q
JLZVxOweYilQwiZI22jTqk47qJefBa6/cUTIyrcQkHN5f7z1sKCvDMhzrZkSHhZ2
lK/+nZ0qGQgUXJRhPxloOZEvzoVaOO0iQ1OESKqHCi4HZmpEQk2nGqWkF4J0pjm1
U+aXp3bLXN+0qDE5VSPmdAIQ2rE5tZWiiZtsBWQpl2DGTbifL7KE2Mbtako4wI1i
2JZDtXgLf4mrTHy5aRg9DpizXBIlrsMq3I1gpMxirUR/5QNftrQG4KyK8++TL4ar
G2smTtNUwQ7AR1J5ePmAdH39XpNyyAp89XZy1vUuInB/2elMtCt2t0LxCZ0Uzwey
G6B+cJx4UOSA57kneUMV62o91eHVdbvk57b/AQObZ/Xa0onBxe8+8A0BWrRxYXl8
pnBwxHcvgUszdM+GYgiGTcga4Dy4Cdhdmke61a4oxcCVnwRyAK7G/sIoHHIw2iug
8h0nRIzqoI/546xYI25CRPigZ3GZM25W76NLtfMrIslWt5SAZexOIIcoSpZULnCC
oNR4kd2jfzwP5erQxrnoqEIZgGcEKQ7qRT1Xop3ZvOEbE8G5MFmfIcMe7moeMVGO
MdiTG3yncutjv8336woLOgUnXMtCDZU4Saq73Hq1n0N+VXUCtqmwJJcuWoP/Nvoc
lxVHxkcj0eoNkYjg4zWHUSSQi+LTWX1rieKJLlrDU436l8FU8zIBayCMDhYDe9cK
yegSR3c/t0K8AeJl9+QBOGz9BFHBhSacxsH+7V4whtQBcH7CXgdgMIFIRUK/iM8A
BvmJnve4UtEc4BB/6fS8GYAYynDenuHmFzNMOuLmbi8mkrCIqwRn003xPO176n99
ogYfLXmmrplqfG4wVe8Dp9/ztK+nNQjYmEVHFenYbqgbIKlwuYgUFcjDL6bvHgJ3
OA+cCYQYt6tQtMgZ41lcBxMc6OCg0J3DosiU9DydX4rYagsgyFfQOiCQghSAKA1v
uCdBVePNBDgkrEmr7U0f0mENw/ed4lU0ea+OHuu+O7ip7WEQro/Nd6NIhtU3Q5N3
BX/QLwJJLjumuXf5lfmSz8lFnhOV9NRodFg0ysGOZDA7e4PZPh4pCOte2LHRCjTH
Wuxis0rs3NaQrNCAtWs+ALoMFJI4huQBXK6W/VnNgYjhkKc7aYwz1ibk7g8qmhFa
qvk8Bj46DdXD8Eowxbe+foLwUTgmPERYYveJLdkDBnQwiuUFicDu48QM9UGEn/l2
NAoOwSsOroSExTK7uEZDF8ypZ4ktG+KNDeoHV/gDdpEINx/yTeRDKwykx+web+E3
ZfroMgDixQrbJzOs0xW2H0pNrxzjnRgpaWSQSBgg45iblOa+aE7DQLyhmMXY58Et
tNEFLl9kjXh/n2ggGoLa1HBQTnsNwrmvl5AY7uy6svhBiTfV71x1BKO07L69781l
7xX0uVkAvAa7huJi28boFf3LMoXy7YRdqxAesUddkW5rFC1Dbf+Fnwq4P6xHJ5oY
qGyCQCI+Z+PIrLfFktz0e1LQIdpNB0/qOKX9etKGqEUueNkgWkig2ncyNJ8/SDy3
zB3qX9Ck9LsnksghUcJ1N8kZGW3iK/15L0Mx4/4vXnav9NcW5trkW7CDPyNMyDSg
1loNtbgy99ir+2KTO3Ts3Px7fIvGrffMf1f3Bm6epvP5Sh6vbuZlSek3utuN7yMy
A+LH6TpdZ3L5jnsoLlwqyYlHIV7Uf8wX6uzJMhmBuOGe64pd4WyNNaIXhd+njgUl
IFOrgz+d2HvkNNLwZGHF1xuXFiVHufa+guIVBv6loI/3q6Qy2stPfU43gDkCV+M2
mvlvsrQDFtbIrzRWEX8td5+7hVY1JkUuBOfq9LczivicnGBopcOJgGpLkxFXdSZ5
l6DOO5jWhLVP013LcKcSw3UNBbxBDLAmI/rmtJiaUEGkHefhqKO+6OBrYyixu31D
g6m01xja7WQmxJGNiOma6mZOrVFXgD9KDdJCaAc9xfLs4PxFHZMvsHXIZQYpC2EP
U7JtNHBv9GmUsdGhlNPYiRUwssy2aR0RSIzRstr/eMYcDKCeGe25vm1TabwV3txu
QNZ8T2GFjWuH8rITD2G6HfxtSeMIZBBNDuSPuKu0mW1Rk6vLSLaaUF1MPsWwSUNR
3MJFoJy0Nl8l6v2ngyyXL/8RturcUjYBYaLnh7KXkAl1c+4y6oTzIz3ijPWR5OTD
PE+wVyRzNGWvURxmgFvOqP3HrQzB/mkOc9AFfqalyNzocUrYeEKCki6z+eiNbozB
8ip0p/ZuZTb0wNZ6TlEzbftUxNZAA0LkdiBv13Saj+az5PrASJjTs0oNtvIfCoJ5
Qd0QWv+R5yzb4vKridD2Ml6B6oQiPnl2lGrFbp2pEGMnLZpR+Cy/WqRVNQEgclLY
7fYU1XXoC2CcU6OfLJ2YwOQ9gNng3iKxGi0kqXfFs/6E1p4hIbh+RcNzt1hnmcZA
OF5Y9cFUbN2NVgLdyaqQI0sfyMJeUslz4qQFlODUT9y824CLI45mZpBVW5E1VeA6
ZzS5pAdIM0UAVwSPXuDJhKh7Ee2PPNgft3QUbV7fLva0+WZRMeL4ITecJciT8quW
OAy8+NWSned0aBXHNiqufb2pC9q1vZerB+ubpmrdfvfeBBKeJt/iI1FYq8Dkm+Ls
u9HjnZbLBdeUAu2VHlZ6RApQ5IMtiyBCIh+PFG0sw7GForyi6e7vOcMEhrfd72cS
5s+IxRgpT2JHElt1SSWaAsVG54f5G7NkNVvZ25kQfYeshe8oR5CG0kpHaGPLrV0Z
H8Uhkc+pSjDRE5KBv6u2XC58+HewFn+YTksz2/6hGG2OyLuFnAzJ9N5JBWweIWmc
49kOO7CdxWZMjwVathjanw8tVbKDW1Me4F+wIvHM5c9osRW7wqXykoabTz2UBdUX
DLjSEHZLajM0lkCdeallYnc7mMeQ32G4kCz5luL1DZ5X07M18TzblIS/ikZ7bsfw
v3IDFVGC3wy7dEL5KQS6dabmy7Ra8NM+F9SMXS5+95e1RQ2Mj+tLF7lvPFS1B4p3
TdCeKh0P8X5vuUp25wOuyflFDvaYlliey0Hy0I4Og+4w/WpC1cYXH8vSge+eFZPB
dQsW/FOdeuVGsgradXE+enJzS91N7ze2IZVgcDdH9gGrRrmkE7LZGvB5k+pU2U8G
jhUUZsM9oyYx2jHgS3P3CSAOy/8P4CIL7nuWApsegZY77aghTIZTOp+ocjmFVSHr
xT5ooUGvupxITENr7tNM0IrAUHy2N6Z6cxMnDVUky2jTYfJX4b1utdnjmG8cRB0l
KKE1mhPkUX962MQJcBOdQMuOPbL6GFYle1/L08WMkqMvsSa+mfAmeTcrHjAZyXui
hdnHCPZX38Tn+8MkzPLsI8ZYHqkwFZVcUlBZVGs1ofXLU0G8z87rv8nPuiwHjEEv
AzQRlO+KgxcjBdrNyjH3+h4O7Y30qImW2uP4gH1nL2/Cy9VgAlsxxj9RsCmKNVvF
M8DcsIG97rjsKJPsl5GuoczPgnhV2tB45IyoHKk33lYKr+nedLvQ2JYnvw0QiGSn
6glStGALeGVFkQ7FYRu1H0jFyIn10D1y1DSsbiau/VaFrprabLUjFTgLGEFpWfg4
N5aliMh43m5YJGPJtMeVPq2MJq2O1snekMPH6tUKiLSMVBdfNzgm7yy15PqjUW//
okZ72xFWq3wrg2UyiC9NlDDxkGSZNQypTQDnnlkXnJJwOeosy22/wpcQQCLWq9kQ
hkXmWPfjRkZN744PyLhYLTVR0W/NyYFfyAxAnrXTzcYCQwnlO3Lm4uO03PDQpv+8
7RFhEkM4UVuf3W8//u0hG06T5NGK02rPQR1z2+u5na/0CCZfZP1yALRCN5SBTjgN
VspyuzQO1LZe0r8tleKXJpclT1jLlunkt6VsuxPt6v8xNLRcD8do/YGtqDhYjWbT
b/MkQr11RHA0eP8OgOPaIKXXcXYDmoET/xKDObtb2BBx5pjrcsynJ3fwYQnS5Riy
QLgGgMNGz9umhvBglXGX+JqDsgW/FAZ0ttnsq1VZWp1neL+PCqHNxL6cw2Eatq1+
JIi4OF2FC6j/hASwPuxB/wNn6jqmGwnh/L0W07mdrYvkfq2wR6WaAX/WHDnabSqI
IrGA7OPfpp4rnkE/xRoer6QYCDlub4u/RP2j6dQNj/Vzo7yzB+yr2D+pp7By3NkS
km5eUPqz/zFexImqyGngxcD+xJLK3jUa+5p96fXg9Z8vgBI3Mukch5txYpFWX2s6
3M4gsmc8HXHy6+Ub0r3Y5iToVKp0B55HmCwOT0JbxUxzctrW2mZp/vcxBPx5G6UW
rgXCV7RBemjaY9kSxZhhkMk52SB/JZvBV9dfP9KaHtHTjOtj3SYbjY1d/Uvsc9Zt
Q0uNBE2OGRxlNHQhyG7jTEZqlhRLtWE1eUPnbQHsuiG7FlOUuS5ZF/Xsz4Kqdvdq
usxpTSl1YUzfQXQoXDWXlPs0LqyEhnE9rY6snX/VdJzrG7S7+Wq2452G48jSlr3V
9Gr5E2J71wgDntPGJIu7AexDKa4yCekf/rbbfOlle4k4B9O60PHKaHjd0D7fj9q2
JhjrYdPryAK3bt+c7ts+rDejzsbc6L82anWNY5nWeLaord3hQ5IBAtaVjmYERnOv
IeovaSdz4l3uEhCZoFXsJhW6POASeuOKolz2WEcv/jj/NCBnVjfV6NDOYFNY5OQT
IOLjsEWinn84vtm0ctZr66UHvt/uTzrHQ8NTqZ3p32JIa5WaCbYsmhVQupOsNzc3
adUCxyiKBp9T9EZo5QDK6w+L/J5a4Px3lwt+ykEOxsWY984L1uNu5f5Xt6XF/nrb
8UvkyKXSBhq1zp6stchzV3BHybjUfpMo0ndK4iyJFW/VZsE0LYv0ZralSx6BOWHj
QPEYGP3/L6dklAHu6p711MZCVbJLuhzJKeEUXUl2XftrMrYs7s3rOZUPHuTHLW2C
+E0YzrVgUjyBPQiIYfGe2sD7UkMCSx+gd4EqhyU7TNew9iS5cTu4hVLLJX8v/56H
vNLLj3T0QTNI2/uHYK5Um4j7oabO0n2Cd6kAzob+NbaF7tYOtWHI0ALPqAVEhWvx
Lx+qzpCy8wZqVYP1wPlr8ZZnU+vltFMWxciFed69XVGRAHAIcPYpEA+Z8uS1FkOV
BcHXNwUHNP9k1jNP5Owu5vtrGfGhM6M1OIX0NjKDTqeVFG2wT+vX9+I/Jca3zma4
IngUvjU9J5e5pgrfErCXTGQR3hkC1Rc+ya1twIwd31ivAorYLsnKyg2CMYD3Xsje
bkuY32NPJJF6da6QQ6C8ws6ksw1hnS3kb9TkwNo1uVyQA7GfE3XKgn3pYV48bjTV
uVx/eiQkPWwMk1FfhTuqPPdsVc5T9yPDper/HQmZtYL5SQV+TVPPE8tKHnvnPC5R
oEKPvPgv+GAUWSwiLZl1jKGHn0hXU9WcTQ+hi83SK7tu1uE3YLz2zyhEp6QSwGUl
NcEcmLapQDvJ1PohucnrN2Ubh0tXf5OEmWIifUYrcAxCV8cHW5pdh4tdbNBv0Noe
XN2Qq2uFOQMD+BB1E6/7xDRVWMoksK5JL7B1t1sYdmP4nyO6HVAs9YcvcG2JfymW
yne7rxw9tgM9bGXvwIC4wM/qqNwclC9YP3or2+i6eAqfTpu1PVRonert3jaP+Qck
XwKhkFEKGZCPKEec7Od+aYFjvt8dyYZFIaOaQhj3MmE7AbDP5hU2XsCoa/pI79zX
+AYm50/qEU9XCv2Jvp9gMu34nUi2aVDbZHztVA8L0/i9DHQ3ntsa2I//fN16dr/O
rVdvRm3iaMontVDuR3OpNkIr70yCcoEjz/qETKbr0ZOQ5ln4PAYSGlV0nWuG4mFu
1y2/YvktvE8T8Iua6uZ5Ej5Hwkd7U4WdnQSE2K8x0tT2FiAYxy3z0bvlWkgQJIZG
KH2sa+FtKsc988NoRnCEmzxOYbbOLoz4piFL7z0P79supqNBwuuL9wGgc0a1t3Hf
R2wohbdUtleDTBOIXUsOjjoZ5fH83fq+J+0FaoHaYs27BLE2UsZL/zQGZ/maxVsW
sJdJ7fR75yHGw+/+usKBBRRCti5Zq8igad7rhJxUMGx2s/JKwgFfzBNmfeA/LAKU
dcvlHECvTTNWjN6Eflf4+COkV46i9xf5gulpcL3Mi7e8CKVaNzsQcrNJIt9Ybbcp
Q+8sYgSv+cSwLYdM+ksexTgoC7e78+iUf2AqOUSzH6rNMw8lP+2wojFVkJjaM1CL
Q90SIhLMpCNPgk4eVEC8/K63NtX83wq0xWWXoSeP1pxb8kfrywrvFBJz6tMzBsDC
xHHK20sRm1I8hRDkT4XMsbaxc3vXR1xcUSciOnc8P6l4fz9kqXtzT9pszPLkqUfQ
K8twC/gzB7UuW62aCPPmE0BpS6w940sDHcnoc+ThmfDWUrsUH63jQ4a1LbmTkCf4
z2C0ERQOmGAnv0NLOVz8xfJ1q4BtBmokaEofKvGCBetzVaOwRZ09B6tnF3NjoiQ8
5nvA8p8/Ny4ZNl8Vm/mfQSjozb9IAZCAaNmfqqMBsp5EBRf2rU5Fci/txKjOjhkH
Digwh10Cy3zQ7tAD6EvvHr4XtptErR20hfFIjwS9OMbrJHvX8SPliGintzArUesR
kQXkWXc+P7FpHKgXjXV1mR4z4i3m07m9wNWdOzGXpHjAuZ9tUBPibKFGG1I+iFCh
wM0NEjmhZCFzEcR0VJwlOegL90iLNS9Wy1cbzOufOGmXaTWkJvDDLhK4K6VxMB4j
vearWtfHlNg4G8sNHD8pmx96PUTZ1Yci6QemD2fKmHbtOrrrT5pT7aFbBn2942tz
LmOC+00xTDFofakfks56kAPOWMFUOiR1NOtY53QML0JtnstkwBoaryrq9GICMxRg
KmDUPYUzv6q+1X8xYS9E2vvvP3k+urQSijZk1PFpttx7qNdn2v9txZb6EGSCyt2B
6SNxD3OJS0i12Vj1vT7IBAzcPDtMwtkJje8l6kUp0cGlCu0Vc67XfGY6t7lEm2yS
r2++d7olK1OnXKU6ePEWC5X+HQk4DVzpva3GsRTWgF1gXFMLh+CJudLKHoAwQOZZ
ot9E9QafnNnsg6bqL0aoEuu6/jyFEBnty55CjOw8CN6pdoRWTerjvS6IbQesm1xW
0SoG5nlYS6LO5jjNWKUXKWbgOTzfmeGtg+by3jR5TUpfRjVBg2N7yu7l/ozVCozA
tqcw3ZPr6qaV+nOBXN+QpjEVetaUw09UV0O0tJOQvzVibYP77tyIhPEiSJFK+4WB
9Qvq3udOcWnGv0F9W2poQubnh0ME1ytUBi6092krd+p2gWjcUW91IJfzVYTHzA1n
awQ0Me9uKUPeIH2B+nUfqwdFQCkMD9w6SjDAYArZNOzx7STMvNI0a+ySA4h3SYM6
bCKApIsUhV+Tr70NLw3NbVb4GCLf90N46y57eZBT6K1+mCnFH7Mjh2eqTpTeGZZj
iwb1Il2FLAuyEzzxXwLjvgJS5U6gVZoSkFlyQip5plGaBwGzmueGe5JZqIyscWHr
haCqLhsMc2qR0SG9xgMCSm6yfwwhyf/lBrwXL9QNj0JVevawh3ZaEi4FYF610nWu
teFVkkppKnMD+t1pROMTBPGJKAyQwTdZOAnW8eogN2ugQSVdO7UJNSYTS5uWKiw4
tWm0r/ZZzzkanF4ZhJIZLPu6o3Ht/eqlKtMOOsrbVaZjvcXlOtEtY3TWE9yykqMC
A+RbZUWN44FDvUTibuC9swOo1QTeGT0HjBO/GuAzCd33afNNGqz+l4P71aBrn0RT
Nl1HFgVHUUzqcJy9g/PG1lvhV22gquQGdLUsGzgkIz5bjEEALzdiy8mcP0QtvX+p
QAGUmVVwN2kpo9/I+CKZYdPw4zyD8akFKtdcoN5P5ZNazSH1nMJaNQYX9vV9/waC
X7UMZfStKxubXaSVJhFyRpSv+0whMay5f7din926IBI9RJjNrdIBbLjNfNv4CP9y
PsxPozLp5Na5qDuF10HQl6Brhud26ZQRkPEX0NHqXFFv7Q0rAgs1srECEbOy4jj4
QXYF/RcmSpf0Eo0ALnw5sxWjmYgDou58o2QcXI3ClemiPWQtb8v7Z3FV9uAsfSox
9F9XSUXgD1Yk9cQ69VUGZGa0kXyKcRnovo0sR+k1Cewehxm8dQyZB29Dk9rPoEMl
qJl6QgsY4KgXiPSD93JkvzzhxCVzQTYSZdmc3TlaTzpbgV3MKz4nBj1gHAe3bsVx
9jod6foDdsxhKKSOdCNl0iuCdo5RpuDHXNyYnbllDORjrqmM7ifkfwWJGBHWUX0V
1ke9G72LH5V6qFFO/12NoOhVzUKzDDr6HEarNVnWoHc5aPpdf9X300IzbrPAJvyx
DvkmVgk+Pt8dIyPuArIhnOi/tymTxYfZYDZiCQw9xXqvEudXpPKybPDYP8av3KQy
Yt+sIynbK5F1nXJdPaQcZx++D1A7YeYaz7aq76ll0z79J6zACWeBxC+ySqL9NWp3
9mhOOg0TkzXWc0EAmcrsDWcmP2I5NI9qkVnTshfotbUBZvjDIS5nShqlJ/UqOejl
rWQFd0t6MBgL7e3vIIgh/cRKK6eF/XWCBI7yCHYBB03lhQcpDspQTEjUzH7Bw8bn
w/6duqd+UC3YmygQLYM2FRHZ0auaj75M4DkOVUVadpL7prEyaavik/dik7mkkd9V
nTdTC4siMpw+yV72I+9G/YUalFF7/xkNeh29jZYXdZc+ZJeRfPRWdGbqjmhqL4Iy
eMVjyqiHnVGyscqituYOpXoBmBXx8G6gd5vducBnXsaHw2ZgmZxTwbCz9Qyl1Kaj
22hyf/Dd2ho7CER/JmQ9YJJBNx5Dq3RLFuRMeGseRjKJt9nOd7e7z1CLmGjYuNLh
bTR0A0oaGB9zFsPaiEUFNpupeLQI7HTuM6OepnGyje6WXmRBcHy7D1FiR/6w/ocU
lIvr11rluKVdsv60tjbkY12+3W+1uRfa4A+sOGc06LN+MD3M3t/0z5zjXGfeDxZZ
/op+SK7tvIP/46UZibcqEFpkEeuBUwKHOeornXLsnEOEuXbiR+fSvNSZvUBVw3dP
ooZh9Se4w6AYhla3a1Sb3AT0O5FEBqG5FryiKWnskzqWE3OQbfZdqPxPaBsnA8kd
l9RbroNzyv7bDummfwfh6s/FfyRmkweE5VdYWAYm6bTEFI8dZf4dSq5kv1Q+R0t9
RBgBkzvRX4J9CjiX5ZfIGZ1XDSubfR0pEhAB0VW6n2/G0InjuDWhspwfLJmSfhy+
F0fpWgFTlnjm1JCr1uwYia1ZUvU6SU/zYbnSwJpZ6KsoWEMucUb0CbIeVWME26D0
mIMKtAj9SzyU58DpQbk0QQk/RW5JjF6JP7zJY0ePY7k906Lf/eKy3Q7CmbHYLPdY
RCoI8EcKRLblKJY8HsJQ3wtXVhf9gvq0CXEm1R1efbB5QVZGI53HlkzGEhP0yLry
lwl47MOE7gZ1NhiB7AFHmGRPc22oVav+LX1fMHHEaLtdbidHPnZDwXVfJldwq789
pd6ZSg3EEDiNtFsknosjoAvPE5DmHEWR8tcrX4NlfA+emg6V0rJVbMM4WOblduNu
fp0gy3unudTkd8cJ7kTFDWPlnDvQpujJuDcIzhUY1G+MiGiooC5dt6yt0ekfMJiD
8zZa1tCcsC2fS25RxmNFo9/itl6R989j99g6BaE2or5ipU9/FrPLPktr6BRpshOX
KrkF4RFIekAg9xZmlr2NHLK2t0MeUyXMIYyK9T+01KW/0QawQuiAr3vM4cvmYCDx
y9PYTxL+GPr/zyYNm0ss7SXptVCuFgyGrHyhqfbcMlyKbNVtSIucRfAFjgfOYN7L
E0xyLA4y0ODuzBlOcCwR8EwaWXLnlsAh1mP2zJUxzp6AIoKB4NB3mSO0Jk+5NNN1
la0w9vc6Qt5Ir7SUkXgSSpiEmDEQc8hxuxnFayGR4ju5YjprCR9IJyQgtNRl8gLy
9CyaP2LxTgKAZLCqyD4tHaExJbKobTLrzyKmAF127updzMkXNNrTrnOe7tItwPRz
GZLDPs3jgQIgyqckdAH+CmwwzTK1pbYLFGsHBtWSZAlOst8Tyh/otODvr8QjY/+v
6CGK73SFbI5N8ejn0fUfxfrfWMzDwfXp95Z5Tp2QJ8OSVdfHfxkkTD/+PfTSLwHR
ahTMPMdGubx3xcbVIS1Wruzx0hhA/dDFTmQBOTTreALe17iYv1qKBpMz4KS+iTkL
3VEtClLDdd40JYSSpRGV7ticBzcUP9geoqKay0slfAUXQg+gkTHnNmzozOQexHz2
Tihs4AIeVxgJ9hCjJalVxvXmtqGsyH7VUAkUdCT4PJp6LhYeZDoR+MEfbUIVmFcK
mo1HcDgmQgO9SqtQx9xWfDO6FQ8ilLNcpOwcUnGtEzcD6JxTasd2/uoQVCATqXI/
AMzF87DdVACvcs5ghVR1tkkxznzrdSK0M2OusxQdb3VFjClJARhXyuTnt7ylNWFU
I38k0s8ZaWo/fYAli5itFBKV2UZzAg/SXp+vKuNLj4W/QBMqsCdpTWJpf6rcGRHy
NMn3sYHJ7VEu/gU1+YKb8f25DcKlNc2w5kcCmFgnhx1h+VNjj1ktP2kRwsHGJ+uQ
tk+CYb5oGmjhK3ZBDAIEpZwSARi0sIWiyO8d9KX0sbjmpdMDeDvAaOLLukhk5Zvi
WW/dvj53iAuNRgSjJb21i12ZPispXRviuwcE4AY6UXFtBxAE0IvtHPWSZ0sdY0I0
+4lj+A1qHheVikdChChRn7qR7PxvEkD5bYz/DpAsKvQGcS1XqS9nRbVB//tKAqPq
U2jnFJrrHU+leZNAMFBF8HuyKJzFPCTa2SNgbYjIONuvJAnncwGL2nkmEYs11lJL
XzYDt9d8lrXu6QvFBIuJQHTVh+E99jA6++rxJrsJsRBB1VuD7+N6WvmYKpQ9bHnB
gNdNUDrIjkfkpH9qAyW+RDP1PlKzyqRVdRwWvnvyiLRZxrcJLR0IkjDLG9a9Tr2e
+swlh6cqwB2f5jWmayheWc3JsPCIprpptVjHF4dTazUaUR82KC9iW4ohRpJ2vQWa
7SNNGRU82ejgEMHVErqsbar4bnwzJQtXrIkdizVvyKazvqh9j8sap49fImBuMuTv
IdmAz1m8y1Mch7jWDopyKmy37/zUWIZNByG2/H4KJniNGjMVjekD83EqaZvaav9L
J7KULJIyp40chc1+pptnnepwknVTO1nh1DGiF/p3ikHrCQmRPPlG7Nd71/zXVuRl
2rzMfuBuf9/P7eDCsIBpXNg3s6hGbTMXMwsmNeA2yIJtmjBa8ElrQihAhe9l6I57
S+ZH6vZ8xw9dsV0cekQuwCLvEZ/KHaCIRn9ucBltx1Yn/YxP9dL9NO4tofJgx1ev
RRQZveb7grtPh7Ai0ZNy/Wkmt6T8MV3wQ4lzPGxx1KPD7WnudJ3z3OG9cQJUdLpj
p6Dzn4R0sxkimTa4Or0SekY0MgXUJjwj6jojXwJDSnNlvEGE9vwjM8h9NSBcHH3R
1LezuPhzOdpukABhmxbUIcMWdRf1CiUk4YRVz6Xaom+J5j6gZmiWm686KCNoY2gF
MMDI+Vxz07I3KLb+g7Rri/jy+GHfachPpBgFywVxnVi3Rw4e4uCdE8er9qhBl2zX
FB/I5L9HgRN6uoi6cYdWEWjCaXgXL+1/00FBSw2XVHX3DNUm1KO7VSw1U5scb6el
LSuKvXnTx3U6Ssl0/35okUFiKEJYha3oJECwW7zEOTfIrD402q0tim6JNIr0ipCO
xngSO5njhpyIJeSpkwlgHSEP0ss22C235W9p0MEgUp8hkt7/bzsh88HAwfZu1uSm
OEYG+rVREYqx7IzcinsraTg47inIllhWWMZHtQ4NhlXi1u2qIlB7/Q4aUwkCskZ8
LSgOZ+AiTTzWMOB9gs127WDx0JQeLErW5ZRmk4ioJ4I80tdQWxUStn9M6KaJQ9gX
DEhi2MOxdHVrlxKCKGA41CKWsItAdyPoS68GotWReOAl7v1YNJL4lgG/7i8hAhBG
O04OU0m/08KH4emDsty1QaQj9DQvb/w58DxIF2ahv7nie3KI5z6z88WbzkKdM1F6
eHrhqYoGwjoX0udHp1nj28CbTRVhSDCWRWD+Oozy0AB5ewLajaxnN2qIn/GXhUMs
fv2rj6Kkbhuzd12z1vtIwhrFeNF9HjBIAZh7MZJ75vzOPPHASd4x8ekHlq/ly56Z
Y1srkyFJQeWx8y4uSZPbuHEpchPKSRK2BfdaLcHX0Z3myR4xrKFvWv14H0Gnm0F3
qQze5s/Lf3njPzN2IWc+DccSlQSNPC2xz7L45SFFXttrH1+S4zN//04RLidjnann
yBZawvK4uGBJDYECbLTBMB0l/opekbbM8lsCL3/pIyZEimpHTrCLYkexA98QF2ei
NOSiVVpO7cPacjAqZYFq74XN0rSc89gYN1zOtFAGEXkpCT8qDnPnsU5cXWapOlYi
kzjXn7fuDD9HvZ1cjjW9evU4nj7krRoTLWXk+s4ZuRcNqOK4PxVyZWqP1TArF0M2
CldIFXevUsHyRB1ZUS8Gyh+nTgmWCFpGCut7ywT6E9OBWsprGBEAjEADVza23oHa
mVLLePB6amfSlMIsxe40V2FBfoBvcPJ+Ab9V0q/ukf1TYht7gbTYdyLjokgLdFtK
/x7Tj4Llpz62QOC7URTA3SY/XT5W3u8nC+EwtoDHlshIT8QNDyaGugWQbgosyrXo
LFrTXD4MEuPWDMbDxXTII9vsvhQNUBsyCOOtrRdjwneF4Gl1NxVA6/9krRx4wyfr
GbBVMEsNCivbU1mph3UmvVX4L0xeUyiiDUGHo7ZCBxA5/XWhXK/t+nmPIs6A5AC7
0WsVEoJH4d9x/ADinwrfdv6fROZEKto08jyxErMP4TTyqXMR9XHta1C9OY01eHsy
lQlwppOGqZfyiHMUjU6GpCfAyZr7/defd3OXGTBfPlmbl/al8VN1Jx+LX2xznKd9
fx5Mm1Zj3R+3IVGAtun7VgHFQjIx2RskHixR26HX6LjHthKNNbYXcpPggsCbVKWZ
C0RnY2z7zRRExQ46RFIZJXG+fj1Jp9yrH/YznKxGblLpedNxndFn2dlUZiI3qTsq
aWrktdgO+6Lsb9E2kvWTOZc+Dgbh2RcvPCxGplmmypOYRXUMTXI3lA+PALbhA2IQ
UYJ+LKD52XMjcecarZ8UD56zhiNAVGN2lUAjRuN7A+twmJxN3ubtjt/jEwr6lIHy
gWPjJ/ZXdwAAFXRG/4K+AkCc1IX+nny/vgSJ2B9jrEoQWMZug0RQ3BN+FfdL4KuI
KPXYMNJmGwCXHi/6FGmu9HO9Pxy/umcZ6EVB2mfwTGRLwo6RMAbScQpssTV150p3
IbA1nrnPaKKuyW/hk21UUVoargddwSLyP+Deo3ojtAfSLN0QcVcscZMOHx0pkXZQ
Yx/AtnKr+zuDwy1X6zgdnPX2gIhybkHmokmoJOmuzt8Ye0x7T1+UN/rNtU+6iuSE
YxhQFdAasqtyCMUloBYK+eXQEw6e3f6cKlr+btdDHVA2/S+i1wXTN/3KcEO20ad0
pfjIzPpAFvkbl/hGHRQrAF3Sie7VrAbM5Ksq+/HkDT7bBCUov18Kr7MxV+AR1COz
H/1d/mm5lYBdpLxn8jWUGEsqShOFd96D4kM+Gv7Ak42X09FXdej1Shstd6bdtN6Q
4QVR3YnBmIivMyhgTB7Wtoyixu01PVdHUbMsPC0nIkzbtXIJwWDnp0zcz6D2Osol
jT0pexuVFIDnsMJR2bXVmIh7WWsPA+E00UZD8dzKjLyxUNLwmFWDdULbRFDGXLTG
LS+gntqztiI4iNUTX2byfegbEA5AUvD0q5kdFjaYZew8Q4mMZWEGQJCVXLTEML/R
V6e0LrI88+5MHBt/dnipC4sPkrJEMj0mdd58kQ0+qn1uFHBuVNgaqiNgEfeDx/rc
1YXWgGXztDnJQyAL86uN69NeTIlQQVQo4uVqlVyYBOEKsKpZG6dffgWdYdiMlgEK
IxQyo8DCf7X7ndapcN72QCCZQlEx5ViLwVqi55hV8DAlFLIeuYEKJK5v5NE7VcaH
bwigIHVaY6d3KS5ugCN5ce0fyEC7bv6lc7MRVRAMOdiWSWA898SGIs06ke+pkMW7
Jy98mmU0hD0E4tvWudKL8ESbAyIepFcWNQkWWiaKte6rbgUYfGyFNMFLtDAbcou5
kDXj2BQYP2QWOJjYUJLv79YOgUZevWq2PA2Efwq+obg/49oA2CCxmhPifwtyEtfl
47Q4aHJzMEsx6bbp7cwvBSk+6Bot3vYbJlY64O9RIIefuojeihOh8sMtYB02eT+B
axrWa0Lf/tZevqZgpn2ilxcq+p1UEWpPuaiJeVzrCMnHXc755VEqfKijUFrp/V1A
ZHCnqdheiLUM8lhI1jkczKsR52V/1ixI5i63IvjD9HA63DfG7lVhru33ZC9E8VRK
XFnsF9ovfcEbQjkW+VhwEaBT/flcAYbQgP2MrJE/87RWN+IY139dQwpecX4sZfcu
Zf+psuh6iTBFd2ShqiXzEzwIhmQqg6Ecn9jT0nkdVc1QTG9P5uFH5lRcoJ7NnBt6
z2B7/lqZFVc1akEWh9WtDJIQ/rplyucAYPdw30R1JWYHmUa8blv2peoJTpjc2au9
bOtX18vszs8FYeYNrM2qO3zwOQf8ucAcV7VmgWT7pXyte5jreWZfRxeMDLx5L9Cf
IwlKDpBpKVsy2Zd41bZ7MTYmG3aF5jQdtwaLeedgm8IO8S38KJvefjgUsatwKw1X
ok8ueNRJKwSjSssVG+rJK52KEapH6dpPpOyomSJ3N7oPt+bSMxCDZJkw+ZCicb9G
c0FzoqhWoYx5kmHbOHxSX/wBAL5hj1/JS1zgE4o565Ohlca5THAFy/BKUR4Kwibd
5Wq5xqikdvx/7nNbu4wRqehRXSzJRIZrB6NP+A/yKUaOn9pSfeLI5PBQDReADCvb
ueatKJcd1rezTLWElTBVG//xh2ySq8JxpL6gm1tPOuV3uVWBHCbYMZzFSDxYGmJO
4U4kjMGPLXvinPeRtiauP3plq7og8eNdtRDV8csdH9SI9BMC+IAUgTLOej0Rs7ht
RNFbL5u9oUTNQJ2kHYIxuEugJ5MUAHOLcgCzpS2TUEd0NcPK4CiGTVWDk8blk868
u/KorCnsX6nW2yePxn8y5PcOvxh1xSWO5ippqON2fsN0/W6eyjCkHtwb768IbWfW
3+95hiDE2HIiOxdc9/JniDzKEdV+aG/UfOF+aXyspAjK9J167ocomo9mJNsXkNXR
bNWt1fRCv5EsDXeEyTVrY+5JdapSjsqgN0eAZeqeMhzvPcDID1W/njbcrFZ0nk7s
pCGUclY08bvVWyYX2mmcHl7YsUPqZM7+B0uzNh59lAENObnwIABlMkBbMjG466MS
JhgP/6dOEJLYWAqZ09vu1pzBBSF7CcloVjG2SZ1LBMdwFd7EegJPjm3iIv9KCUtd
Pg4JRfmrHhM5d555aHLkgZn2EK3atGjuSj0geM1Uzio6wHOXdMphAfqYDt8fqzTS
whjNYGGb1gBxVOvfOCzxJ3SZ2yyYsefKgwzpersCWDgQPaCgsSVL15DZBC7CwIQS
Jbz1XfQDoeJ//F0FMECURdYWbYcABbJ4qpkCW7+Y8yTjjr+fVcPIN9CePFsBK9VJ
es/zJj33OrYeoDGaKTNPxNutZTWMmB5ktpuEQYa0zWSpcHf+dquO51ooPzf56gRC
NKZW3+5aBeJlrPPaGfnluZLfZc+vefTwm6Bo1JXhPghHg4bH0XeT5LzAHJcal2vw
TzVfMFcEoyE6b273loTRwy85zkPcTKdMhe02OqwD+zPuaV3sp1SKiPBLVQLzOM05
yMCQ+cwCIJELEWLPuZuPE88FxDWMOvUcWwtaKLf5FuUCeRjawBouE5uCazaCW7Qh
rqiNSZ2Md0Uvyfo0n2Yt0hICpiEYYlw2R19RbnFEddF/umcLPhxNgNbVYc/UFxRr
Gg+YGd0HqPvek6Kh9Eo80wuIEZCtGiGRo7meZGhshf0oYGjK1X14itOqbDFIWR8c
9ZrO02QQijQ4gnOrLYcsyfX1ezfXa48ozo58OPIPPNQhl04MZhW04Y0y+kv9afuY
yBXId/zdfwH2/dn5gVnoUkDdqoFS2iSj0PupFuifiKrKDpjuVPzBbjOdEQ1ZozXr
wPkc0jJGa8+uCw4jfitrszZs7/taQbvAniK5YFZxezfpwDDIGyCFSclo7yfT8H9m
qIfdSK+YadIGiwEAi8YePHvuI+yLMBo3rVPrVPMkZGgKKWRsT0iZInzm+nE/fWlH
TUKGf+n2JenkatI+7NlJcucIsGKRRc7IkQkJnt1RKqzaEILf8Osfd/DJP71yoSO6
zcHqIvTJ/i4jT/pfSpgStUrtH2hrZIocVjNT+s5KiY0mKCzkZ+lpJhPwB5/R5Ot3
osNhIykR9NNYWq/n2v24RNqSNl8x1XNEXqQ4fY9/JqiI/l7xncRVZuT7xxKFNJGr
SAKlzAROePftYGJqi+cb/uw6T0GrkoRHd3k9aMyAlBUll09RY7c+e6YAYU5KP3+t
YHDpbzRkxKx46duUGkrR8ONXx33wyIkrRa+j7itkRAG31ZIySc2f3pAc/n3W4Fr1
Ipj9pTUQdYqR3Bxwk/bNVhEreumG/BopyMj7Easy2iupBvqUAaX0+KgfFwENVEGj
OPF9rtHmEv8QErBEJ8NToaidnc2/NGb328M7v75R0XbCcf5XqUkRMHVi9hmZuYPa
9RjdUq5gBkuXJhFwhflxf88H6vksSOnlWUKAPZdEXWylMQkmeX1ilO5vCohui9n+
IeJ2fjqFVfbsUr0XZz4tKmmtrcBcmIjIsX0b+3ZrjrVX6xVlcDkl1b0mtQ96c79M
R9NV7uJGZ6lZZSNks3TSjyXCZyvUCr2n90/4xj5MvHRIhGEo1WN66t7w7Y+Wjj5M
O+vWLuWCw74w97glOVPveoOP+pIO3tCPwaBr8G1OqgZNs6rh5CpSmzRIAYRkiTjU
vlaTok/zv5Nf8OevAHjcNxEyyJBwRDjdm66GYHNGBimNfv5svg9rU5R8pGTwOlc5
cPcHYZp9MWkAIRwx+vUmGmRvLWfCmJp1clVGp/Y627yDniM4hrfE4gX9d+p3DPzH
H+VPsjIixXGsqr9XAxUHVxpxqT8FW+xRSfhmC0rGxdEmPP9N+fxi4xbT7uyUm0C8
BHmY5ZxYUc80rvZB22TQMF9iz/xf5OBKgmSnvwafPRp9XupnBFp0DgzmHf460YwA
vZMI3VUE+6lduMnpdaV858ZONX2p+bqdbsX3FiVUDxLjQ6TvSHUjCRnoS/5M5LvQ
Nmo3HSl+q01TKbahMfJ2abcd+2JRtu9QmssoSLRVUbxW+QiPvi1TVP1lVVD318No
Aw9hNDUdBBGwFtg/M/EBMjiwOU0Wmoe6BE6F2sLRPtrkowdLpzGIk86F19xfn1Uf
LB64GV1oNj5Jt2QUfWk1C5m1kckuekKnc7NUyB57HLc8CCXp2ZXkhQ3OkXQB/v67
6Hg+tGGV4rhwZGnpKBIM1yA4JpKjFZ2O2KkK22CUlbtQ/cNQVoQfKb4u0wwz43bK
n8bTDI++2Bw2cW2oJSF3/sF6wQdop712d2R7ld04s2WpyVJ4pPmGn4Wc/kUocCwT
/svNJ/JKtD900j7JNDXK5JVLLm4qj54/Zj5THfIdcH7XwNbqR2ZQk6MaTCkz0g4b
zJmyFO/P7Qz9TYW5+r5KdUW+xovnd4T4/kGWEkacQNmO3p1pkHAMotpmbWbgs8k5
+TBfgzEm15JqMjtLG3q3Bt43m4qQd18oPsU5K6ApJ5ceRLtLYN8zTP8JTNlNverv
R9aVX3K5w9LTTBeaXdY6yquBGRepQbpjHQTEW+CW3LZ+RhQS6Mxp9B2DYQMglJc5
TQoqp5i5zHy/VDBg5FhFAeD+YU62yiDaM07brzOjkUyCMmDxkJOTEHfD1OOwB37g
Q78iuTSLbF1TdpGnpK/6TtRV89Mgb73lv3zYorpCeg4W8ZlyeWjYHAgu6Nj659Kt
mjqarvKWAw74ofh+hM7ko27pQ0HOEt2PdjBGK6RYDwx4XxnjgP+7WkuS7eIUAyNB
upamU5hCk1Hi3eqU+DnLcHz1PN2wCmhT7vGZabQdqfJt5crzDFQhHM3DVzlj97wP
BGOkma4UW0gk0ZyoKmBwIb/AphNb/8xko8XOwA+RAIKuM+Y4qKTT6L81gWM8r6Cj
1QtyL/I1aMKpovDyqAu/TsgIhPP5JZrepH/+1ZlIjM6RT6Xrr+gTU8FBed1wj7TI
CuEp30mTBpjgXmY9jicLLicBBr3fhluW4T96gcJ0d1oY4I/ClZ9ctiuzP15QhTi8
sYgWVidZ4ce9Q/FaRRwpQ5vzWZnaJQtieMgYhfeBAVaojkrqgGBSBluF4KwBU2+a
bJeUcvvY3W7KDkGm/bZVkr4bRSfuUnNsIB8Gpddxl2woSKL8GWWI76/o1u3ekxQX
oWOO4CA4RAoU1Ddp6WqdhUaQq2Z3CwPV2/HqtKZqjJazQtT4cWcYXKbg15MjEAxe
kmfLHKhH/1AAGhA7+sqS2X25TMf99PmgWEh8L7PT9lCr+3BqHVe0ldWVe1g5btI1
ky5fLvMaYPvoC5L8FJODLG4GrDTQNM0lqemarih0LL9uEobYsXCEH4TyefD5S6tg
k4M1diGe2piOC22qEvnETJR9ovqr2LA/Gt71MUdeVPfSlKzxGxvMaFx6B51vp4g6
3nXjm3r8fIQ3W0vuQm0So9k/OsBc79XmKrSg0W+UbInJQHLQMKPNsrZosMUF3rFc
rOTb6RQkotLAKw7ZurLeDeuOynXxMpGF7lHxTvEFxp0M6v7l4SsV4HQL5Jjo9d+l
Uz0VD0T2hnB3wuoFL+xg4wFAAGsx3qneNP87Eduoof9SEIlW9BXyEvo4h/iH16Qh
rEDI4FbffYvBYLkllGuR+3Q8JXN//AF5P6+IGGo4z2JLr3YuiBAcXepqmF99suC+
cQIgkHiObe4lHvemiVtDP7oBaYxEkQE1eJEatv7H/SLuTmP8UL5Tn+tCgLjbXd2F
hzhB+pR+RYljm0vejevNmErZlJUY4rz8XHo1GDp9vfw9bnQsnDLpkLLkrSHJNqyW
ZuhTVey26yyIKnedWApk4WYoQjUWwKHfUy5cTAVTQKMHQ5sY/TA43OW3Ly0hSnV2
gLci6kGxV73N/DNjnyNaAXThfLrSHW3a8Kb8vNTXt2jv2BkFGBYWz7LXNgtJgK3c
SQFgywTvPXTls0LZQ0CoP0ucBdeI+PFflUbGa2DA4QxQvPQ7mF6ZsV3T1uGvsTZr
WjzNlk5nrFqrnwCa57Eh6MEy5E+9mtGKtq4Pv4dHI01pvwASz1+rJzJqg/CQtDIH
Z+fFS+CPfNVV3jiNDRCw9yr0RS6MaNqeYapLBH7NOgxDN0eEV2MuFL1nHRT608/m
nFsS9cXBH51te/9dtuIyopb9OkHAUrkxdSNuYIBDxpFjLToX5ifEvRia6hL0u9aD
n0tOJERK/MuRMqSz0A7uakOQXW8QcbT56B8TYrl2TNtEDossJFfDv0udtcu9lCJd
4ZfxNu5B1Lj/ixLeNP9YQ12uHc310S23RPz8EGI9DEeYCdOeOeQ+UIwr5W/+bvnf
TSGw3JA0M0HgTLS7U07HrrR9wZD1s4SJfa80kYShUspqg/4ZZQ1tmqEk61S4ihWV
QYgeyf/TwJcaOvEGfELkEtxZMIl8fpnc6y4BUo5lZIK7+iHscGzww6Qp79Eke/Cl
1WgXvwPsyhaYkLyMjAk7xEtCEw2a4FYF+z4dK8nGLNYC59gsOd344hgW8ZxsIdOd
FA2QXV1IQwXw3SuPx4wHDVGBc1/lVNzsvH53FmxuqSTUJdrx1F36Q5jWDIAgS6FT
qil0eI+5QjPhHTHswJExlP8p8KNakLn/dmrqantqhZRE6ldPZAgRWQxxx7Kc6li6
g9ELiwISg/f5/1V4Irtc096W7LiDJtHVhNQg+VXyJbcVtLQNgI+BOd4g+kL6EwYg
SajNYcNjzQLzmYgTsq/eKqi/l67FFQ+5ZkbAqH2UKlxthaeZyrg8awSOys3fgvHK
kULsyX/0/SOG6eiznQR2tA8l2GdsF98WVvYkpZvUuDGdizqaHwIIg3SWTw24E+rn
9p7CezB+ubVFjQZEzYgk/M/IfU6ijY54LmhunDyVjL2A2co2FGCVHM0pNQSCoot3
+w1uHW7cFHDOKQ3FfKgndjtHUnK8iz9lGl199HNWlOrjhc+zjbYufSqZ8y2nlmxS
VejYBQzBe6veRXlO/re6/hy0/8V1wmwCX3GIxTjp7gUFmEUVTxJPU3hTLEIcjWSJ
wYGLXOwgT8ozrL+c5XFW0FjTPPydeUSrSSm1+ZvnRZR+/vE4XuYezWsCv4j1EBXr
ed82s9DNDZ/HpT35HstBLhZ0WABmWqWR0H5HMRo8hz7a0/Fj3YGdPohBFZeMX8M/
IRVKXcCaJ6+oc+SPmXv2eiJ1bKBoS/0Ap9Uwi/wh4MpyyxbvuXbSm7ZONiV9+oU7
uzWrQDbZIPb/4vbzrA1CVH0fwlRX3Wlxp6JFH7lIkbQj4vgULif7bTrNZy3hXH/g
i6Jon6BvkbzoWH4uH80IsEx2u73OAwdudP2W9QQBWw0MYiXgR3UGyF+9g4Bv+Ybe
n3xEdsXMmTSHgSxuQIwtugILJIfzES5eRmeOTcWkvSBwaKVW0fdqi1HrmRoT5B/7
/M+RNIxL/3hcBNP+Lik5JRt8LyndGCzIpJZokdCACY+qBFRWxORudLNhe221znCk
2/2q1Xi+Yla5q5S7u686ichBdHyaRXJQLhw4icbMtzDDVUv7c+mlv/BsiJBl9arc
yjPCxf2Xcpr9EWTwLSZDrxbO5/cVseWMsevaSfWV416xO7KtPunvV430tzRSqKiV
Uyb8+p3yfJmvAIq9YDAaQpDx2J+eIrQ0+rwcO6+qPDmgDYUv7OZc5jVJaMJMMwNU
V4zj2PxMz1GbcQZLmn2YZmE4OMd/E+j3nAOnzlylfEuMc0B93bEnNI0wYGGkj6W7
tDsLWcbhxG+xvvOLbJr51fCzp+iG0AGqgrzPri1IGHxSbyIRW+ZCIqBttzad7zh1
lxU1Ph0FJ8RIIz3KGpfueTSnhk1Ao0nNK/WWsXeGuPLt9x3mCCmWwT4Oc091y+UQ
23FiR3Xb5k+XA+NoHiWTXLNktiGDB+ILp3X7qqKzo9HHiffclN8P8jviMZmPjGpv
Mj/zOgiuOIRj1Rn9LwGfynKLMPqTJKqGgqHWOEyXIGDGzZ+7ecZY5OtmyJXZOfS5
V4F7z4ZsV+ZCWdabe/9IizmxX9h1EJJK0qzU9QfaXh92Ajm3uwXQsAaY9dk4UFed
sgy9ViSpLyAIyqs4k7dEF0YgJi+qD+Y+fai1YC+13hYV2ckasDGckRjQUrZ1CTbr
JV0T61SNcAcyvFw2FMoMQQJrMwSxptgZ/UJ6MmuikTgnHWAhODMBs/4PhDVWD0Ik
Zf32MloCYkPTU6bM6RWVHqwDPF1tu8Gvnzj5wDY2xuYfSrmXW+6cU/EYnJLs6sb4
u3U605SngMpQUQGwcb5qL05gPrrAS/vcUuwl9f1Ih/7xV83AbjPJI31JvVQmRdgC
OcDsnIBo7Fg3WaBReUtYAcWqwBD+CDsvrQ1Ha7GNd5van/0/z8EwzkmE8lgtVTok
XUSMJge3eK1W/dUcAJ9weuZsKUqXw1tQ94oxLULEoFaOAcpUDsTy1BiklfCgsvMv
0k4NzJQHk47Hof+rfgJHWaznPkYrSh/YCfGl7tNSZzUaTNTlVGgWyx6EQVGEMqoU
JQOTgVP8wq4jZxJDZQFpcaps4bwaRJLnbijwWTH6ieT8/3oyOn5bTRsMk8DXhtov
tfL8s1LabwO12upRwgzYnylh2io80IatNaBQXHcSeMLNr0hioJ74gZ94OQZkBy4y
U+2nI3gNI6ECHB0XWlKylEh+Pmjv1EW+YYlfb+n5HVCJCe5ENeistMPRj1tsYqFJ
+SesHoiw7YLcS9EX2iuwDewznwc1DPQHlXtanPOYRelRaKgbfTWmrvwqudeMJEOn
/Ci9ei9II3UWMYrnwW69xgDPmy4AmsJdyx174iL6B9VSLEhpG8zkltrMbUhM40Aj
zjz0enu6QW9yhQVRbN7TdbX8ibXd/kAUKi/dxMTdDZGdGmvE6J2nQnuUSmKb1F7l
yXuOIeIuxtXXbXvF161FRH/AFJC/RbkIjL2Tow3QolVLIB0h0waCAlf+CvWmzZNK
5SJ5+cdaMNdL1h7uiPgI9w==
`pragma protect end_protected
