// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 03:56:35 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MIrRyskgTEMj9jlHKe94ZP/x7n7JazGdqim4YboKbDOHfzI0CPEdWWPxnRxou3z8
bhs7fcm7R5Vr551vuEzCSvWXrDSNjIXuwG28PGKdRC9r+RlcEXgZhR1NxXvzVwfV
x1+hO9r5G8M0tf3s5IBTbVAq2bnmXaajQ/6GlffqknI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18368)
HuV2yzb1WTq2UEfNg3kHzQkPVygc7aW8bdUVx1mDDwdC3eKOW8MmS6PH8WeAnJ2N
du8uHmAp1AWF09Du9C8cud/PjoN4CcBl+PVMNfg8PthDyfecHRLr9rY1L1s9xlRH
er3jnQpWX3GWAJP/dPbW7nVu9KP4nvIN7b7ma0B+gxTb13rcZSiJQubpmOesC3Nm
klcH2fkRRT9MxbYbwk+nkw/LKdjMpM9Rst6Ix/vmWCrjLJVQU5JxvtT2cnUDMRMp
9JOP0cBTuDMWHWHWc4JGbUqdSH0xRygw5gV4Kkm6XRfeONzQz6t+LqcoQfjasAU8
98dPX0HgFc2J4QPWOlMfrvEjU/xo6oc+YCxVHUir3EL1Wg9rcCMTD4oKF6yedrz9
Va2qzdIQQpLs3SnIE1Y2hXIi4AlOveBnqROlSGyu99T9DjYdFbHuXpwWY73lzvU/
Q17wNGpB3RPlADWehyhHeY4+jxhJjVW8UZLz4KlnLEbQHoUee+u6gF1Y+Qucu0wO
5jdxKBvDJCgI6NZ6CYZpoBUIj3PnljZfZvdJrhBDyTyFVIiG3YAIVdHXAmsUNAWc
f+nMl0RoeHi2B7yq86dnxqwNfkuEkG8/Bkx20qCLQ4g3XqZxjUOuVnaWyNARCluG
AqajJvxFV8beBrr8GMqtZ17QK1R3c5QXqBh2281Hei8ZcCNyO8EwLYSIYhquJUSV
ZtjOTxZ8jn6LIxXs9IEp8GrBKZL3TcS5LtEqrKA9uoV55q9pHzOVgG3Q9P7ML7Sd
Zu480O3E8djcIrpzs988S2w/5+5BlZW3dNGMLw30Kqs5JIxJ2mBPZWj1p0HsejiV
ZoTIs96ftv8w6QJBrmDMMtpEiJApFk7od7cJoc7sIhXB3KxIdnm+pPT4TZInEjWW
XsVCIMhntMi18SH/uOceBGm8q/lVVJf2IMjFMX3ns8o2eBaDZNbAo6T6K2Swj4QY
9/kkPh50idPYV5f6RkqiBtiLcwXgvb0hpP7dJsdWS6cs8j2A+9HsJIgozD8FVI8D
ehebMQa8XYU2hxuVQzOaXJfSxp39qQTWI5+5zd325ctPCMUk9OTGqCvCUyWdRFwB
GTY11A5vhAbuRBSvlX5Y7glthuYEq6px3k2WxWvFZ4ApcweOwnedbwrawkfyAU2s
ICsbTnMyLUkVkKX3fk/5kHdRDaVLdS28dcfOEUAFvhKPpePR7ZvDfcOK+M9SiDjc
Fo/xuH3BXzX6sXyHU5NL2PS9RypAchF2DVlDmG5VeDFLRVevl2BZ/PoQ4dqcYRr4
+GdLaNEhlLoX0v1N1ssmdt7b1K2EKYYfmaXxnTstIYq8nMD739xcpbnvyi/oFjf2
Ygc8nQjIimwTAPizuUqmX+98PCSYTil0bqXZqn4yPD/9ORYwa/lu5VfX4VakJhV1
bn8U9FwvrMg+QFnHq0nbI0+9LR4ckEemxMB3dhx5sQ1Xmj4VANsr2/A7LuEcnHIQ
wjRfn2kLNCvalWh5VvIXALRi6LEX35ej7H1Mxx51zJJT2N/ok3wQy02qi3S16Oit
Za8FaX3vLGW2IA3C/birgvRsU2BCpJemIBQ7gqxMHeX2tCyd2vQv22rsS7rvWBlh
cLWzG8aHZgnk6kKoMeouCg/4qHV1Y63pzpnsSoyoAKvbiqYfrrRs2u3i/WZ8v/gF
T+f5MFd66c6UT11Vkiens3xP5h7ZsrE8n9fd1pF82rvpUd15okUc0/NPwB4OM9rh
+zfZ1YskiM3Iblyg/h9Lzyk6OWyl1a5iAgMYZ5eEe64G4fYCC/F4T5z9417TN3GY
+qjG6exR5SH9jSlCqjzi+7Foox+zT1ssrIEyjuFe8GBjCPOcbRQtjMCZPGv+eXwl
rvluqD1FzhPfBuxCqj6c7FlMqxu9OOLfUy+kmnfWhDXs4tf/lNmlzmnB+5xuz/X9
PoLZ4ML6M0DxmhQINFqn5Rr5arfDlaOIqp8LR+d4L1ilf0oHwbL0hejyafJ7qTHl
L3q08kqwAZ9vT9VGiCNDoVq/JViNeXWagRepl7HEYDTsHROaDgGYVVCK8AgIZMFi
Bfk0UFvxy1TScCHb8exou5hIlpjdKpDnptblgj5cLwlNKpoUvOh9J/AHnj5hR8ek
ui4drLBbzeq49L4QGBTe0sDOSeAdxARVxS/Yw0F5249dpz4AbPyI5r84DmXj/Rmx
HB9BiqKOE9e3a2Ciu7zeY4durz9yMdOw+9akcU8zqPaIJPUXRH7CcCjXZ1W5VwS7
GiZuB4MahOKctscBr0pYl1F2HjaFAJngq/uIoIHPeHDMxcAQekBQtXeV5jtTWbAZ
8Jl2cfxTnZgvGU/f69K37zZ57sQRto7OeFMrfa31SbW+MyvOv4OymykLmDvj0Zdq
X8C6Dx4AHOevkJL5BMWKwWgH6aL44p3c48EnaXE6aqARyIHAyxeFZ2IX9/a7ozpU
zYuEJg1VlryWdERhApSJlQ2f20KIRmCuN1zbQISK1hJI2utRiQZOErUC4PeuE+Cv
2Vt4PAKPP6GstBl4h+XBUzM/APQ+Su8EeH5g59cRwyIlTzoxJhpKmapyMj+G3kf2
mcZeWETMGgMQvfM3tcs0/f2USjZMVvC3QFL/dGx63ncDCddjEtw9Vwi3aSuEJkBs
G46LzUFIZsIicZAfcWc3FtKv66jqfLSMHH7x2uXhMPVu8GqLIWZB8rsrmC+HR0xP
dPO55cig7ciTZy1O1re6d/bNvt7aemsmCQio4Her0ZVfHdSyk0+0ZceTBdpdjKZJ
HapXmVXzXOA9tT7RWsLCbhYF3DECKMxA35cvwaMFUM7hJERFIDvu1Y81FXK8uMXF
kh7w5u/ykbK8ywcVd/daztw2ueOmqizLuqbYuOE45gwEpNP/K3dw8PVl37tPWNdn
0A+MnaBh37SMvg5bDDLGqUuJ4HjbWI3Kea4z6wx83lxQ5xbvCH6UJfySBVhiKqrQ
UH6ieMp2pwA546A90LZ+WLmh+7FBijd6jw6aKv7Q84m/SnfDWLSZzMgGgI51OcdV
W+M420XPPHqQORMsSYn1zi0iO68ahj/5i2HJANsDzRcu8xDXsL5zYCNHRk5FtJZo
BNPr7anRU49tdhCb7PPGQwN3TIHila3eC2UHuUDpRuBRTOvhV3dXN9slTVyxb9V4
4hajhqwnnkVYMtIiEkV2JoCMvYkGNuR+p8Q0HuUbFi44m8QoNsD3XLbyYFEBFgxR
Tbsdoyiu0T5DrE/Lmamzufb8IftgvtJp59W6XMShYPH+LXvotRK+hnSg/AGTSBvS
7uAcgGjR9rQNCqAc20VdV+bVycJk+yFM1bgckZcxdMIpWHzTH11ba36RUc0imoj6
o7wy+A2rkN0DmTa7PNkUp73A4X7+Qx1XIxVhrHFMCVT1VoW3TXXisPvVjHJr5D0w
6RZx6Mmk5Meuzxe7qUNoMzNBMLYSyr77hrfc2NOi4DtWdWKuPR4OYevkRktG9ge0
MkzrEJ1hd0hIWT5ZASToFvuPS/fWvRkcKwLRLz//EAPsqYe14EuvKuEpZhLRSG4T
QwCGWLVAzJTGEj0mCSFewmwx3pEa0dfVMfpdvcdoi2HckcAL1NfC5Xe6ZfXtQiSD
c0WFBWArhVC2v2iU0RpCrgnArvTdu446V6FhzE/SVYRSjoePZUWiXDIYQM0z70ww
oE8UwIC8qR6uaSwE8KizpsWp4Ujsdnegiv21QsOdafet3POeYtxfkX87GykXinOI
HnjVQYAkjnwYZ/kbVExtfWXf+JpM78ihCdcUhAMe/C1KSDjZ+8heatW76ezymfKq
1ZqSp1Lmsj749B156dmjSm3AOueJhwVmPJXEi2u/W3qhDqJm0QD20xLL0sevIyyr
62Xs3IARquMpSoU5AVnhCQRohWfjCfOa8XWba33SQdMOjyVlUrWX6C1CsvmbeRQe
emzHyJlfnue2l74UPWPODZ4LvzPF5GnVVG/WR6G7+Up64vPiRFEUk0QxYdwV+wUM
2iqqEFtN8w2Lce2W4chzOkT+EZx/0uLOB7fk8O877x6hZygBVbW902f0lAfrEn29
IiD5jGn3VcsxRB/VF+sx7Wj5EM7o765FJTDeVeTFdfMXnPctxpwyvI7MgwelKnLP
I6iE7MpMcHTOe0InTGCG0eT0prkYBSq8EMkTiYA6Dv9NuYAQ4eAMRq9aYw5VsFjG
PL4Y921Zy/1Jlmwmr9zsm/OnQ+gjRjigsdC0fHsZZZ/5W6H72WLab/YmfjlaREYy
cM8TDHNf02R+MnEz8Pnq3ibe+557u7FDQ9pq7gNsMktURk2etdx1euiYeeWDsTcp
6FVm1YU4pXguE2a771WkFZdY4bEHP1piCkO/VkV35QO0bAEQ1+M5Q/pAjtXG27oP
5G69aksA9xgtZHKLp4uqpv25hazl/RrRx84jhgZmsCWF1dYoIZEf/eh94cCDcAZy
zSiWDM6mPj/lCpFNdXjUOn7poCykMXyTrz+AoVpOophnN9QSYfG5ypYcl1kFEDB6
VjfY+whk5VzP2jj3Cb0EzzkJ7MPiGore0CHqSik4nWlfDuc5VMB4QAOpPkzBiX6K
4Al2DVGfe7KXU1AwP6Fd8Esf8ZqxFUtXl84K+umma4Tv9cpPxSVl3jJGZNBqdbbE
jVRXasQQDCBL4VMfpXzEjMUXygmj+S3iXtw0C+efHzIQq+gMDIgCI4ClKk4t8hRQ
f/PQwoN2ethSDXVrTH82W6amSw0EioAJVqgy8g4BJk1seQUXt5Y+srFzSBf+aqMO
vAQe0GutaPWlb7rvj/hYiYfzWd4xCyDtwW9USx9q2AgquOiQMt9L2ns/r24eXrUk
FLQ3ZdG2hss03IyTuykfCyC4KoavO3dQqYajlScaL1fLadO4rK4bxylrTxusCj6V
RGoxgV3CQijxnz7F5Yh+FVjurYDmzjwEcvBazfHXr29OnH/rHSdNzVBjKmEgj2Hx
DqkIvWZyiS3PDq0DcvW4QWpbTcbfYt7MAtiyYe5604QEasThV3UATnXWqu7SMPI0
++t6vJrVBgmtFBJHbEw/K4dH2lXJ67IePep5fdgHLAISPtdQlzvzX6RatwEaa/A/
mOoN6ECIZx8qGW603jYtTZesyRpq6khsHfq1xgouZeCmpPAqRuY4Lrcs0IdYmAnH
pc2iFrpl9JgHnBmi8+3809Ity8IsmrqhiM3UdKYhQnds4+6XRiHc9/8a72JWbLoJ
4vzylsspFhCfPnGsj4v/sDSnv8glHVzdc2mnnOX0z/cPWfXYscMDQ8966l8jHsJ/
RA5HKJQRA05IdoVD0SeXhGs5yEQi+nPSvp/Pk1838ClvRgRRbBqR/egsxAnMyr2B
ZPUteQog6TcdeULkDuGKAkvpGCnN8cz9E0vVvKW61+6PrALnlsn773K6BDfja+S4
uyfSBdv9OHzu4RGlr5UhnwoHwsrINDqGuxYaCMYHVx+Evj9PZfU7gopJpXwRhuJi
J6O0ilv4Me4MWsWMYeC78eBcL4coLaSiwAfVMrwRFQfQ9yRNS0QlCW18GaUBIoKk
9qRcTWSAan/0oykYSW5FbQHcnsNfAedttNlLcD51XXhpO950BrBu8QHkm7wGJ3iM
JwjmKJzui/aU429ifwZXeeAF+g2EeGnn60exoS00Zoe0L/tW7CsQNIp841WOZMbs
5D37pb6OP8Q515NO2vkdVLtctGk4iBwM2ZtAzttrqenGQzqGDVdyftg4+1WsADn+
OxhJSslaV/dQASP0QJpIffsoq1FSi8lUecnDwEceOA23owTSEei9uK+ERDLNSUli
lJM+7MVpTXMC6sM7jPVVKwbrKd8Y6qzOxwNMy5Q10FmrKkgvmrbu1w6r5yJ16ZOa
r3dm4KG9CVWce2gyX7KWOADGNGQHpahX++CD8tJ+0tOYG7yccp5+EFTtNY/3QyB5
0aQsG7738+jhgafBOvKxdgfCwO4GPtsd4tgQ/sd73nHHg5IdMvmkOQnV+k9h5WV/
rZrksZY+hNWuytV0x8Uf1cN+dC+EDKP2iUoScKDiSfcntRmpXY2r984rxfFz2k28
CU0KPi0XpcDSJ4BszXtnU4b/Wv7nF3PraoQA3fTmMbqFqscyUdPSyh9x1Fw1nG5I
ndBoKcGdzdTeQYZkTSdFbwk6OntoreTlaJrkZHz7SlJTdAvBnXR9yo529ZyJdJ4B
Ao0T/ajnbgJslzHd++sSBkKVdL54onRaF0VHtSmHZyHLDCKfqUjF/bZ7Bn/Amr9/
s+iKPooV9mNfmcfX8TjDsJ6Veh2VAf3LFCIks8psnL/SkRGCbRJlKH5AwnzhKmKC
qksq+R+KeU7ctd5DPmJlUtEEV0kgkf3fWlgmJYm0Ip0lEmHt1Y0h3t+miHGs5b/r
cDXJWwJdVGxQcY2kWwi/HMaEzRv3FiJZSMcSO/V3V8By8kbGzzgeRLgnW9XuJUuf
ggz5dKUwGJNbf/P0sR9lX7T1rl+00HbHJgHSDoIIoqTmH6MI0yyh0Y/OM/NSa8FI
gAseenYFH/p8h5Cq0EtIDAjj4QxCAEZxxtEX0VSdBqfVhphUax6mvRroSOBzBhOV
xMdhPZOmRxcvnpgBSNy5Fy9uDPan3CWPfJ7u5rfvsWywjl7PkrYW9hWH4n2dfupv
bkOS34AL8bCqiurP22N1r/yJNSgeNK0n7xgo/mWqzaBnm2zv3zumgLxQc1uKWFUj
dMf1GV4/c67euxZKQBr1wRbYunz5u4vxVtJEOd+5Y6/BNX8O8zoNnymwrtg5MTmh
11RVj6jPifkvgn1KYUoddLL9nlPbsBS6Xv3IYrlwcamw2SAuGsmnkArI4Ajb8H1H
jfaLhFDkUgSfyzYVREB110a6Uy5zPEbbO7izeD0BwmDV6QWguyyLPl8Fm6ZvQwLh
E6mTBvB7db9rJFJTM/G0KPxGA4wtU/XSaYuWYdsuAGa2nknubFKwCShRSen7Rx/M
/J5d24cj7FnVZykQJGfdEFh+Gifn+Grdilj9HSJSIrLk9K7V2N8HT6cynZNwNYbF
ZydzdRpl9T54B4w9XYFsHaT3UDkEXJDSvVochbjvwi12ds0JAhgq60Jaj+749KfO
DsjKs1VNukOLvLXDDT7ZAcudGwNwa0QYiumqCXEIWppEaGlYSf7sIur143QTrJHY
5mGTVZja+4CSrzlwFseb1B/h5RDC7Lc7UcU7MDAniTcBndZ35CtqZbdb5NlGCXnz
PIMoxTVATbxfhCHTL2WS+tkFLhV0YnvQ6/T4RLH2Aq7IznCX4WZCM7hLMU/vYS+E
XHE0XiBGb5xlgZWtrzU/rqJmeC1kcpWFv1bMISzyBV7zGZRtCOc0iqla4RfMmPXr
gxVljbBr0z2Uk6jtI+i5mlrVC1qJJTZyMpKXyVqnCD3jE/KJMcOgM42LvIDV/qQ2
CJSEzbpi+czsNClytwhtORXhOVt1OsFAfQ3rWdvAPFLxD3OI1kOx4TKUNPx21CwS
VedwJPlKdgqFsNqSs+upWcZqhtPf5m1DC2/0Doby6ZRPZfAZCikc2xzWof7cAhtE
54VJiR4lPLUmOz6r57UA2C22L6KJrT1M4KLBNs9gxrGyZM+8Xjh+Y6uvsw6rcIxE
8oLYTqiYfe1tTvRqbrcBgqfEm/hPI0x3sKlxTOgC2JVpBep/4WtL201sBPdyhMjG
9LqKjw55khpYSKbcR/Tmdrq/zsAUAiWL1WlkashPgJIBCNjywiWKqq/0kV8UlzkN
8JSNWaZ94sXMb5tEpjXOB3yWh2wCbAteIoOd7j5/guxZf8H+Cwg3wiQvcI/JOJ/h
GX57e5GjWxlrJ4GHD+zWmfwaA73AiNbu/pcgfoW+vd3xQH7MrvU1T+/Dx/zm63bl
LpBR60VAt/Reg008UWRJgTuuzvgKK9cdRGrnODYuwYKgpttvpK6sqDKtuOseivqE
i+1HdN6RP64T8zrNPtrGTM/HCQGvCY3fPJgcv3C/tgEVs+nDfXp4L9Vnn96VAp3/
5DaUTwgfxHQ9xMMhAEOb5lVUUgkKTNyPn73MbEzPHTmvvL0RoRBnAnu0s1oKvbCW
JKIApiez3sZMugu4s2gA9aOihnOJeA/J7dz7g336wJa2QcuR1fWvg8cN3Ynd0KI1
5gL5yETLSZoIo2IPTWW8oHTr/Xrq1CBOXRdiG0t9DN5WRyIkxlUKWYZDED57aqUH
lQZTv+/P0XhMKi8bO/boRf19cWOBhj6n1QBo+NOiPdGpq6rdIGMKCZ4WX46kV7RH
oFicY4zjVx+nuHA4v9R+f5k8DM78QYH/5f9J4uEZwt2AbeGVsM0YfqEnSSPDfSww
Q3yMZ3Zio7ajfPFFmWUPOc0psUG9vO5HMXYhbIYz9QBi8+Dfffr1xTv1NtNgsAKL
lULzzVrIkIftizZN6/2HbNWJsCSNPtsdSMDFm1KkiqMl8gzYgKnV4Y1iNAdLLKaQ
7egNPfktUuRWPPYjf18keMBpG5daZhpDuMQdzbaSHZRL8A17hvfHNb4hCZ7Jw24y
fJFbA7iaTOW+k6CU3txZ/Hz42hJb+z5SK0Su4H5Oy3sMFWryA984kJMyeKij8Z0w
I4umNT1rsRjooQM1FK468WO/vbV06pBGUBXy8hS4OYCS9DNWZq3d75mhySjbNitM
tOUpjQdCj9T1uARqLS+k48zoZ2NekfD1G5mDlR8KZG2T0XyjY+EpNY2UHx6iLnPj
bgDPx/2BL/Hux1q4cMnNyG+GdHyUhHlsBfPm71XAKCf0x8LVv5Aa5wYyxnFWh8As
PNKJUnOgyUagw54gzVMWY+jI5VnFWkkbNYqUf99ZP0GviQcK+Y4hF55j2xc+TJMr
vz5Ioa+/J04ytG9ZUizl2QFffTIAo6+UIPk7pM8ImEh4HDKyOWc8LQhth5ykYWX/
ggsGxohA76FNJYpUZv0UKKtD5n+tebnHKcEjgH5nipyW6rlx85WqUlasHpjRgc4/
XBWez39YC3ksAZvPZUAcqEUqojGMj+RVHCwH2RUiDxtv2TD//GMzXRd1r/EoGJhC
TRNq6WQDGHZcYut5S5qjuUzptaWeGYi4KX4TBiLif5Ks6E9uWn9hNmc4wtedGiCg
U2xFKquSI5y0iaZMrCDt9Tg7Q6CZLZK5WO/0Aj6iKloJWVg/XpItvtuI5Dao4pWf
mhdazLtnjCIys+RVe56Jj4ynOE2E0FgaqYaOQ/dNrUo3FcxEEZFniraVz4W/S2XI
ze1DlQJOkDY+vC5Lwy0H31x89vroTrq9LibOTDOl6G/qnUEHsUHmJjB27hbJlyRz
ULzGqIfiZEfhWZSf6YcKpRIPKnREZc2GQOpTTd5OdTlgJDnXRg/xvY5kEgiVzvZw
s5t7KK+2JKBaJXRizRMeBaB9v1O/1gaUJNLXeNFhk6AqI4GGbk0jwUYOOpGf7nFk
TzYEBHKuAF4qzL8rJyUhorX/6xV6C3e4kLCa0/D2U314TjWd1sqOKBo7fdrP/Yvh
4gzTPM/GPB2jiZIf0nuke2y0onyCrn5iZaH4E6cFNwawJiLlwvTCPyJUrhGcyJVl
VyX3YOeADDQqv/iFAvY3VNhVVrAVKW35OBGbsuzP3V+fpGKAjmXUmEK017iM1cI7
gcMSySQhBXvDPz8WHltikwkBLvQnasm+G/bseqcULrpFK08RBDWycAPT1SQVhESM
W5YY5Xy6m0WiYq0vM6XDuRTkmiX19qmuwWC3E+BjXQEut0uldKEWcvA+FtZFdsbs
WQrx5zbhqtn4qvI88ffRNpMBRk2d70wOgWg+xxjCKi22ZWjK+yYKrUI1Z94T/MFK
sWxThQzrHyE0A6L/yo1mmKVEKXSIHSayV6thXrGWPvkfTZ1lhxUReQR3vRA6/O7q
IJZ/pEGsSHgmBVZ61H6lKU68wFEcIBATPI3TO59O+juCi6XVH05MlSCKA4ZWCEIf
Vv3uPn0e+baZTSAbL4Tik4m85rTUVnOEXjE2SCPsE3nlEl/nGuUobhXgafc9IHjA
ybyTht93T2NyJiLClWnpIUXM7TiPy665y8WjGVMH6u4C5GSyAU4PobzC9qIVF3Je
0fPY8K8nPCYiBvBRX91vGvwFfvAqJYsMOMONIqan9e4/W1cFDmCivW1ziEc9iC2A
N2TwBhj0xxJKJDbl2hyvxBss27HTgKZ7c/n/njYguxLCD3nflJWiguD/MEsv0/VX
UMjIBKrCpheCraje1ezz+1Do7hpmShrafgliXODb5tmIjKQbTP7jnOAsKkw3c5wK
VZssnaAul/TjPMsdM7bSKiVmF2w3kiYSJP4WQGypOINv1GJ2EwieTM89K1kwLbFN
k8HDgMmOMBjQ/yNOeS2I4YKhK1fMRr+O5Kvbr86WQwGGuceTN9NJ87YHR2ysA2hU
AHhiXi6uq+sBDDdDiMaaDbHX9V/5dLlqaA5+WL6R1g71n1Qy9ramAjGj5LFaAsDj
ayed58dN+ekXHqJZndkBKdod4Y/LO+fKqv37qw/ekMuhBCQc5mQ4sJvjSEU6MuJs
ubMFyMljIxQo/ZxLmNR4QUHb1cRl5h+3ILpgbJErSJKk8D+l6WOt9An8RUJpZJ6l
0dVVlbImVIVSnYhUG6Y2OXxchwkYLNCD0b1+qSS61PR5GoEITfp4vssoTgvX1RgE
LwW1ibIOvAu+qIxMZ6J/Eu5sHXlB//jCz3J50jhfRjWKWBGu26LNscWNdNKN3UFW
yNhs+RNhEyVqCw9zrrOVnI9kiTll0nx3P+ORTrYg36cKTwbYHUO824vA4g6rVP/p
Gd4Zyl7aKw7ZqOa6rNefv248JzJN3NBQB9S1gFU+DPnP0EytDi5ZvMbbFEh3WE+U
cWPadP0EtZxvK+nGpD6/APUESk+gluyMWh6/vh2Mf+i1DcRfkxATVl2iUfzxIroQ
peGr2mxM2dL60R7CCnxCubDjHLXgDt0ybTAcJ66QpH65UDJzxJshW/vKVoY/i4Pl
BRPaMBqw9cughupT4BEXDN+CATutUodpS2oTbqNAbkMyNmR9gukrGUTw65rmTB6d
cSmFNOZ9KrrCeEDuV5E13V/m1Jid3cBC4sHeFRN8MiE0VMIida0Wqzp5xwHQeJgA
ezSrMwYV9EXowko7zLKvr0IXuJ4qhC+oRO9LduQeN7omZGw6Uz2JbcRw8nDhToj0
45bep7Swop48mtPVTjcjsiQJeme0yqvCqC2orQgu5kWTu0CSQfklaMnvQiJAIxy1
W9UxeegGXR69B45xSl4cpsrBGRRGTThu2QFRJBejcowM0CRQtH3nF1RZg7yrDhIi
bKySe+Y4gfVTRm8ObJ9m2Ocrimvx18WqyWqTFgbOp3ly3uJgjQDr+0RhBVIRY8bs
uhaqol0LLoG/tv9tqrdO8YsNfJ/Sxq6xrJuNpAV3x5F83JiQZma4coSHOwHIJCYH
DT7qjwc3bwYKwxIc0DQsIsa9zxC1BFQDQZgOLmKM4df2t4WaJ/aGAJVITMqv5No1
MXcvh31e2AdD5gY/37XVLbnlGwyoKmnYg8r1py5SErpIMIHjYAKtKE6Qtc/rpnJr
ljigsnV+07VGsa14+joH/afhd/4li9wyNcx5st/j844/tn2WqnHi/HZzwyRAmplW
pFnEY+zLfHPgY16VyjG7dUHrZjYiJiYoK8tR7Z7Ht/jBkZM8W0biWnxA8vID76ld
gM0FJjPisaL6oE7F4H19M3dbslBAcmAyk1LQ4k4fRrXX5OWoTm407dgLLdvoexBY
Crm32QPvMYWeoD3ufTFl/+0O4OmAztLzuw26R2y80n44WYcCeoh9YntguFBkfnLj
FjU5LxqAyUw31LMwYdhFfJCh96ku4EsWn4mkKa2AXcAfeaS3ZEIdAO5b3tyUNKKb
pKDixr/R5POmUDteSa5rcMBXshWL/VbgJKdQgBY7+HkJZUNOQzxCQNHJlGwkKj83
BikNeMU+LjM/bD+Qxra6bDST5YpB4sYjaBljb4gqVBYbY0spax9FAYFMFPe5JbEP
wAQgpsaXNFygZqxkP4fSdnzbkR1abjG/yAMkk3/16OQImZ6+jxLS99VP1ciyIzmm
APTglJ9NunGxSPG6hYBHm9bN3oTKN/hSVYtsPYKJuRMtNOh+JHSSICwjXnfIQW0T
H4cRj9mIjrVfMZQRE76Wv8lE+QwlRe2GHB0OtylAvBSJmhUBmqxF55tx04J1gXbY
yA85KH7lh5vxD6SvVi5sXJ9o+2nBURqvFYhpVRSfZVgfdUzxev49ciBCZR1xg+87
20mOylGAiExwQ7nIMxSMncJHUo2agg5qE9RmQlU/HivnRuy8Qo0Fw2Axhd3TS4vU
TqHNg3nH+DS5xtR1mbMHzsCoYi6+tfbzO5Cb9z6OCYILx27fjc6EY6li6nU9uTlD
uPV24WYm5KEQeUG5WIXbn85FaEwii+ynPYrBRe7yL2Tnl4ZHc2JF7Aj0xd1TX6ju
CSvw12jPADnq91b51kPCy4T5XF8mc76NA5p8JHbq3ns6SY//saNjwxYdOcPTWfiI
dzib1PlBipBGj44nvv5RXyN9Kc6PFSnmEpbDa3I3FU21KIoAuZpGFenApDTSfmNj
WDXQi6E38WTIC8HWLRJ6akyEk++86mDAopw/bPQ7aaU4TZLGAUXfzPTU3C8UulXM
ZP0H4GijlswDHTue5fWEXSRamsJOT845nT41fxcEuk7gABz0T2n1Nf6djsi6fiye
+R8Kf2tUqyrCpQYNQO3aryARmSpaJZDeDJcgTC0S6hXkx54bA+pw/kJlDRDNKJ3S
atYIjwXO0E9Zu8HPNSBFGY6JbUykIIoRvqtlZzJeFGrG1XPb+qujwcjhETh9oOeT
Dw3QTqmR0m0pVTreM6l1QZ5RrXXP9VP9w+6UfG4BlDEF0n5qHmLISw4zP7En0MgB
IkWCeQVJHE1l6BxnEge9UnfHbcUWEWBgRjDczijyMncBrG63NQDZIFWHFrqB3xHj
5AAsSLYRWeHodQD7hfMCZ06WY10jyxaBe5iDptwiX+bMTo8ABo3lb2T37GCJ8BiH
iYH5trZt6VlHmjaV0oF7z3hGzPRt3JJD7ZpZZk9Gjcxa+EkDS9EusuMq0yBBNzKY
tXviWvNERkt2MFWCpAi5FcCPRxqx9B6QmQz4Fo/EIjGyKRhLA5WiFsWftXhaDX5n
0xqDlD2uZc2XoXDGZC0lu3+7Wf7ANdaZUplhNorVAcUHYlIB6fcoNPWTLbfopqGA
nmiuFrHJt6WnqsO7EFPM4lHZMOE0v7XSndDsWlr5XLt/MwHSatrWcQtF/+IHroAy
cqprIZ9hRAipyeGZPqX1lyDqP2aZYBUYmeIYiC+fmIFJYnqO/YfiYMrk28sOHM4h
POG4+xOusiNmL1q/XC7N5Cdy2/N0r4eQIE4VTPvL1/vfoOq98EalRIrq+GVLYDVd
DtAthjssQ582DPjzmpgSUrWkJgM6XU9CxuSdN8HEOQ15H4hAaT4fp1DQcrRTJg2S
TDGmTFfR0DTaoOEWPkYWpF8C2GUaJKStfELtQWLF8gSS9gytuqqqtb7r68xpWa6X
2J3OPO6cMGS1ZUc1EjJhg+fd8K/u+OMl3tm9PWiVeol9bR0EzDFRk8joWY+1OmSX
bTpwR4qMrb5sJwK96ktSm+Sy0iihxjLYgh0/Z0kCKIdo5rEg+OSklZmCRAu/HjWu
K/GQ9S61qMyZ/i8STcqCUT3SkeMX38xuVEh+7Ld/shOstsF5kRxiUH9z/Bne+2Jj
LqWQTP7JDg1vIPcSruPsfBJSyKdzK4YGXac3P+XIoaroMz9vTDUoUiHhbcMQdX6V
6wwIvv/Qdm2/h1do7Q8x0dYYXF9OO4OINWEXN3igpRi0LCSTC3w5Q4w3PDoeQci2
c8//n4Y3uUWa/n1DUAFh/F1oQaruvE78ySnnybDUlAd3+x5KkjvED7SGMcOTKHZa
XFVBvWm7+9qYs9iy0tE3lkrxaax1whq2E+sg+5aQxr8uzPvFh1WB8cjnd3gZbLSg
8WqYaIFFrDrdCZfUnoIYxdTxJs7CmH51/I4g36CkJqX4d12ZAmwEgXjWEYa0Nsss
F9AqJLFv298hcd2tMHLx+WUuG1plGeAD9DgcbndaIwHzxocXMIW49dCMHQ9jaGE+
oEnFbv+UFZJXko8I1zLSiEMyd+580/R7VeDQKLO8hV/e8Ih4KPHEFBzat8BIhS9a
WZOMOKdQ0uWDFx/Suxkh4DpwuBydVUhQFaEm12kvEUdSbfSexjI9G6+vm+x9Nh7h
qKNX8jjcNVECJ7IFM+YONkXGD6atg5WkDiK7z2NSdtno870GCWOHQUVWlZ43/Twm
pbbEMe2cI9SiAKKYZBo6UkR6L7TaF5rqMTa4Hgno9/I27l1ljxLyKy2SPEa9NBA2
wIqeE/SiZ1AHF2dwKFWQ5NyBXKtSdzZNaVSMXJ1o3i6nuHEJB2+VvK5OlYMdKnav
Bj0Vg/zhG/8yEjopPGSIraIoZIBFfqOlwYL/99Ky0ZtHn92yJOU8BRQp8O8sVZs7
VqIVgrNL/7r/oEUAJUo3cv3/V8PjHH+rteIZ5byx7zQ80PHxMqdBN0WuCHifFDS2
tmNnAw5/RkUH+TCTrvq2CaFFVFAcs5hBmFDcUxKS3ar4nMI5fGSMDbZC2MyKvSto
QbtN4SyxJhVEoTOcuqLg4F6DbpX6QCKPTkBQOvJRUMCZ8TgkhM+tTr8IwOzJCtAc
UErcTxNrFC+SqaryGRD5rCVgCzCZ54cbJ/EaVjEu5NToOJ4xAn28s+nY93tri/o1
jkhBxCtGB/dTpcFcJ5cZ35B+Er+J28UeF1am5Wj80KByhxEHbqrESQkcPNVMd64H
DgVWZDSEf1qqshX1iBpq9w82lQTFlZLvQkINQBj3doiZT9ZGeiO0Kb9DeeZ221xY
P4MP5dnNvkYRM8MFr03YRzBFEcYOWskM4Pf4SuFbsVzY4TFqQZsZ0d16aHlseXA1
19U0nJhYs6AVyx2+72qjtYFb7vm9ScjA6fPOBPYOo6VJeFdAGfshtz3pVx4NDjBX
tKMYBgGIHcMQNtjgmwG1tlsb2AX7DLKcpCQN9zi/FPXghuy38309oqxdn1E+OKkX
jNgheTjY8xLxAzFArL2H5JX5Xz67M0TM9zdefdqgPRu/q363BRBxh9b+ETkA7/pl
w0suuGgcCLzz0N35HzhHMyDsBBD5ZQjGXA2E0+i1piT270wPejiFOb8aismOQftM
byIbevkP9i+1Mvhw2cDz6FlOLxucVJzj71gSyCEZGNrauYRC3bY1lBjgHD/8epO8
3rNKANYOHWLbyxhVu4IfQGyYWfwPyN/mxTWDHcCAm1N+eSoWv4eKq0ktfXUEgDoD
pq3arDg3IVZEJJ8atvqOtkz9Olgg3P2oHjt5C5bjYv+OEewx6Rpzmdpxepzxcppv
yZ/KDfszeOQea3ZRWNWJiyZxNyB+qhsj6hXdDhIdA6NQ4ZPsCAUWe6f4tfMoVtdv
/PGXZ9HvaHoDIoq1tRP3KWXrVF5UCPsMEPSPDakpLLfDjAVsNic5h2vyW5G9O88E
4iYpKj5iTIcPLiD4OLmHn5lC8NTMYNFl5PSMj87Ex2w2J6q04TvqWCFS41OJrwgg
4NYNqRuvf3ymbvRNe/HmsCYFMDnh2XO4J+NKseh++VNmNdqcIwE8wBc2BamwY8hr
9mYhGDlXqXp3rbznnMpN16V7OfQvRIP0ByK4xGpHo3kXeyVyV84/J+FKJ8STuPkc
qnr6EwcpCz8p1usJ48LC8sZCWwQ0Svd0dt3a2PWb3XtcEVTGISHFogZzIyGfpLui
VgPfK6C0WijuL2ezUm8zvoahteBhRMUuwWDKkXz0YcSqh/VbjECRPw4RwIdWEPAx
zLaKtBQukDfpLXQ0fqt1tz9B1IqezhFoNw3pvv025TneH40YpLPX+03W6VtiwaQG
8/pnjExctmCuohNNjDbMpj0v1QxXnvZ0oI4wzoKXaFECtlPIWVejo4knQ3Y26rxg
gor+2in94oRc0l6G5ulPAFbBEPSEM12Gtf0zbx8tz3hJyIgloeWNpAtJ8T69LqDW
ZtgZtEU52eam5AQMgnHzOQfFoReHRcb8rK7RWQcq424RvaRO4DGNJS+WEn3cr7Te
uPTFrEaTMypcX8cxAenC+uyf1SnKvALteQpuV22ne6oFT61YlB5ziQp5JeiOzd5d
mPrg0wxQbFbe+IW0T/eTYjVzndycuJHXN8fzg/u+iR4BNN+bIacMJplN3DunObxc
/DkH2h8l0V/rJvdx5bz8b6gnLnt6YYlQ+WyquArjDTh2hm0n8MV+WdpJED1++ANZ
TkpE/uhbG3cD1fSdiQqsP/zUWVr2uCzdq3VD5ep+1ucYa0BJv9B9qJfoTig6yS/J
VKCGLdJ/3+FE3nBFOEafDcOFzgaiTHU30d4UWZ79o9iB2SQtdUuySBfhBvtvM1it
Zb14/xeBGR5jui/k7w6BzygCd8D44rUggWMGpABgpcK0pRq45lqkuhDU19sPoUGR
QrobkGZgiwf8SSfs7+bF6PA6U7NZ+Eo911mF0M8e7WRFCvxppu2Sk3hr4+pSHG4k
NiCojGsSpJDzaknb82M9Ptkq6XCXZO58yUtX9CMvZeMVuhAJ9T+ZwRO4X9MASf97
hHcuoY30dwTihY1i4lBhKxrrL4PXS/ytWfO30zNVgbOmkcn0r9P+vb9hjLuhVml1
/mjwUQGDS+OLN0daX5wCH6dwj/rTE6ce+HawoVEUOyvnZRpZrsHrZd5egTdWgG7O
7bXLrvPsnmLtXT9Fg6CdPbeg7JYb5J7JG14kCQzOvKbhQwN+DkyOLIbSsG8mu4K+
gXT6XVBSep/QW+f29BrnvI9fFAUaV2CMjybFW9HbTI5hUIL2tQDCqEbN89G0WMEl
ONgwYGLIWydlXESjLSPbJU6YyfPbebGTjJ5LX8Ha18hzGEM1ekZgQVPPCYZd3a6M
deaw51YmHSaNf5iE/O75q95QGb8+6hCCV7iGUIOO+nFUKbdMJOM+odWL9FBYcl3K
IBWV7VkKeDV+ddoTsBYjKC9DwAkwAWWn6RIXOm9PpEJUGdt54xMuBKImKsGR/ZYG
3hqW7O2asnQEb028hxAKUHb2kvY6hQWSskU2dMpEAZP0bu7kRp13AA81nwIF6D3g
JJpn312qVyHwdLJH42sQjUxKPQce3gubPp6VsTqqlqUkjR12UEhnWbbltw/6PEQx
qNIqJTPdVkivzzpDYiIimlDIWq9HbLUaCTRnfPYfSKNmzQnKsdP0yN5+3TbyQysd
yDhQWtCNmJI63YDamtEAIwLNiKWZ+2lpvvnL/8Fpe3tD2Ovw8fYVfU+ukQhTIpLz
ijja6h5Z6ZIws/zW9/tof07KjEDNLQIUTRPJYmwIbYLO8cQtcmypWM1dZjQW8e6j
TJI4nymVx3D5H3OuC7Qds8Z1iUtULUCi3Hxqrpupf/xZqbhDGwxuPk6IcgeU3tqr
Ay0xh2hZexwsKdzI1c9r77QrUEDqwqNFF5sUhx3SkUTGmsl8NgsoMrqlIXV75Lse
HgXTwUC5VqBapY8OSHdVe2WnokHl7jSbaiuw8+JW/QBOrnzCXSQeZ1gLaWLwbVcw
dDawxb1KiM29MaVWjAp6K75WUUrkar6LTMVBvs3KE7jM9sdzhkhsmE8LGJq7esQQ
ixPumGY2MOnWIAYxkCwaQ6KkiC1IZS9yNg5WphuVhsVb31f/bdPgDxfQhbDzN+3m
EBT/o1WsXxU6112YqIAdgGoVQqt10xclsw8Jj1KPSqWNqJJQ1+Z3GVmC53vLpNjC
OBjzI3oCj3BmzhyTWcy+5yamVffuVvHtsGr7OgOZnUxKQdiLJ6x/bwBiSgXWfCEh
Es8aYaVd2sI5g2/qGeCFBFl6OietyIdh/4ZqVuS6SYOTrwYycnRpHx2OkJYQMmNj
OAL720dLwkVRAfeBWEYg0Sj00GaReM4wIhMbqYSIZlI/k+phaMdwog8hvjBE2OXq
+XK++j4sGtUUed6ME0UMlCzJvsVK+C59Ff54+ouYfci588p39Br9ZiL+TZd1+JmI
QObvZUsXvn6RKRqwY+CfpVqalWVcoW/MPeUoKKGzBJQyVepaQb35ETgOZcw28TMd
R6zTgZQS4+/vdHmODl0aEiKAOiLrq9yNl+1POij+tj1YS/c6iTFIgws2WhcjlmEg
qWhjnkCAfxvjQxAVSCcdA1s/iEyqxQeKnPc0ALf8XFkHgqtSajb43UpoVGWNpMmx
IxMTYiyGPMN1MYmbZKDBiBYy90DdSjGr00m13jpOxSBsJCY3Qo5WZQ3/5sd0dFKW
oBVf/9L4Tl4ADCMpadG4JXvmfp13CBppKZrYUwFQ0+Uer8CKDPkcg2R7KkeTqVlL
7rWwE3atqtFwQede0/nxGgy259GioVTI/8GZWU+Jv24HGOYeUhLNd1NaaLaw9nM/
nT29AR1l4PUR3u489f6cIHV/srvtq6OC6hgvRITrb/3LlVV543KkEaV3Nqpb/K+E
9y/BnQ5DjPd+zdwdariUFdBYlo1r42Si0Py1Eaav6mJg4AR+e8zO0qUw4dvKpT8T
HG/TJoPN2S8EtzblZA+NwSiVI38Ru/QlLtMtrslVPYPphGpzkTMpIkrvOMhA9IgR
C7uAmvhPM4TVqagWCPr7tq31aphnePVOvD9DVFkMa2SMm2HqhJIUsfl437uRxnh+
yCOKoeXhjZ2/yzzOTu6mQK9dkyB+k3EueZKeB0fCblFg0nctwhYmF2NSR1FFeRpQ
HRNOxkyUKTd4FN7hNbNhRNVwNv+Kgty3Xnk4OYc03sBFLd/7lUg+PK+K107PNOKD
A7DX1JgjDyyVpaaxKkPMFe6kWd0i8UpMDEPk0LDa62gmc8X5H1ms5HHD/1MeHk75
pozQJT4BUwG7e0qhqZjVC1K7ggMasMzAnQVR2B57E1idbyMuL2MKrKvHLTfRH7lz
pK9EF0KT82h+nZ+hJa10Oc3Ypci0M+t2uMrJCNVILM3p4iIW7uz06MSFh9uCJrl4
6XO2YBioXu8zBs4r1ukH2PqwIafn0PGlA74moqS5wqcgF2pb1fa8h5MH0KpxWLzv
BN+UOuE6ERzdJZFDv01OSvuyqb0FsfBENFengrTBzUAwaOzsaj0P6Bpm4tSStvxD
ZbB6NIhBChQyerjZl0WGrWlCWQnW111+qcMZ1p2WEtvDQttSd06YvJvxZn7LZuUg
9J6tigUnYhWZ6YBwh9ST8PSuUdMW96fIddYx3bHRxjhS0ehbiw4kr5q0F8op+Ws3
veKWFiuMsmk/M1aUe+L1EXIKUwtohyitGxIvcuWM1iy2Kq9q4m3iwLW4ZakXBc8M
xV1p2lqsu5I40Cb6g+pFhsToHBAyGIsMm8kYifT9WFIEMaKNiiIzefluGcmIN+ye
4DtYs/gUwtlW87lKqsmwjkSu6TBLVWOttehTsrwY9XtT1qDQGGY40PHHpOybrwaP
J4DUo5KNUPzanmproHzBqJ5JdopWYm9gD+j/tzAJ/6mfdT48YFqEwQtNmnmTUWjN
b711H1pPKOcUZmZqg5CSBJzy9ehrKyvO0ZdROH685Utajg7pomLMgC2fAfyDsLrK
PrJESKmJVoEtFJWq4beQ/aRR5tVeNg+1v6XB73pX3yER963RI47Ky0y7wPSWDX39
5cbJ7+omAq6rpY/OmY4DHSVAgrQx2mibl9xNFE8uvRjESI16oaoYvEBhU9dj1FXc
BW/tbUiECQbhIJZd9yRvTJta3ulxb5fhESPcRdbE/Ih4dsuaxMQf4GfPn3d5QBIr
ZOR0Z7d26UGg9YOrvKz/W66yh3NMYvxwXQGcJvvUN9zgTFO3ejnfhDm7WszpZTsl
bSickmhUvlagoVo4rbqFniiCifLuppn9NhhO2AMKSNJhbg9AO49QlduJD/wOy0Va
yU9HBVTHXdYlpigBzi8DnUbIXCk8oIWAsQwHt2M0S+SQMtbQcG5SQXF8Rq5W3vKY
SBQPzOnaWhShFx1uJG4qYXvChXSy/+9HLdrXDpRO2Co0U7RVlXM/G0h0Pzfm2VAe
3Vbf+7Ys8wuQrkQd79NeAbEIduD6QwkFa69K10yug7fxAdG2fXkEkz+wloATz9Qj
ykSDFVSYVa7k227pPGb6EOF3ugKQvLeMfZifaxAvJXr+9bn3iuvDsCBhiht9Y4jI
ZvUm3O3oXLgLLYqW2DRhcgsH26KIaEV6KasxtGhNpVDvY0p2nKu+mA0wq4XGBmL7
ZpKTBAvYjM5Qedn748eGrU2BEJ20ckBpYDjVqs7hMD6ilMMIjzS6Gm47JkhEZgV3
8qeQiY9vxVUW45hV6c3sG9gu4kaC2nfqxRGiLy0m30f7gyU9XaZ0y623xtEWAWdG
IOE9FlCBkjgz5XeaIBg1rAHIsovlrQeeacbuNajDf0fyIn4e2mAQvSNgmvoAEeTA
zX+UNto/oaFJMkl/7HIvYGuZDV6m1UFW/UcLarVU9l5kb+NszfCMdj1B1CPqMUli
j7lbFD5tYYe1G4VUs+WMan1vUgmMi52jIJv9rqJy151Ky/S6NFpaknCpq5AiDAP2
5agd/DMTyL8bQLbKZFK9oqOjDuoM1DYJG11kqDE+FQeuLDVbGsui3MkPB5ySTpLo
/0nAINApIqPg+hSbcSc9QXWaRfoiy5sMIt21LmCAXzRdMQTbgRsIzta4cjrogPmN
+T9aCafaYXxGDNzXwa2vFr7jZOry3KWBMvIjs2dixgqf/bC5tksGkyppWXDPPZAM
FFsZqrK/phNAS2VwPVzvVrHcxZ/rSExMQ7vDMvMr2wsN7jobDsmf+eogVIe6aqvx
P/DnNk9128mvvnsZeLYbqIg9tZv1sQ/0+r9nm7iSx02mqIZJppV+AnM+OshRvVza
b1u6EBhRo/UriVZ13x0cJ6M4WOM6njt37LXb/pEXHGqgRrKSG73lxNrRzaYjcglm
Vj82Rb9mYYRSYXwnIf7NmmO7EbQdejRzRzmZg1uDUNMb0naDqrE+F6Ylb+tBr0kc
ihsVAySBGUO2YiFCWfItaKsOLc3D1agjBR2x7rAHAFiNPtQ+JNuphhZ+40RVd3aq
x6tbgNmlPWYvdgGUBFsfXrKvBKOt7lD1hJaggblCsF8mHQDLYscLauVUtijHhPNN
dh0Cqo+mKihb5MhlIbjlPOS68SPISh9S/E/RnbQuHyVC0A7uSxdofOfFxHaovFGb
YFTRmAu/f2+jXho+wzXtnbrJBKooVUISRwGTWCBhH1ohBc8fZIXjt3d11gkT8VOV
Xi82MdRFcZB7qW6ToQtBbwMbwK2aCqaIXn1JUw8/rm0QqZund0PKoFjgtPA4id/9
pgpbPUMtO1cbs4UrC2ASTWDtknnFUlUipJnfbFdo+5qD2T2d6VdvoIiKzzWoPGOE
L6j8IbryDFyLBGcCxeFJmnZoApMjsluQj1PwiwZIJJYSofs0Qssg+tEdMApKJ49T
7Pjc3yEmI6HyKqY+Eq7I7ai4tzmyN2FwY8O1i9TPLZjk7U0WSV8kEgMgAd+23EbM
zX04WUlldExPeoMVTllwm2+iB6YQKvuaQX+TA1ofCSQ3wqzkgtQx/0A13sqf/TC8
xIR4V6SmpkBmv+DEyGSGnHeZ/AXRVuPY7N9PQLH4aUyCb6IUMyK0cjpve71H9rkT
d+7iGmYjJvm664lUHIcvL4RN81gdjRtYn4QgRslA4tnn50it2zNjTPV/i5x8CwRR
7/sUVVZuBlCMneSKtJm2052N+v7oT2Y36ulpmv0qK8szDPMfzFqQhxIVDf7zSuNp
2HZj9ArqIIFu2EtBPw9SFWNZvRMMiMLQREPVK7oITurQbZEs0vG7ryS9baY2NWfq
2ZoFPHcfub47CkiSxfBAHvyK/+8d2maiZmvDnT5Exh6HQWoImkRa2Dl9jSmpGSzC
JsTgVwW41qfoTUXxJa2gOKiAPCJdRbE5Wu4Vqq7m2LOVzh8cJJiz773IFVe8fC0V
xU+O+6ZqM1JhtSfl1Am0ulcflJfbc5M8pT+dWGKsuPriWlrEvqkw/FH+65Gd5F6H
AdEkRQ0IRzZI/JEu6juSGgUzXXoofLG2dp+FP7P1qdaFz2pgo1K496zH927nyd1d
P4bYY7v0ztmVDpj21ydYxr6X+aLzUOetaxb8bCWwE1Z8yw3HTf1FxEKshak7hyqG
/232rTcb8Jnt1tuzoTjm36OX2I8pr77urh9jr85fUQKzehMT5bcuDSR2DomAEJiD
RyUC+XgxV3qFa+DA14LJKpbY8Y/5IVf5gxcF7lbSNBB4n9P9s7QNqpWzg5akr65t
TQvrxpymDUXO531SSLBVkAxkyIemS8ni3DDK/YRIBnECRjseH/fePK2048LHY5fE
9mOcNr8IV/uOn93aSjlvy1h/HmA36ab0nBDxtfI0TQKsaOM9OyuojZ34rjQMt/NR
zmPQ6/mIDJo07qv2+TSqzpgH02PvIGuLCvJRRMMKbKgitGYQZMkcln7mwUorx6sB
s7nPeeTA8aJGOfh6zldm0i2KPqe3G6jKmdy35Re2Hr1o6PTxkn/Mp/2Azhyl/f0k
45G1kDMy/69ukqyl4sOylBxi/BE3SY+vqwWinWTsrmlUNmX9ObTT0/bTeL6JSvWL
lMByZxYIeHzyU/lnpxHgBpDVfrAquRaTcRmaw5KhmWp7Of2E3e7oJZ6bM+2XmNDP
Z1eI2O+SpZKSdLPfzYdRtsqh7g17cCvnLQlq9bpYjzhDWhth5zQlzDvUSkSBjmz8
Is6Ugos8uEljmsZzQimIqs6Utw9hnx9roAT2V3T2y9g00VgmMSGFnTOy0DSDlEfA
dJWCLGbhwndgZCE5gKX5hJb8kG2JlQniC5zsBtH8P4F+LDwum7ZIgh3Bw8lfjK//
tDH7VqHUPXSKj2R1iqYxKabmx/3jJeRrFOjwiN+a1oehLPynK0Xom9/ryMsDnTKK
CFfqIckZ41QvqZUlB8EN8ZVFIuSM4hE2jb5sWidJhwiZrSJKQDM4T8woX4yaNYwP
98Jxpy9UeWVBY1/VTxZW0IP9EwU8mkwTu670UQ+iFXNNtPRDFJd6m0N91bsZLdI+
Dq6q2n+JsMJjUG4GsYkvkdCveoDVCkuWt+mMUlNoIh2CoFbEhH3o/xZmNMJdspUc
ds4he+ewk++hN+NDW4jepeypumSuTbVElWlnOEC7pB3zylDMNrmfEZFqzf+ydShN
Cj1lDwgPwVx5DhhhE/Sxpv7HF/QTz/UVCOka0K3mz6rTumvaZ9Uct68KofSE5dWY
Pd1gLqUkjgb5KAmXGo1sR61WnAq2P8vs1fUDjxc6PTkCSRcE5mv0hN5kRYUK6sgg
uvCAQbCSLn0RVNuWzkFTtot9N0tVanqC4jV6SviF/CMFoiN6+4nLXFla5qwRlAf5
EqLqR2960BUtGT1tMWwYLcll9en0lV8GCzW5zgwAe/B75awvvGp8HINwyocB21j9
kIFkv4znvKT33JoUD+gg8y52B2PW8BWMEPDwP0/9okbvoAm4N2um8n12chGSPW9p
+XshTJyrRynKjNrU8GgC0KnfEshrB0CwsdXPUXS8+3TNCkDbVF7e2KTPurM9jl+e
QHXV7qr9jPn/0T2ZThqGkjR2GNNPaOyOoUy9FeXQPxCkwZWYF0WGrGFPAre78mry
35nRuR1PYJA5b1REh3bUldAYlkO+49n6qdo2B+FepICwav86PcJI904hEn/dU3w4
8wrkIxRPqBwCFC1otJbskJTeIISOrMtz8y0DerYxTzg/PnVExhV5h1epa2M4s0kT
MSNi5Z2drRACumGAZsx9Fjeb7PvGPbbFcouMgZ9WJMyI4ZqyNvg5LzctPlS706fI
VOVIxqDQ1o7nF0a3BX7v640wiFZST8ifpUWfX+2vyMqsIFebIj+s6tz5m04przjz
bdsWLJZm0y0DTxQRljeVHJwc/PQzTzAOrqsX7/kkS7cZzgOc7pgl/z9v22Nrcc4U
zvbkL8rKS/fb4nvBEQ0h27fiRX2mjofH+Jw/F0ZCH0zVYbPUKfLfZ4S4V92qeE94
/iMsw3xDyDGD6O2ER0lAgO0UsTYJ5asn/6Ca3/T48Giihm7gqVrlXvkZuFre7G8Z
3MyH3HT24xFvvxhK1ojE7DdGqHQPx/e9qv+hlO6r2eQ4FBsCd7ngbd9SfAXsNy33
5iDjyxrD5VSxiPskfCEXTd4WnTax0ItjT1rCg9UI2NUcHSrX2hgweFsPNheY8/uW
xAyiNlSyb3sYnyxF+SbmmG73o5mKdvhOYj/xCcT6jGWSYv3sHy8YAotSptSOJI6X
9Hly6ffzfYPPMDC4AEZgNE+DxbCpYp7+B7OhNHjS/4SVD4Z/l7ibUicNcwsQSiMf
lZ+Dx+ZRNhWOQFo/7y2NYZneBWDc1/hoiSnSoIC5sl8EWsZtgFSLy9e7wemwdR/d
0/kCsZCn7trY7ba7UQWYaMRYjoa3TPkTITSdLJsGVx6RZEPO+wPcuLv13adWE/cW
NSdTUxYL6E0ceSiSrANzLVuvTC7knSylHn44XvxdFMkGfY5mFfUfR+TRRWtFLrYi
9Ocex85kkfaUVv9+60eYzR5n3G6UC3ztLGZEmBlVeWt/GukPwMgZH9dJWRm17Oq5
xtY1W/wOuvQPHi3MySlI+J9UNHyG8e5kOJQ+om65s7k=
`pragma protect end_protected
