// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 03:56:37 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qDtj1KsMVfSPkHIxEUiJiouhXf4oVGhoSDZ61RyX4sudWCmfbn6pAigKYicL9df/
FXqgNA5Fc4Ue7IVgmbdyfb2JwCzRQWquwZhWcIT8QQ8v9aHYvezZm0FmlAQRePcz
cpX8UW5Sc0ONEO9jFj+D9p8xpiOMOWrr51R0SK9ty+Q=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15680)
r/fvVdTX1Em+UsuAM+0iuflZKu++a7g/MQdzz/aYlzxY+BEEOT5OS1uAEy5tOh4D
HM9RvGRLeqQl1QP8ecUcXjxWcVL8I9Pwj5DHads0oLO5Sv8NjYlwgE1cvJspSKLE
haA1FbDy+SpbussG8HvZIcEnhfyQaq3VL4er593wnOcLVGackCBu2DbhoQFRnZJt
8AHTbl/lP2wDvFhC2Kci9+krlJXNFx3+NR1mlIBYzYPu1PDPDUQqhrBUoRH4aYkZ
DNbp7BWOMb3b+ULAlSr13TLn/iki9JdtNtAZgfJ7alVHVTcMpOBwMbO15KN0pfN0
DNiBil+z7H6+NEXvpEgUqJI7/NRi4P+h6MNDCB4zomUjmK76+ILD0tsTgqOtVERh
JlCuR9xXNe9kjxOyy4QqWd83cL37PiIHwIyCobjvCVU6cPbEOBct9/M4rgNqwC/i
gBbF+xqG40hyb8l1mAFcJRFzlu4T6DtTRjX7F2dcmpjtpfVsgp7YmG3tE92lLlrl
At7LP1p56V+wqOb/NQSzpQd4N5MvU8mhvTyo2d+n6dOWVtMSG42IUli7dq5O4F+O
n9nV+2CpgbCrxFAu8D0G+puG32ggbYWR7ZO4JTlwId8GtKERxZrK4AvJYnGO2+NI
2yadyDMsdwYnaOdo1sampihlEzfPA7ZyLB4I+hQd8RsnO2uI1ZlkM34LDUyJJJuM
1YD04uUSj6F6kqXxv4vbSxL8EaFy25nuFoUKZvx9t0RMyHMT7823xWEEwvqGda2L
NaGbfezmUkYRUdLgX1jdUHN9i3EI6jD6Yn6/SScSuE9li/6CKD7wlQGGOeENz1jB
wE9ICPxoDuxQXcBlw4NOoZUKYAUj818tVl49y1J8X43Oid2ZcfZmPer2lTVd/ncS
iiEnT11pdf493OVlTMfrcAK/mjL039SAxczecp4kDHiaerv3K38a0641NkLwqcAg
5dxflx4rjBSTYFyHa/p6/MrZe+N0jqmrDfLWy6SSeLRpNf8zEsVotd06jfDbcBh7
4YS65iIz8IViwWv2WTztvJ4h/XJovKyw1ytmVBAeJDQD4vt1WK5aOGCKB5o1UfaN
XLUPCUPGfG3Uw4cAekEbzMM7udJZfNtzjdxkDI/v8x0iwJAQoxZEcHM9zcBbGQmE
Sqagiee49CAEQoK1Bhf2lk75jB8VJ66s2CWIY8H3wi2DnacS2AxQcYVtiHTE/Vyg
X1KOGe3oL/26EMbLltIJlyV6n2WI4NgTjPsmlaaYqJoh2I/+vTDCbp2ItBN2Qnov
bOij0cZAS34KBDTjJH0giGqBcLyt/pBup52UmPIbI+7j0SN2OdbsTMHDL72IE7cG
yZIfvyLVxQYgcV5EAVygb3foeqqaML99J1iXSPIoFyWOEPaOttYIDNqCTFpn8dcp
nSNHYR3wdEGsOwyJCAZ1B78H3WN/+AmU9DZBYIlWjPfwEvN7BqSd2rxHgDnFvRST
gj/3SS6yKM1TCTplrViKkNrtbVRruEvqh+YnKyrucPzQrS6UyIISMhf4gdmOqhyd
G4qZi9+mTe4mrHS2jSE/ZPO9iZGScRDBsWGt0WVfVaTr4hm48VCCntvPqSpXfeQp
AhWpJQ+bVIswfvDoM7dB8n24pLqp8nR3j/ccUdY+6jrVs6cmM0TpGSYTQN9KipIO
Q3PScDrYZ9Mo6yc1W5B6QgVgnifJmpLoXPrdOEnhNkf3vJj00s0CtcAs6/4D8931
2kOnbQGGU6xqwWp2JYktgol8C7d59uQ3OrWkdJI1rWfjrNz+uiQMRQNXm2B2x65N
sCCGwuMv/2nHG7DSHSAFxodpi7bdKuvdLV+qYA3Uz6mKoubvH2qY4jUC+Rja03/I
TRkPoFbJdLQQIIuPxrYlteQ9dG1tz4Y6Ex2MsaV2YvZzmmtSO3J8m5Bo8GY9xITd
16mNquKznSWZB3lsWcw17b+Wjiv3pyCrmrthI7rQB12jgfHjHmnLV/eVSgrbeOdj
oOhW5H1qCCdRH+4+2Ai/s6pHMyTXhGGRGkyhhdZ9B61tIkzcjvd0Bekj1RDMPgWF
SXcLjEgdRohST9cZc/JTcctsHi98gtAeO1zOmn+DQwMbvADZdttWPnaD3DoHQxM+
NGf7S4In8OZO7BJryFe8GBRFNSKqSVUW0EqeUvco4dRivcsDIvYtId2wJL54q4pZ
DIYCpTGzWHzllNcXbTuAc1Ca/RR90icpLgf0qDEM+K2K4prj9IaVAcJ7wvb699tv
s3Tpp94IdsBPe8xh3ZOn+oTgl+6nKzyuhLviIZecsswDB3UGQlKlHP6rwzeGJKT6
oDaYpuclTbGHjH2DNMw7cYIX4ipG8YXiSS9ead9imrUnzORWlkGwnGq0Mz4Rcq0B
x+PJCwGwPlcJPoGPN6GO0YhfMKVBMANM5MDH8pj4vQfY4rEvMlKach8nBZ2x5Kld
D6ClSMBjaPSMBkx0/zCytwzRtPOh00KmUMGrLpeDHxtlG/98603+frL1FuIDMM9J
VcwYNYBjmUSgFTMcDbHjTA2CgMFc2WHLN1AB7EqLQ67+ZTuwdn6LpV341D+DYF8p
wZIPRRmwCQroGQM6o8oLfQMoigmWi1fp/S++cNx2Irh4xLEO3qAePuNEDLmXOsu6
6q8qJjD3lkqPwec2DXz6PoPHoliss10v4/GHhbYS7FATCe+tqcQj2ZJtaX6OMGSb
hAa1aRgexKUVusBZAlAZAwg643PcfNVAaItUYmbxBXwECayPGyjyQz0NDbSERkOm
WrNnbBf9QDKzpJSkIx2TCknaNBSAYlEiJX2oQs5VV1o2huBjzqUfERCO+aqYcLKg
jKWCniDByxKMwQgEbFRDO18ksytVaLKsXZqL95N7uJBK61Uib9EsFoVxCFUkO1pB
/zycG4uX6kPEqrOkAlr7dt/CMsz72yci9f11/uPRiTjKoKCaD+ubeN43EL7gKpN/
Kgm7CP6BAyFZ4ay1JRMLZq5LrrYa5wmqXYYc3OvUG3IFVRHGczgLdElzGceHy8WM
XQI/fsI5MCMPlgdK3QqX4Uyiz4hYOTCEokUbxBEB5Q9nBlmelGyZSkynDyanDP6C
RcdHQNc5R59GytqfO4F+VYVvf4uPe5cN3CRvj5HFSZZGOivPrItjM0sN63saix7x
3suJ+w7dvdrFHAwZv9mydJxd7O5MJLUE8JQf1L3oZVDC6AaBYy/OrKNPfs1muu1y
tjAc8yvUvaMMdQz2PY7bDqSnMCr9LpN7M5A2qkh94G0GPyKDmygECLf04Ta2lkow
jcS0Zo+EwfuIIU/Zchbzv2ZoeguUTh/Pq2rgqqANK9tnTrMSFdyn/KO//7q5efJn
+Ox6JXx3lzOuwDBqVddmfYUahxQh2+VDNnmmvkXTd0E2uXLzWA+Islap0TEJsZRe
IbXLEQfZU6k7FLiAverSez6WhYqmoDf9Cr3YSTOLjBd4fNRk46OLUbGzTr4M4pyI
1S21YzH+k728o83bg0aTKbfl8DQN/1a1wcGkr9dO+CJ4LzbudlJXtSpOXs5a45bB
KRX/+oSJZoCXamhLF47+3UjfgsRJwmLCUo1Nxj5qtEw0UWhEkk47udRrkWxRLy7z
TJaTQWseRLWmSneHYl2QciwWW3Ul5LyGu7LmZr+1Lh16X62/qwJ9IH9LPmayqasK
rxsTUSdvS/uWc/DY3yGto8ccVCsBSpWQMFeJ9RIceU0SeDGxjFgI5AJLww6fx2+I
HNm9ecSoNfgfkeLMgJWazZ2wV0SSGPVCWpf/JrpPS4oCGG5dCirujx/JX14ZywXE
F4IJV0Gzn9IKJw190F1j0zQTZ3NjD53Ql+By9CdfSwtXpYU71SOAkCrUILX/5xwn
kh2N3ubtYftBiqdF/Hw4WjKTlNwl4EIp/++dUMOmnQtNTzEfEHwaoZ1DhblfQm51
D0gPZZyGWaSEzGylzAPcBfrY4EFfLS4nR9RYzvytnBfa7nw51yF0YCnkD8JZc4RI
oZFMYgVA7QGqTLs7YQ0+nx8foT06l3+y4u9rvzjkjkzjKwDbI1ik7MJSbQtawKah
mWfZfTB6G3zJ0wpZLukCdZ0j3orNZK5e6RdYS96rj0UZfI2zb/EhALb1dLZocriP
rq+B4yjZZagIe1YXDZcx8oHwVy92v/9Pk6UiWu3ozLJU16HQ14P48g6js1qykf6w
Uitk9hlTZTfGXGZQVYDwgQRnCikzBvRbWabjH1M+Ole6B1yBYya465C0RtozjDGh
q7pcWIN58mR9O5SSWrylqnS7IA+qB2kRbrSpyrmsnx+cBMdlgDuY0RMznGDLqfYn
sFJ+GKZD4cN3RCwS8+wKZuUpvKg+tJb/yb2lWdVa5N8ODXaKVWTVoPgbJRd3nthu
Nw2sSp4DFgwMugbKjw2NMD2/QU2vcIFZ80JPsDUU+Z5rbvOW+qxKAUobxKbGoirx
eBM+lznBEZCbyxlTbo0gxwFlptiGTX0dmZBR6647nGHvU3rGh8LwxYHbSJmTkHZe
aD1Ifvv9nQam6cxPiQKfU17NWffjJhp44ZI1LPfBwmZKt7vbEvO8IvgyjTz97gdZ
/UlZd91abTnbgPLBXv8GaDotaaqT7MkEMn46NuBrQSicJA7vVpIz1Rjfgqz7Z3G6
hZiy7HPYOhiVJsV/ZYKn021kWhzoDachZGtZArJ7Tf3JTklaUy4WmsfigwE0Agm4
HoVZZhS39+dZjYydYxGBfDPmoVQJIGDloNV2Tm7fNol39ZYehZTO55BLj2mwZlPZ
044FWCW2aIkn+tu5bJ4alj0Nyzbi56puh+l9yD6ny+KPIOAuK5V2pOI4XXhM+sLn
UXAUeHPqvvafNrc1mBz9qniX2Z0iI9r7lP07avdbTSmk9AgR9FvlcPNsgmeOarWK
0U6MGR1Ck3VGA2y7jzma7t3PvQzuMzDohmkZ9EX060zaXfhIeOy7CAto+ZeZ3Jhj
qto5A4WbRVKkwL1rzSI/hK4fxUZMHivwO8JA4uX5xMMKG9gXMBW9u+kKco21Ks7v
i7uzfmAfwGMEnSbs4np1sqGiRhotlYe3YDJ26CL3LIfkOEe2L89dfSoNhMWqMPHd
tdinApNhvckU6TtVCnzlUtCyJZvscaxWS2ExZhGxyVWoSc6PFJzv1o1W6Xk4OAF7
G4o391P1Gnu9vzLuNFcCeU9mUFVbIyLGwo+Rv/zcQHxTb2JbBTQGOIAaN9FbGE/P
KHFKO++jekioBI+hIwbPnB++Pf6LwBqU707kRrhBfzKaybGHNDeBFvsECVJj/qJi
KPyvmEjrZUYr8e39gMwsoNtBiiQiYe5r3qOgJBrKfI65rbsFV9cRpsfrRNXE7wDK
Zw5b2lwUew6BQzmKpOUiOS+ifZsYEST3VvGkojRxGzaIdrVJDTjMSW+tHnGkEGib
CU00ZktklgUfVSiWdqrozsqw4oMOBJkCpjZRABNF9+z5mM29jkN2NpfDc1a/xlyX
gsu6D8IZ+WUqGJiyHtQQgSv9cyzWMzo7VpWIUj7azduWYL9KTekO3JZ4F13k3qPG
7AlClYfEFb+rNgjIUZhIs1AddMJocp6bxSWG4xcv5c2y3JpEY+TRCg9nXZJYGm7R
h6Nie+r/RfuK0SNpJ2BZVQb1ZxCgvcJLPDDCGa8Qc/a8qRx+ooC6uES8yj+LRsvT
AFKnzadfhJbeutGKk8jdw8D8TZ7G/b59Ynj88eewR8Ri/y7ZmPksJtT/y7o+EaVd
TdOXwfuWQyIUbJbNFY7xkLjum00uSopuAb0JjGjmaqpDLVZIy8l8VpfGErA3nC7u
hvlxlmXF9CYTb9V5/zXOilph6Ud9CWL2KNIwb2JLI+WeZgBaYzqyUPTNizDzJEZm
KVEAbNAU89jRbSiGe3aUXGKKNZ0Tb0dYtHoDSBvJc0QjlpqsXwJw3SsnL1z7mVsg
7VAk1Um8ijvdK6rC7q4vJKhi2hc1H4UogyjrEAs822HG4Qn79a+NgELqCmKYOgJp
/EDNrmeh7LdvXreDlFq/5jR6Wso8tVcmNzOJGDQ50qrm5iuhzWPTuDdl1T/6j4EZ
cN7GkUiWFFAk27qpL3g/GifrbdgDBm7MJIpkN7BQ0oMfmdAbugmep4BHJ444eHUG
3dSTvaktY/uD4oSVSAgZZCq3UWViFfLN2+jEvawbmxog8Lofpg5BVhujfKkbU0ej
Xwdi4pE85dKOeZWaSnyhSjwVj4JxEUAIo3T9A+JTvtGRi5ryTGrBHadD45PfAxJu
5uhzhfAacG7T+W122bYAvzQDUzEwYuQ7+Ebguf99Z3ODvvtMLgwiaz6zcEdtgtsW
mwYXC45bZr8D5ZrAHPFjpJfXQWEB43j+KVmpv39q4Vj6ucl/4K+6zUW0eCL+YP+i
wZKqv77ocNS1wvri2tSnKRse7sjuSDLTKDMuzOVCUcTXndUHUUZFYZXEi+M0wUVk
WOo5o5DrkvaQNjJdfY3PVXAgfeQvv1rvXn+rYJZThBFWuRG1CQJLhRzwiR6sRDoX
emk49YwiU3rSP1pLyURaRhd0eWmckOMTfSU3/ZLa+N0QMla4lolguzleyT6lgBcZ
AYjrR0kGYxgk7kk1fGog6cK6osi8qMG56of999SydPGK1hN2/5xnrxJm5j1PmEh+
DlTqCb973xHGwml06Z16559DFH1ExOh23/oiB8G29KC/5L4xhIm1XranFqTflS/p
g9WJH0626NrjCoxeN3Xkh1yJTEtxL+C8Ydsm7kGbbVQ9e2AztWhPJ1mvgJotS66V
1k4Gx1wUGSKScpkAUn+CEFev/G+LXrAeDaL2pKELRBs2dSsOC46nKxq4WIHvYot6
o1oPQ1TzU7q4IlTlACuH/JeIht9Lh+i9LcftNOcOwQ6lckN4u+TbYuCzNsBz1gPH
rDpnW1FX6pyFWZqF2gYR5G1GeGRc/y2M0BzqfTW02UWw6MKzdRT0tVgUHGhGnSh7
QwMtU+nSDPN5FHUXN9U+g0L/lvR3XM0zUZojWKRZMeTj8lAHQuGu0wxv06+S5m/9
wrT49vTxMUaB1nJ5bBH1eoWT/vMkvCCggVq9SCKMj5CNiE06lfYFSac7nXkWRDGT
iVGZumO5mULcljh1n+EyJrYBuI9GOKJvV7oXHBk7jmiv51S4w2A7OfNy/eLKmbLK
ABIJg9z4hyuNmy5tWIojr94Q5ULzp6QR/Ks5omHFZEAhKbSQ5ZYHAfJl/jvSV7R4
sjnHRWIlFXqlgvygUxHNe1ubtUSludYWx5CKYTYzx4VifIBdy0f3uyLdqOYVywFh
0j50A/4DeWrc9JyXz9avJ4zlz93TD6MS22MS8KGuX3KRLTUj0FCSXzLutUaoytf2
Fv1hWLfL/XX7r06oQgMWgpfW7z1nJrrsVTt6c75Ods3Lp7IfsxIM9b60A0Yc6g48
uJJepDIB7wZtc8B/0My3WPAmQy5gOu25lv8OLC1HVe+YSq9prY5WR46hZhntePVm
XbL3QHYRH1dG+dzTy2YqxOKQFu+3HayWoFZWEOBzDCuPgm8SU/DaDMhNTApiIkHu
7fFbsMjRq7FT0BQwLU4dpynv3vqcK/CWP4l213Z27gWv7brLHAUwx8F0a7IgtLbV
gGtv1VPWf0AHdTPGIMrCpOpiWXNcP5GWf9lCVaqUkeefHR4RarVTu44tHx2v7G5H
3yDDSUYxEeXZaob7Y5UCJe7cer7hShRC/qKJ0bcxqhGlp2rx591mguoy//CG8QYm
9abp1YmnzuidolNkwJSaAcLiZewv6L/kN0rltA4trcYXNatkkEi2ToeAphQmgOk4
ib2ADq+c9Lz4Z9lWjkoezW4y3jCQB3axxQhTbPnO4tOPWx2fTuPEOJYHJraP6TJA
dbiA+/N1M2y4BK0wXAPbEZkBh7sAEqFbfV4MDQWYyPqOKyXk6rOcY4LNe8vOh9c/
YTnQadjJdCLnl3/g6/z5roZMnrKevm1jAYdZMMLVjmjwuVXlpwz2T67XsWL/QY31
WimR1lZhJHnQFoo3wn03RicmETIlP5cKlmMa8wC3W6Nklin3IXrmBkvNN/bRvd4v
i8H1OmMXTiA/9Hih1ONl94W9nLK40mZfEs4/7vfj5c5y6l7SiQHF4zwQLWdLEbth
svQrW0tc3uDc0hg5m0UhtbBegIsecHS5TJ89BbH2oFPWy0+Y7IulOv0lmbIjwBD4
I91ac/N8BsUnwh0pSvG+ioHHAegXLpISYqyWJr6x0foUvmW+u10KYF2pLyCTF4O7
kn1YB5nCHMgpFUCMuDqnrPGRsOmRwCy0AmVIisksnLXt4kJudgoqsJN4qCNZqfGw
1pbNM7aBwDKDZu/qab50YvSRLbSZ1Q24kkS23teooq7OcmceeO0B1sB4614SZH9/
pIk6+HHahqIYSLQfD9nquJHRhD6N6x1lUoSpr81RwyIGLQyZIOf3jHgAsT/AAXVr
RwqebyE6tv5iLh2Up/NXDBjvFbTV3saJFuilfhblVcxsT3PQpLdvgYQiBZVIosjK
aI8+3pXG0/+Temge2ckdG4stI1B7SYmd459XBdxo1wi/aDns44mh71B23GW30HsB
6tDOTe94QJY+jgsEzrwVPw2WmyFoehgd1ViWvql+3n+SYjyjO97PctprWWT/aRFQ
cl5RNYsaHYtS/krbwI1QpMJBzHQGxcg6c7UdajSGXKf7Ib2ryHQqAW8MBfhP6cm+
UNbtscZJQy9pFzhMlGYgsU/gBFvKsP3ZOKD39TEvBh9MWJ32xqcpCmuAHwxvgI1o
/S0zGgz5gnPnbtxVtu+5hlqn+o+2+lpsJAcSJvImZV7Y05fiVRkelGX24F/LSgG6
LUtVjJ8IuH3CePAUDa+0bDpd2qBxlS9ALZvdE46Tc6zWPVSm3Oo9M02Zp4wROnsl
CJy/H/fvyR1JCgBLPE3LwVql5lqrwXl0WPQH99KSX/zFsM0Dyc3sB9AFH6/sso2u
M9mYZqAOPh4i+OSdgwcKuGa7tl0HvSIMkoxtTzaRRarFlC0hNuyKkBFgms7rL4kI
p4wctQKgLB992n9hJCWGFY2ymyvZxesq145HGND+5wDvBlD38Y3KP4IfdQPDt6Ed
UtShLtMB4kB8XonWCKcDEsjwWxvMQlJKipvmXJlvnei8Pnsmqz7lIe/90n0EmuKi
QCduxWn8CLWo6NMAOwhf+uJSEytINmQfOTLZdZkuehIZ2bLHroDTpkIv1SGZNweU
hf1DCQ9V0G4ABG7RlcpbDNnK0iVmY6f3s9IcqXuPH/6gsYP43b/8A1LXpdTdBj9i
LRcP5G9HyOHgbrq9+JnjwLK8Lnb3HCd2piuDx2mq9ZviI+wZAk76R/ok19vVBC52
VNTAuZO6t67Kl/wfMdsi9IlVFs+g/6G75pzmBMnKJSeNwfWzqh2afc2yZWfhpGD9
PqWT120OhfsEBbJw3N39Ltk05k4jXrueemhPhWKRA0CwBDWTyMK3nG/ZxdAwUYrp
oS8YPFr8l/8OetjQG8SgNRa34t2MNXpkUdJUCZM/lFZp8ilYa/LSyPio2rTLtwbn
aTf8kySvJyhFEsS7EOVNz5Fe5mClbOSUtE/9rKUK3a4z/yun/pork8Pmji5KbsK6
GuaD1jy4OsXEJlnSYHvYJ0gTI1NRwOjvNpbIMfSHZYvb85IDhwIP0+zuRER4QSin
sabhFbevt7IRD8gkJ+Sy8P58y5cAAB6N3xkNNeuR8u+FWMJzH80uAwyAucJW7/+8
4zrUXaMUmGQf4Qbz4qITXbYFfgVYPfFwU4wkvUXjaCM3nmiVSmbIMTVRA86VT+67
/MUFXhUe0cS2U2bblW7jTCPC3A6Az1X3C29tR8QepyMHuvYkVYrEHww30nlEWFFw
68+CoqEEpJYIxkHL/lmbSzFiNRoF5qoqtG9N9DzbQb0M279w6afQg57H5r7f18Ae
CCnzK1sHAJZu288xm/DYOnjX6qksYPqZ2+yKTZOAkg+yBaNsNWDxVPenCNfFjGYV
RjTB0zcfAGpXdeN4qUT6D5fMqnFpA4Tk3zc7dQDJKITHZUVTWekhufZr/0Vhce1C
jpzZs5fL2mxGrD+MeUeVEcf/Xa3dyPhb6Sk6JHLFtNhb20N6ssJTwtKtLsyQRH4E
3PIqi7LdIQsyqqqXN7rb/hTrTrDZIuUWT1oSgzDGOrrEPycBIEPfHTaHQmHQc8Ki
+yIiHEzvOVSRtF8iYRoHZJKbCNspkkaMhBerKqcftllDRZQiJBC4o+Ka1RHZFmjv
vBWRSuYYohJByvmxcEPH7RYaJzQLpkfIi2d0FBq4kwNdpdEMDMJ6VxwidZ83JnlT
zhwEneuGLLZF8TlnwL2Llgph22UNfIQSjq2dHGXAzD4nrGLZD9vR3/wHs0vl/8dW
dojy9xkOPSeWMaacjX+Q0zPpNFM6JUkmQjQiA5Ab8WwHPpLv2zn+lfbfpuQ7KC5O
7h3Wc5ObEOZRuFkVeKOSS+HY/+eGAYi230KyCofRaBEQ1cQGv5NuGLOP8E5KptA2
ii5JfKDeGMlAa8JZXfhsFM/OWhsEl20EaL6LKLG8lLFd4pbBG8leRpN3DqVqCm8d
cNkIp0Uz0LUoKr2ybW1zWywClo4shVdS014JtC6fgf0BPETuSohiYrV5oz1AF2Z7
dlom9XZg5XiLvV8NDC33z9BzP3MNwrqOtdcemsklxiyqVGf8bWtLGruDpQFidTWZ
MU1TrJAhUbU9YDzKBvnif31bzmPu6pdkkU+OONT4VidjH+RkXUZiSGJSI42YajFF
XLWcmo/uaO6KLgWbwsT9LnxFBmtZOjzYcbwlqKMY8KHW2Uy8M6ewlU32C4XTUoM0
QrSLbvFUhEUMNBW32glkp+YsKWp0eOAgT2GlW1h/KWnZGXlS1YXaB05OEX4bTW/l
g9bQ6WlWBgmP2ivOEPRJed6zX+xDhs2oftVG6UDtBcCApABYY6ZDu1YSlYavj0GB
cEqCjss7O0DxUwYz+7M9euFjlCr65pQBEUbTOkT29vBT52wkqy/v+A99/UUXW8j/
NPmxqCF0bg7OrdrSSn/kr+ZlZSlsdM5TgZvFFeDNoIoQOhLCgLU5M2BzP4xsXmfX
0vpffhs6tH/O5rzxQ2It31PSGZ5dK7YzQdkG8JAvDNwjzS/vKn77K7cW5UNJu5Fm
Kbj7ryj1Wxi98n/WyUbt2JRiaGfivb2gf/e1d4ua3ULsKoJ0zWdZA/dPjiqCCogb
Q/sz5HVMx/cW18Unb/RkTjROX/oKrthXtuVpVbr7KWJLVEB0YaetL6OSkGt+a9ij
MgrldDxr31DVi2+ZceX08CEk/WQfwAyDVCthMip/MFg9PcwjM/BJt2BebibLdD3t
wyL4F79Dym/kUcGEYx46wJnvfSockH4J7bhszdZYjUvCXNSeT8aUVpMjjOsK82gD
Xy/4hk41NJhxisUzvDAU49srIpgxfsYINR6tTEWXms888AWmhBhweAyjqw+7dnjc
GJGh2vkbKJiFNvU4wry3VwXddDXkqtktMNDIUuwvRo1EB6Vo70czNAs+KrxkVl9y
YvSB/ck//B6LuIwo6IcTAj8dh+4CHePYfXRKtnq6CZeiANADHKyhapDt/w7ceZxr
FO2o4P3uJjvLhws6MM1vg0jkuKe4AqsqiAYPb5A52Pfw8GbXmQB/XdZuTUpxr1K6
dLtzp8elUBcR9cYwdEttWjjiQYMJFa+tglBcc5TzdA0VHKbTpYY5tiPR203ZxyFO
LOo/ZT6/IOW5+ZXUPWBphccWI3PYPC3ibfcA9CUqIF5UHQiLRe/FjFOC63npnN80
s4eab1cvMno5HB1ElnUYbQ5ASxoXtt2EGn4hksfcXm5MKRSvOYK01B23BaBXsN1R
4uIvVzluRJncFsMt2s4A9dZjV3YAM/zG/zFXHZtk2x7o58LAFjVwv1iC+zZlXDBA
kVs0iuMS6AcLTKEu+jewimru333BVXP6GytEJmq/LrHdjvMobSOWER9H6AurjYAv
Z5jtIHFb6cv0I7nQz7nDCnPDbdJCg55RY5sPwMdu+DuR9XHUHDBYgjCq4c0gTdHr
TcuEL2NcVnZFtYeJOuGFu3P2kI89oftYf+JDj8JlZvwLGVtcN7+eNRSgzw18fkBV
gfhKDXjuBNQzTXIY61LfMh2lkb785RXnDhCECT4X9VkMVFzDZ85pY+3UXPCrH1vS
3lhewCKDRIYVT2UoWjFi7p2Po4k/OZbLxcFXAfRLEthQzcKk7L+h1kcgX6N2Jj9y
Qj5CjdfrOMSlE4cGirFbI+6/MBdz0xtI8DuDINaKBQtRdi30v/n2LmBUD9QS4OKj
DwbNxXto5TZA+vSg5Yf7w1UJfIK48BsnXKFcZuegOj4/dssQS/5phnkSB4NmwFP+
N4RTpsDJ8nQ6RgVGC4hLFgzYBpDx7ikR1BVeXukbfDtfSvKxRVPDtiPh3T8YGOqi
Jgo9U6mW4CVBg1W8uXGkPkpsrjCsvq3Q3tCAYfJ3J944m5yuDECIoQbNJAZBNEpG
cT7SmsydxovzRk79MU3Q5eVpFjEaSGEqEx3+KsfiB9XEGHUdo0On37+zxZXX2roa
ILMNiT22z9forrj31FKsT/uaIypFdUhjEQndhLwFu5osHRtROzkhzLQ74H8gL2gb
kIaLsG4OUjxZcgmhuSaECoTlJ39/I5av9YZOP4MnwKe9Hk/JoYiBpDrz9RfF7irp
vN9p3d2i8yF6OMNNQAoyFSTz2SipmO773jp/euzhFlS5qWCwLcLVWY1hCAFAiLkK
mz222szx6XER/kYMNpugbfb/6sTIunnaQElbDwqCYdIb56w3FB5eJ3kbgJeN1aoD
Jbd6ThNqK0cWqy6A3WPRlcSojieVSHf8vlU7zoq8jixtopIDEJP+V0Jo4E9vKE49
UbvPVx9/V+o+49eG7YfzjTO/KseubNSMJ8vY7LP3ZjQNinETp15sf/0Hf5TaYFw7
79gnZG8WX55dpEu03v6wNVtq5SxpXYPlTZ3C/dng3AoomFZtZLXz7PkeNMEdEL+N
tJysOf7sS8nszzWYbcDGcVgDr5oNMuttCHVx1SsBnwiUbfhpIbsVYvn+hEVSyokQ
aU3pmRwLi0d77lqigWS4okRd0nkFPqfDQXFymxBsC7xJrTqa/+WV49dtxJGK1zD8
Vay2GhrEgA4iCXyz2t8lOHYzrfWajTx74IsG+FqdFABZCm5+CL1tIexzmLKyHBLC
XIO1Om0jFoJ5Q9UwkPAKo/k6n9Tr+ClWVzzmiULvf6Xm4hVk9vcgOTQhPj7Zo65g
zrtsY6O4EY5pJdMcJb5zRoqtR31byMzlzHX09Bbcoddvvgn+ll8Qpu1rCAdSd4is
jlEqdd+H59OlBQdHH0kPLq7V8D/rGXxkM0CYhZHDAOEUsPSd58Ww4t4/cufCkngs
VuAE17yDuq7pNOmRTVhinc3tnwzVS78cZmwt4GB8ocYLwAaXmh1nLbVp5fs9iNK0
4KC6rTpyjgQcCZ7gieZNJbXKEkCx8yO+/IwDTTBPWz7D5Qw7wbv1XF7wFlzdoQay
Q/sM1SDbeJt2joEQVVqFMGITpqsBaxVfhCtGodgwqjMPhGCc5pVwUvuVx/P8Npzk
drCt7OD8iVCecB7H/Xxq3/JbmkDBT5LVuaz6TWK+m4qCstw24gaz6NoJXES7warT
LbRC1VXWlrtB4CRJ9SDJYKDZ9n/bix3NfkmvVQIrojpzHVK3qSxfqGrWajHIpiqg
SnmkUPwguZhzIH4DfiF7sBw5D949QCbDanR6NURE/GC80UkQ+3rwpm918tSXBZg4
Z9RyOPA11NZucXoWgBEE2iOgyLkvwSQlqGf/sO9hUmuD6UAHvD2IDxiuMWw7t4Zk
s01rxtu/yDuxvL5Lb3Q541nBVaaZQ9fQSszro1NoYgMHqXCmNB05E5yZ36a8tety
g3Wt00J30IKGbrE3eqZCBruIX9h/cRnvCtYshyFuyDBoFNibKeijya7IE4JEuByT
lDPanG3azRo/ydLbpaaphwVayKjB6/JQwwS48Ao6niYA38dc+ypisxwlj7o+mxIS
cuGq1/TAcV5mpoWNIc3STrblVHbOaOPBrYrGgYbLQkCp4+aAJS4plTLgHxjvs/X+
DfPPW70Jvey3oN4xGub9c0JN05GEULoN0AtrktdiN3seVrWRGtYWkRnM/YJovTOi
0X/wELKEcvhglZjc2V9fk913az7h04H7S5ZqB5s84219eNy2+T+QPOSF/lgLE3yZ
69i+K5Ijai0eZLR3RwysJaiCD97DCoETtGkEeYH3zayZsnwYvwcC4XGmxb0HaBXq
RZgIdutTi7Bs75ImCxWP5owuXZQGN3aFEphTya4Ull8vq8OulQ6inBQNCy8pWzkl
vlH5jgTzhD8Cvtm/Mq3DnBL4oytrNXs4jV+xOvh+zoDs7Zljrqa6vmK9/Ug2sD4b
va8GFKmtl+gbsIGeCbxtqLKhp0hG3NvIXJHv2GsMStBIJwToeq3qLNT8WEDSJ3Tl
o/mXYMFtQPll0U9Z2eekv+GESc9q9NkqBwuCcro75e3BNekaeXDlbSd/ZRlq7KBo
hiKc0vaeJiaBshXe2UUsYNzC1Qi5XSEqm2aWjQGJzpXbQUnNWczgt/Qu8PzB0MyT
6fafBvJmsy2fg5Ws9J/n/ugO2egxSm/X6uJCBjCXiUBrY1rYa9HMRH0kzI+0bjtZ
bt4L9N2Tm/bCQgkHxtVQTyaBN98pssY9w1BAPtfPz+LznELYipS+JFdw3kdv+sal
Bs8srzyyUjy9JtM3piQxW5AklXRxwHQxOtaC4Tx4Ttfpj5Qqua6j9XvMgXcuz0c+
Kh3sRFHNxHcVq4syN08tNMOi9avgIGInafwXI2yzTvUlwqKoSPjC0aiuNv9uc5hK
9MZreKrs2oqLjDZpiU1yJ1ltRxDRjdv5wPdFx4kvGfvXPY3zx7rC3vref/x/7F9i
CIzkYlnle4eK2uvjDV3IiXPUaBWlioaAqeJTaLcxwXpRWpqUm4JvXbmWn5aJOlJg
qUskBDUUmIolaQOzQrqVlrYtgdXPrWHFtYcptaVqSqIPWJFR/N3RNp9v4RbkA8hb
f9QZH26UjoxlPe2UaPzXdi3+vA78eYX5CovE0WZ2Ze6f3WIC1Q+LbJg4M96psuhV
ex8fbYNjTK/0940Od3wit+k7gfFhL4uGbyTt0A9MAd8Ibef+NWT92D7wj1KJ4MDY
etCcSYctKyOVIDG8OqRlrhVnh/Uk4sf4NUyHl3ztWjcAaCb7pLv14jhhIgpoGQGE
tzeAGUzDMOgEUZ7aeOHgEH/bSxPbvzw+ILqyYON0KxXzqe9K1O1k4ePktT/6vE3j
Lcxw8M7+8c1HjpdMpOxIsmuA2kC+FgNwaO4IKi2RWZDXid0zkNOvxpGWMISBNuD/
COEdWkyi8hSEM6xRrgoMkOy838ml2FsP5qwLXE9HJi/wwLxMBg+alavSUNPMHx9b
2Ko4wrOqmCSwaexlcWF78iVlMwMcbS4AjoLY6veyPGcc0V4OxbJfYUILy2h5wQP/
zl7GJBY4lLpq9AXhW2gZS9Xqd94TXNRD2Y29WEAvYv/0ue61Km4ekm2YYD+jA/Ip
Sphh113gdXQ3Oo3YEFxP9J8Zn6fSs7GPC/fNGMp7rki1GRnz3AtvbHNnq4TKFn0A
khqb1h32utAK90qiYT/qlhZMi5SZIEAHqYLuzS1XegA8WcBweSpcOTVw8gwtLEg0
IKV0p0BGuIjfnahRpzrZ+LhTmhR7CmWjIKeDGn8uddQc58WOa/VjFQ7KRI5O60jI
vIramcGMnJiDjNqvLeJRNXbpW9AOPhQGjbpp6bGwFeeSSL0zuBjMR0eH/XO9T9mi
o6CDhpGlv6EmTdU43J6UqQ11vDiEYd/5EylsEnwdTkUu2ayoKIXsU4RZjA5l/92w
f1NNpKRenDeJOqVBFVO3pjsFKhXi8yeh8LbftdCQUU8wv8gagESsZ3bQehkq9rcY
MPnaYK+H4vucEm1eABD+7Yvd2t+HzdVDYMLwd86UGik3Gof83/wjkh4tgwFuXGtX
vqdXz2uFCRX2/7sNeWt3VzCTTbH2P9gZla9CFvuQYOEeOBGkdCAgwQcMeTQ0Szew
iKTchM/5pSLpPVzfl3ChEg35FXr5UsGI/rK87stwqO12m1q9VSCu1Mnbz8zYDqhO
NwBqZb5BHmQpptmASN9MUKjm9sqhNxVeM5uu0xreVX91ap4RjVuwgiuszjxbLUv+
kf8NVoEDpjpZVAVDFFq077D8FxGKYoP/Yi678CRFSqiIuH1S8c89lSch0oeYgZSV
XwA3683MZA2z5Rtaxuw1W1dw5KueCtRDkVenve0ypOVuRwIFvbQTTCVnFfmIe8YX
VFj58RZ5cw257ex4vL/aTU+1EqU3s1kltZzfg4oHXSIyhYG4lJUe+CX+qKTYOrcg
i1yv1Sc1lRNjpRqL8181ppVQTjjZVed3aUpvfAEcgkdXnZjJ2mrLy6W8buQVvA6Z
ICk7ShHk3xhlsDHekkvPkAhPr1mHtVvSa4T2y5HOYJao+FscVQHpbq+JCk+vUNhD
MR8trFXtiwJNbCnikAid1Ij+Zd6R0r7BX8FGNYdZ7ptKdXDGiRRfecyz0ipmzTQ7
VBdPawkYPyjQSUVTfWOAhPXDfDT0dQ1OfsxBX+uDF/NuIb0VF3l8I+3s9xIIDbhP
YAmCQWZmzCxIVaBih12b9xxhxgE633a0U5Nbi+FcbHYfufowx0KRD7VXRsrm02DE
2Ru+jim8TY89+B0/wVKXPAs96bimm9XhycpQhlmgNuIKsqM6ATe+/Wtu52/U0hmV
Lfq1/8kZpHyhzFcbgrRmBAeZ2QuduH7OaAtifyyCvTMxLB8ldHjtvRDASGKNBj/H
nWg94uJXO1dfaV1lSLatnSCqoiNOZtSmK56Aux2Hi97ZoP9AdtMANcGvHqfImetp
8bRmUPUC7lPkJH3XcntqA4SWOVRBX/LF17TdCxiRBYSPwVgKR3aMxBW1bXahLlUl
sZuWGQdsF7orMUyaIymX0GzjZ3G7wmor+VWW+nWw0vD8ZsuRcI2OC1pZSKw40iGM
6cD68s7LNBC68zZAcB9O2SBKw6oalhXVDLPNKw1Z+YaHWqCRvC347Ppx2uyBIX5Y
sVMs34+uGqiBaN+LpvM9XlIuyIaZsIsg35zwno18qQs89LHfLlBDCfU142+RcvfX
d4V7yadjhcNDvHYTJdNH2m1QQqgb25Yg/DeffTAi048MZJTnRoIkMXye7jfuaErC
iVsuBwNHTTLsJt/hMEUXiXVLw4Lu9Ms+cryhanIV+0DVQ6I05Gs8VeRWQHVHAKAT
eLEn1/5Dgh44pWqRpsHP8zZwDpKRMMvzhONtKNNsAgTM4xF7DV7swCgmpOXG7zRj
qPUKMR06uDxZVdatu2pw/VM+nL3hPX1zW2pZfiylSHVUdVhGFS3EksS09BEw/yHT
Vk2lUf4Br55ZQygGaQBeBgEHjKcU5VOBme/sthuaETrPzAWdvOosRPhfGDri8tbp
5rWh0rY1q2+oCGhumwZf9kxOusT1hZmqIzqb5elzq7yPfh3xAY/A3Zr/mqMFWwfp
9rZ7QWAmIpIlKlVoUg71NtRmS0f0Llwzp2+k68Vl5Da7/L+8LjZUDSpaWY+YJ/rk
Mne+9S0K617AXh8bEgZ/qluHTbgo5Sw9iUnkAeXVPP83LyC10NirwQ4bXiJiqeqC
e/AZj7C0mmuwmx0IXMOJ5j99au1P9VthW4lxXcfbYQyRD0/Ukrqbnbpc223WPkHw
zU0LRXo6BS9SsMfMfNmR31FKeXNCBn5/g9Hzgyjy1mbG7l6+JXXK7pVN0UEtt/zw
+P8vVPUQ9a/5Bkz0YqwACvUBJhGqfr1VCFDUj17cvt7vKPXfkWNusFItkWC4FffU
ZPh/6f/dyKi8JUylq9MRTlkxRKAxeVqOfFQFXLZpVKfGTAICXVYS7fdNEgA1LjFG
W4MJ4rKJ09b9OxfponhMow9eZgWXwyfKB0k9jTUB0e+m7dN3ib4FUjriGyFWTBDY
CjFo0V/Ns0o37qTt6TkUWtkw1cz/8qVYYTf70apbzSCjnBIRlp+KHJn+Y6dBmtBW
pdvpz9jX8++pKsMBiwQBpBZE1kwUP8VtddJ4uGEhdC3FIJy5Cesd6WHXemM7+ZUo
J3P2Awg2e9psLJVbtmxkaSEvhpEsr9Il0hIgy/x+Rl2VVJvrq+qMCVtzHBw4oDlF
Tu5h0BPdbmo4WXOz4ODAgo2T6f2iCgG1ANBQWSnaIJJeeHwaysU5dIasAQxzirc7
SDhLnt7Dgyqtu2hCYJvQbo/ZgeOy5zk3YYJWJzAfjiigUg3k6IYWwdXUoR07AvTU
ioajKbmC4Nd/uiaoNmWCNHLaYeGegQezt3h6Urli7SjMSzrEtbDPCEBdYIv8hjh8
qJPgEdWET3Gqy3ecOlGACpwLwrQ5P7ArKm9Bs/fAwvAFXjQFLhzCew4wglwdCFxS
WPbNBoJjLDghXRZtEBP09sfi/Suv8DwnoJC+5LXmIuFcbZQdLbdMMZ8rWQI9S5Lm
WxM2DAXbqgFxwgRKxEziBNxe0zyWZrCPFktY/WZgVTMIGuCceyzTNMn92LjHOAiA
76hPjM6E+K3AG1bL59DlsOna0wBTlJ1WmCGnjkW7p7e76bcnSKF4bo/jGe33Cyxp
Si+B4FtBeUUdzAKHO65AxvGWAOmPw6uaJ6ndU4R9umrc+j8yD6I9mnsmsaGcMnDR
By/CvEa9cGkXyySmp2DbgxE/R2FdmQcZpQTVsMNfyRf1vSOSu4FQ9FdLwFntggqI
7xMFsttOsg0JT224N+scoqgYp6+Pewuimxg//b9uVprvz4mgLDExn0hilMr+6Brk
SY2C8LT1QEHRjIxa0Vmi/4jE6C+8kbMz174GswSDmL07fere4oJqZb+nw013oEdu
AwfEnD+6MtYWELMEPcOmE/AGJxfWY5rGDegh2yPP+ryu8IFkq7iQW654cIIUKpAu
IN2bk/TCOQ+FUmtanMQWSSj+/YHUaTc24rtRyMNSHo877IiMJdRVejFuwq79+24J
jBMrasD53msv8V0XXkxrKc6GgSuUJCc8Yd/8KVYlVsyfPoZw4Nw4NaldIOCKGjcS
ujVB374p6AHzKsK8dq3JwcfxCjbfHsqimmPlDset+WpgeLM2SMqmQ2SjQTrCJBGK
JGTQ2yh43kCw3z14m06dFtxCqpO4WNBzIopQHCSGx1cSTh8moZfqDpfGKsCnF8pA
hdGszH6JJJcWwq75ILR7rFv7pFLgw+eLZfcNsfadadmaTar698DfZ8ezP1Tdn3g8
uNzHSx2fLR8Fam0dZCDT5ejqcxiSIH1QO2yKElBrYNALpdllsf/pTS4kacMkZuyA
6kZ81J42VmU79I1YNdMTmhagtF4YRXEXkaLuVPSz+vNkoAi8zfmDdC/CVyz7JJ5q
VfjJbLvaLJBZf1pe/vZvXlJVsoBMPxux4SoOAkTfelonZZ4dj3DGNEMv+eMjrv+d
H5ENRlIcIvhDVkgqY20RkNNaVujVlMKQmK0sd995EqpJnOoaQ8qaHfx08RYQgAMs
SdEeltHTnIyK6gpr6hwzw4lAmOXi9nypl8P9WxH6jeOhe94pxMUsIIxglLCrtCP7
K0l2JUGAB6Cf/SGWAC2vz+DdoVQ+D8WIDvqJcOMIayc+Z5jTfSlrICQVHkMDJVPe
a1rRigWOEHgClccaErNLFnsJtl9zYR1RH6bNaSwO56AiPNqoRLCcVPBI5sP8iw25
bc0LxGLgWH246+VhxZhBFa01lQqT699ibbmz4kCcMWBe0IJcZP+9bU6StMghA7z5
1Na6DNKaz+h2S8Xk8WZ4k3N1gMz8Z/F2blRClEou2i1nC2JSCHSSJmHw6lMlXWsE
4T6i1gcaYIzKM4BXdmX4L4w0NAWT0/YzQcdAwORsvfi4ChFfQzA3KdircsqwT8zr
9TOAM6ydtr9bUr8KD1dO34I05T0+H6x169B2vSFRKJGPu+HU05wqVPM6ToB4Oyca
CxlkE5ri64knlcWG5XhAwxI7lorc3FS+AalGV9oNCsgd1GN0BdverBkRFS/z0BpC
Fycuwev+xEUk9uCMKQ7NI1FunTrW/kw3z1s6cg6y6aYztsgE6MZx14ZiYD3rvx0g
ZciOG1pSRwoHNIutlYG1xhZ85rc5dkqSvpHOniyn7RH49kIuDfSUPQrtSpbQJemJ
g1LjQHpm1eiN4cwewn8bn2tkWDX0GvIhhhing9c70VMMYkDhK3atGj0tr+nrz3cq
iWJ+B8nce7eg6W4kjGyEdPegNb0feNEfLiv84sYjln/UztLPWd775KGOVmB7beYY
aS7b4gsCoa+gbXKTs1/7QlxuJHw+5CJA0BQ+WuC6JSdZ06C5YpzZgcN1UNOyDi4F
eXioG8IJARK4eVRUtWaqdEh6c7UVVSyMjPxPdPygFBpxpVzEK18g5r9h9QQ8cIGP
uyEF+bqyI4w/Qh8MK/9juQtUIZ9TyGfh8+ahu0IlratPhZHSLg/ODak7KrNo/cq/
fPcili9AUhlBdNGsZcsZR/mRu9h56e1c4cCqnEMMqQTS9aGo6zf9MosI1OHp2RZV
Xsm0YWnFhkqMNM76/+HY5HDZH/nqmBRAu9kKz9/wUGqBqVANDvC28oA7tNgOJiCm
eyOqNq/4p+RP8O3ltrM+jHhPtF2mhWhXYXRIe4KEdIZC3bVqXECkwPCpYykCI4d4
RrxSbES/Gl6zX1UqNtUGolbqjDyjOSUZ62SKZtl9qnL+C0DJAY0efzhha5EXwJWe
6Xa8PGvG4JsG66EH2vtVVZHZRnZG8Guy3RSzO6StF44eVMSxph+34j98yTEsBjz0
dB661ZZgSJfmyKV6hZIuFgeTwZHuvD5LANb6D89U7g4HcvZB+0dKAJM13TVaTW9c
1+irHorxK26q6I2QwMFzrFQXcCCYG54ZXUaGB5EiDrSkwDoqhQX4KCUkF94TJPJc
f4FHIK0JPChL0zrw/urThzUEFFGXU54NpfQP870JGcM=
`pragma protect end_protected
