// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 03:56:34 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UvnUCtbtNaLZi486AQFCGhT2m+jp8/YqGmr4oz6uOtKspFo+0v71/CGP4JP6Mrjc
tfeW51QG23wbzjuoztETFA+mtceD3pyaanibNAn+Q7RATMxm1R72b1d06ssPui1t
GVDDcHAyExV8mjaTneyFjuskDzzv82Vub1emolSfE08=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 71088)
bT72qgURDY7LpBwx10CaDzDd0Qu1FsvMuTlHAi66jVy7JocXeGsLIWmUtaAg5MEQ
R+gQqJi5Z3KHxccvNoPUWd/SGmeZyFiAd4AYmC7zePx2GpQM+73fdIyyHgQlCj/K
oHWpLocS4A4T8cUDr5BgZKduEp7kfQB2RT3/9A9x0MfnFi9hQJuc9JJTSsy7PCW5
h8cf1HAnTMO3IpIIbtd5wC5GTapi/tuBzVJayH+7AocTjUj84xxRYxYkyzC6qbIt
hGiJy7JN7PUurt5noSNCDkpXAn18EPCE3U3sQhDDZSy/9NsArNWYp4xGLzGdfHI0
wBhJqB10SMbAAl+xJlA9YlWnGsHPx8wVLsA5o31jHDZBrr1Xzot275XsawalJqPU
uuy9cpf3tpl83U5JUtOF9YTiig8nnboYF9e3jN5Av9W2cZ5/6/+cldfmMnlq/XeH
6/XJpUPCGkm02ykqgVCyC+4LZjusTW/6fJH2zkXAiSyx1yVNxrRq9W8ciMTmWZCW
R1dQ5Mctny2Zopx1R0FuSGWhkYO9vjH0re0dMquTlSOikWB9UcIzjjwZHXbLmWEK
N6PEZUm6D7dGmsR3aoyqGNDtXmZ9qCEczZllbsKLgx6ssPc8leYgB+6tsiWUWI1s
q9zUITuuKZdf6MHQSg7VEVVyriESprjsuzgFOorBwshQmxRLozc/XjCbE+CNprzk
YrYblP5I4byWNaC/gF3gDTNqbv75Hf5p5HIWGFej7LcDVJoz/tVxp65/NsZ01FB6
+y3ijlpTBv84GIbOKVnJldvsmM3oX8yYiYM2qLJCgyfl253adie64b8jk+GontnG
Z2zECDVA9l3xeJf2sfA5oB44oWZxYzkVQ1gtskQ3r5b5jwqQ31JjZD4mugmHSOyR
6PdTA9oOVC6C004gi78ThUxqLc0SBjJ2e212WTc8mS/9OnBR7+ENtlze5/zFw34o
uBf4RjoqCdW6fZuRbo6jJH1nxamd+O0pGZy5joWInWfxB8FSR3ALhjQ7wCGBCPHq
tbiB1gX7owDlTnl9XRAmxGhGjg+c0gE6JL1GWMBqz1919oqAVp5sKu+4/FP0EUx1
aJ9vCMhBAxwXzzPGQ3yRF6xpfMdWOxlZ5iEVs/JNb3EjsOpPTnM5UmrUn2kibtr+
xA9U7kQPQEo7D42p+GvIZ4CRaxXB8DBQ1HlqJGucx86abJrrDUv4rLUT/IK+yzLD
u6GTj28Q9a9xCxyWk6n5bVMlm5by3TRoeLVIoc+/lvB645LYbBotmn2xkci6Nbaz
QC/aGCkJhz3X/HYi3bmSCj5pgUJBeWJhhLflDhyu4Z9zg2zozprZi6/wf0P0BycV
9rAR4/Lg2isHehl5cm67FSSGTR0tMbX1kFvk4hr3XXWbnk8b1PWhYSfX9KVeyBv5
W2xiiWhrrS6bMWv9qENQ29PrmBp6+61WSB/7tbDcwjuN15dY3lCzWryQCz5z095/
cEXInuTGV+x2EH4c6oyTakFq/WQVTcFkoOEAN81Wy9DWTLXJpyN7SrobkSiO77NJ
HdPyG24CUS6b7TGwzKxJY9+BRPSzpisV/7+Wcw+rGQ8d9YcJ3AKFBCUxvc79imfh
Wp4klqwJxJpFyW7HRRxx7U3gdD+SqMQiPtUKo4HWDkQWBEUD+/gCUqmnbktNI+6B
CH14eQoQFc2I9G2x0d4DkJxl3w+6GQItW9jD8dCsATpuVQu8di7GFcmieHL8GOPi
n6xhhhFgADKEcT+RrwbalQUhzxFMsakFQLY9WN3vmdAVrSH0MJ1PlYln2oZBVENC
iamDeQf0H3WYT6SEXGQpYZAmxU3TqvDYwbjY5org63aL3HzFhMPnSp8ZH1oTbInK
u03waOXxEY0bx/wycFYQv3GvuWWNkiqh660cBJdCAu6BllKidm02d9zPxa0lLIpb
0yVEd5jcdJkOmp8SKI6RKSzrjQYXJ1cPkPSrEHAjlNslYHhNPkjTNbhdQkgCpvxz
FrFuHAmce5mlOXEYFH7Mw5kpJJdN0CK7OeYfS+R/giOZZZOq5qg7vXc7DnbqGak7
Hb5RrLy4DNKVB7x9YY6kGGgnMVECF3k9Rxssr8MVCWXvlVeI8RyaaQXJJ4772Abt
sWtl/u8twQJtimPwniAiHwcGqbaQQZdJLu5g6jD7hSqZ/6xr/sUhrK5E1Cy6Roum
GcGC28mH954bAlqGoUyMa3wAu0QawZwoL113u3UMkso0GXg25nHTYHLK8cThI2oc
ROhfdTjnqbG/2MjslDlcA62Ad4iixPMjetnbHME8tjqNQJCeO3OEibjrKfaN1J3t
AL27A6E3Wn/GB32pGE6FIWQeJ3lKn7c0MBKxfY3+b9wBIheFF273PnqqfJrejpms
U0Y98n1KsYDeTA74Zbyiz4nw9YQ2iiacbvIkBN/Ye7hcpl4GUhUJl0ZNZZwN07mq
jEoiZMLMue+S9hMrjZCVva3awPZd3ltI+b9lvbJey31zLyNDtuI6YFqLdIyvJG8o
IBmjQRs9hiyCz7+SJzMjCJ1Dau6sj42I2zBMC0qYM6VCTGoKQZ7oNWqhSysH7DYv
uyGPepdcROoBLkPZSwPE60NQnpWkwel+SVj4PKPTOvJvY6/4rbBTIIcjgT7DXY41
fiOnCnakuD6quG8hh7VgAyLE0eSFWwEMK7Ze4+pBVGOC88NXOJLWrQTHp8+B06HF
KBfMxI4D8kO3X6jCuv1F7INosG8MsnKDQ4eH0aBlTBn15UlyOpjfZNsjSbBS8BdC
vghOg51t88r5v/XJ7aRdWeuR08WAU88jM06dbxfU8GMJhB5ISNnCenA8gl94yYyB
mVH4/H+1mKYapd77VKEZkkCVnbTzKV4coQnIwrNtrcOu3Nb//17h0f+B5LWuNoai
7JT1Cu44mLZCqufJnPU3i3yQk81dEuj4lZnyHsA5qJuhFOgQANdVtTWgLa38BikW
HqUo/97TrAphQgiLXGfJpFOaZEKl/t0A6+5cgr7wwu1eNDPxTH8kExU92fURFeok
jgyn17bQvyeVGoshhMLV0abBoRA4XmeJPE0Bx6L/2SHVJkIgsIdEvglw1FczHgGa
WFPQ+ieTAOrZ/Z0lW6axfF+QcO+xCpykpj8pI2X7a/YOd2o0YOA0Dt15z4sxif+i
2pa6Jfwc+X40F4N3e0WkhGTgT/p9C4vNfixleKmckp+fXNEhaaN0TZPqNcQjbayB
eoPv379AHOOreYcNbzgFMj4AOiQWMUHafLYv7PN/hXvzcF+rQW9FX/WaTDq2z59w
Bbl0BCaSt9+fTe2IBoqi6K2QHHzyEB2lA8+qORo7b8Ci9uVuq898B4ccJxCQhWiK
+GPYTrvWHoGjCGnOCJ4ek7pX54tgAoD8adrVpkDzem5ppa2B06LoQGDPz42yoAYt
cpMYX0zWHIUY+lPXffZ5RI/lxmtzZhlefsVuyZDmnbsrfVWxNZ+3FI6Y9YLBRfFg
oL+aL2T5QQjMnwGR/j7cZeuIaOh7UyzuOaS9LgMEYmDOBZCCdFrkztU+azoOYlIR
PI23rVZQCfxMRT7v2Ed8dG9eYG6h7n/Kb0hRlQ/0wrbsO7ky8e27j0gwoedoHRrF
rytnV41+Sp41zxHMRuiyzwWyfmGjFVn+EqgfMm+ZoZr+/2eHMsuaFu9KmGytBqfM
KNAY+OPaTR3VKMQWVotMV4O/VnV/EmePR0FYdoTTLkTBX+NFYtjAZchtNNJVnkx/
Txb9DaUQZ5SYFFUiV4DZ+n9C3GdKArbOJX2QXgboZTsZPXeisl0BFJoFYkHbk1/9
+LcJLj6l9FQ+exgBopP0k09FU/B5oW1kd7OX8C78Pvv9YnCWCr98g/rp1Hv8kRJx
IqWi3fy/UEowjT6rbWkMNtgzlE/liDuUElmCvorR18O8OplkixS4oF1VdMX5qwYQ
dtWnf2JMytGseJHVvuNSRkqmLcKqyuJifhKR+fo2WvpmvreM4i/RFkDrPZQ1qODs
tWaxkBSm+baa+vxCnN5JN4H2dKT5RwpZt8Extp0N/5Kqg2FHVeYSGhJHxgun8jg2
6AA8PUFFADW/Dc5ppbxhQ28YNJbFxJLbAhKmUlzB0M8DecFYeQOaPEWBq3lsxfDc
eInkM0xuZBOYiWZ0uSAwD8gn7JndYpG7daSpepTBsvykdReDzxu9pqdMcEHyOO+P
0gTEOM8wnuZmGu4pVFmz2X5MV3uC/KLhSXhpz8XRv3ByOtNcJZtsHh2+cLcPbMbA
eTYmEMBoqGXoUrU2d0H7SD5NhraVoFxsBiHuSkcTRwfpdPIuyh/bP7CNoadNHywL
u65cbbvuXMDUjjOgv1y7c7NqlJVnHphRDHdWqLQLtNr89fIJxy9koekEodA5xDvt
P8si6daD6Hzo/m9XuHOMyhWk7dI5ju/PrfSXVFpfLKdjX0SpVmHfPPccf1U48tjw
8SLVYp/FEjqUwlr70eSBSYcWm7t5dSbEvizcU85bUFmo8aULnmSSYHbQgMF06y4R
nDd/EQAlKaMEyWDdzHAVV8SveP3ORqJbvEmQZDR6rO2SsejJumQTOvqKkp6dMVuA
0jefN7IqJQrPmcfiA8CM5i0VAjabpDzsvj9Zy8WTRQE8+7ilY5NoFOuFbDeqGOhL
segiYxD74hp7TCsKaGrjl0KI4RXbvuLkmGJ2CHFmox8X9gGCuj1GMrgY7LJMIAHH
0HaOD86/kWb9ElvLb61T1CERW9EZsD1Q0rArLNyxnRLj2VtyV+UPSCUmkh/T11g1
vm8cPqvBlnfpt8d3D+PZMciXg6Vj4ZMoPJv9lf6+6fiYjvASj7nW7G6T4ZIRJIKz
nsC9RuxGQIC60kpLnRQkEqEiDzrfg1g8cRZv/V9Gp+yaMg2cglTD+MmQ1T1PMPkn
2SZBUAXPLs7jw1ekTgU1A9EqglR4OljgDLkAidXGRTGRwioyDma9YlsjDuMex70Y
9CJDaYuJRU+ASJm1CYCN3x3eKGAsvKz30ZeYBmAHXrXkwdYJ1EsnV6cnoNgiMO4e
E74exnvyfBuMkAC1UeqUi7yDxjQI4hQ6r3d6RW+NwXY9uNXRHBrobUfiWrcpitMx
zP0Rtt1wffM92cWm1b/n6IlRzIxByZ1uIR2P5gXQ5V472KHagmVIPn0+l3Zdo+n/
Yt6tgrw8unLHEsqriE7QMsxgTAsWjq9bbBYOjmMkDPyP60MNMM+7XRv64u/koN8w
GSi9It3ffb289VmAneWzjSwZqPDNA6L58WrjTPSUJI2EC2fg3qvIqVKIPv05qBUM
TgP7NZu/exk2qfaKq28zIFpQ9jF/Zq/i//gzbAcutNCeKojjueKn9D3WH5efet6Q
g2/qFbq6XpUyqaFyrpdQWwgS65y5LDeJsiFZ9ogiLuri/qgVvmhgtTDiuuI8yl3K
PNDHduqX2fk8hG1doq43NbzFgm5qCF5k67PB0Mt0XhYAZkGE8j1T+YDgpVz2Chgy
7fANtjFCq3SAvyPif9FNgFXhg0Rri6HwvFmkzmWoby+Pj0UR23IjvADZ9+HvUtus
fhoqxCI3N40WBf1e3EnAB0JfkKHJb3UCdMnQaIvaCSOp7yxMXszmDEXXvqqFV9Dc
d/HAb5U33/zKPqa6DvDfReTlK+27BA1wN7hk3gQe80bK3kcb4QpowomAC9JiA6N5
3GTnNKH8Qp2QZWgEylOdE+zdExlNe24XZmSDdtJFK1XczA78W7cvFSmo7rMJ5Vcy
O4W2eO/qxBObNn8vu0y8TP6+V+F4THHMBHaAz/s3EI+KpqN0/ScCQFem1OUkG+af
ADh/gfo9RhG5pGN3ODHvDwLI0XhYwW2CvBcQ3DNbrpqoQ0V62PDM2FnZVppCuH52
vGkaWFMJzGrszeJkMWdxVmvuFX4AfBbvx8YFUrmkS7C+9M3FmhkGyN3/gWEKBBhv
L57csV/9EixX45dIHwdKnWn7EuEVl/9t+orjkNznG9DedB6sAGMud5bLz8qB2W4X
4nyR9j+F6ygezz/UQfcX7/jF6TtQC/JmQKa/Mxj80vBFlJTQo7+oQvJM7P45I8uK
AIjdsBunJ4eAYk1y0eBgsjNaXDkEXnW4P/cXH/plTWwPURC2ly9/I+1NPbu4hDTl
V57ElB7Q/uE/MYMyUqY96BHz3uEX7JzGJyzu1bcnspP0b12V/KtleXTSSbYA0zm6
XDeHM+3H7OwKrSKSAeXbuXeBMGXJ/Dq3elS/px04Wk7c5MsRvEHKDl58Blw8Kpsw
y78Fmb6FausoxBNreHrG2Bvap/KVJC9ndwIRDP0KrrCnRisE7Cf+C92agAloAwdk
mhGAm6dvSMpii78Nf6iBg2DivvTcrxNGvNr7FUktPaYJpxP5i5zTdxvHIvIRylb0
za3GGzaOpLQCUxbUy60QJ6VTy/bd3MGPT25TPgyX7+n5txwxOUEK5yvLyawycyfm
w9aBIZepVZ/T6aDPg3dDgsDkCzbxQDrE3vgqtS8WpsdJCk6mWlUPrBBRjdF6DPci
/3uNwlti2Fjlmw9XCGv8kjEyvy3QTzzuhHOsiHWRmBkC2UHkb2E7fBq6vuKkl1Eb
B/F9uEmsr+9HuXpRubheLN+yVKSKDHZhdc9FnJtfQ6zx7vHdmeh4qEgVhVsQaTfk
30sNEQwQPLJAVDvjezjflCn/vuH5ihXxre7AP56OCZEiDnUqBtsMoKsnMM5qaWPh
90dQ1qO56JfgJA6hU64AOFmMPEsJjxwB/In0blkOeo63/yWZzBMzZKkCqeqNb13X
LhWhts4lGF1HXB9LV9zgVRBn/cPI4YjlQFi08g9SH/zr+lioFC6IsDqakDg3y+z0
C1ttYzYoMA8b6Q8AG9tl6uakCP+Pkbq9vl9yBWZNCm4FzHhYGrDdY+o9Big69Fgo
bNqjVDNGMrjBNnLQnIhBk+MOsf1P9s5iCLHJZOsm4daHHz/8kp5vuDfAE1IQbswd
1sBnKoiFCMqxQvwWGTbRCfZSecJ/UpuUhi2MbooNjTraecoRWtfq7dOFbFMGM54Z
msV+SblkRnrH099vg4mxMDoas5mLdcC+l9PjGP3TcIp9V3lxxnuI61jYcgPvj8ck
FPJczurI+2wewyPfgOkyIBWexK+5ODs2ihXrAKkN4nNjcqURkvIZy2IvUo7IRwF2
QUKAv3F5kJhUIhUoIJtza/v9Mh98gitR4hn5FqfIjMY8MhilKgw6qsMWmeMypfJz
KNdDXl/VscdhZvGbfxOeD/+gSD13sbI1xbt8lZxLhIDtt/OIXiFk6FRoKS7UIsAX
M+dS7eLF8jEYp7QL8CeupKNupUWG/65AZjA6KStP63FIOGE+QAzOcOIJRIqOZkKz
JtOJCXveLi04xO4bG3LUkJ+Tyzd6686ViwulcJpyPcNtDmHhacTT1UAE9bUDwh5w
0FjpewN8t9KLGl0IbRfN1oafW8XwPDzsFz9FCfMDafox5DY/Mtd+9vDR6BVyZF4c
FgJekrG51xwzhPP/brpeolmvfwAj4Vyvyl6dBEGCMyAutgqyG/IqLh0eo2n1floB
AAtcbOkN3CMRnqWGuf/aSP8xUw0kWPH42YXGkvUlErLpzgqnYfFTdU2Ib2aqIHnP
sly2zH3mBoaUmeSeUelsm4MovFhB2giayCTMp/tZBP6zQQPh8cdaK/UgTExdRb0B
85lWJFvfqOD4lJHtvnnv6Df9cXioExOaY8Utzed7QVq7nIFElb+UBnz5pIma6TY2
mxKp2waTP9kyBC46/ClOwcxhJhUJZDmuPj6oLK7oqiUBjwPpmvjK+c/F7VW+izyL
832IB1tsxRNY1XLF2vDzSaJ8YQsyeNM/E7mEk/5MOgrxHp5/MabCF/O8ZkrV5o0l
dzQRY5mC8P8XmdC5ni17S8scIrEaGimMdbsYwI0B3U/7QZ3ypJwZ0eilNSQEMeah
cS1Y3P+TnXxxIddwNdz04OYvsW+o7HWxztgrk6WbSgyPyU5o1rtEmkd2D+TDshfH
SmbDnx7uft/CSUCZL3SCzSvXtb7R9tqO/b6RoL9tFPr/zcWdcwcPnhvg0o57UVSC
OxWCjHSFnGuwQg1nv6sK1GStTCeujf34eJLgf5QmYegyQ0mRPQQCTzjQOciRlXy9
GT/UMKlyrJpGuJJRqe8oQZx8lrkS5p3y0p6PY4S8dIL/LH6rwN+PbUj7T+fuXxDp
cR7DMi9EIasl4k1d1lBxIZcHBgbxJfgq5VSYcRiWoZvqtAdCu25zDzBIkVpyOSGr
wtMgsPZ5IuFXounOTkZ+3zqFkF9vjdvysX2B+8LjvnnhBJHtwcK1xkMZ3SogUecL
sLS08+CxXV/aj2uVx3s7tRw/iav1lm9zZqUsUrQklsocUePLkpIHZSV8gwNDFRez
S5gwBqjxBarCIXcwUQCa/89LAtpdmEHuQRCrI21daGABZ8A+GN6Qu32kFDPceZFS
z1aSznIaGq/OpG+9qOo9TVO7IdBDMCtgIjghLmBKpOJIgnQuu/fhTvaqeEeJvoID
9qFWjLC8InRQ9xmuqUvS3BYcki0ZblbyaAxLlkqbvajQUNNsj17oyngWz1DurL4l
FJn0GTnX2gMb/mYe350tiwF6NQ021EVJ4SgQizm4nERnV7N4Q+cx3px3Z54nVgLN
YARAQdoOJsGHkR2GW0Jnhqeg0gzTE1fIvi0fu0aanjQXTzpplAkb+2c/d1TBcMAW
1CQKHVKbivm1uQuIkVh8cg9R9WADohUtPUpT1ATM6zq9sI+Al5J2dF8fkkLD11MG
npfkmeHDTzJxSQlW9bj/vNuAFDNOI0Ls/4z2oftGyKWyTyS/ixfPZnoXV306x6V1
jRz9A+X9zgYccU16kQNmHhKu2iFnGxvy3uXzBVR3NdWmbubLfScyBtwGxnWgYkZ/
2eOq8D8SfZc+UXRyXUDaqif96r6Dx5mu/7JKGblA0RrSH4HRVAFZHPbS66ZC1+D9
BdtNWWm8Q6iiInBh7iZ+gt4qimZaaYV/p/hcoBFiOHk/3G2+I7ZJKb2W25uSzBd4
RdRcDiXI8X3U7U4hetmkFAINEDT1+sK07ZOLW/+I0BIcFrzY0wc9cqXqaaVfIKAY
5cUd4SIG0UFA/mumzXmULLejZnh7yoYOgCtD97Fg0PbOxkVimznTog6UQbXnPYr2
BbNFAXjq+XyxinP1+giZZZVGyFkmCMt8fIrv6NJBAfTgZBpDhU4cDfrgsjJU4myH
TA5T214zbSS0/4f7COnPc+AZtRUuqLqqGfG3+AOl9qCUqmgPEeWlZQB8f/Hke+6u
NiIdHt7tMpoQxBSxdwv+nRG+udPonLv2o4rCMNc9DOtEhwMVdGFjT9UQlM1aqiD9
SjhAItcGifeY/vFdn/kxMMzmF6mU2I8mH51BhKAKLvqxt0inOJM9w/7I4Iax3II8
2bPHzxz20C7z2WwH6vt6yNKd0y3wZtNVJy/xbs+BWZjZ6YInkpeMCvAwu5MNuGLn
HfD0WspB+asOQvE+6ZT5a9JgukmBeJ2YgvIFcoSYQgIzsvybXZBAhFC6hNAa86zV
ntbKsBIKZ6e/Zl6SjhKkO72Vhe6QgjZuxmhXKeJp2/g24G98ngx9JS+t0vNbdGEn
djCitZyPglmQGDgD+nlimv8aAtoSOincoj2FRoNfvh3bMNPfdZ4cJhmbbxhOfBoq
AZXMKLsDHCX6Iuy2u4gJSAo7PCjFpUq9AhjK4q+sfmQ1qgXzWk3Sje1wBnKYig73
Nq92kR/ixNyhgMnvhSmuVGomJ0uDGrPfSlaOosSNGsF1cZU8+a2OUlTIqkwu2T1U
SxXOqXDIjt+DsaLLapTLk9TfzwgvUFc72orgV61TclRUIv0NlPQLMnehH9nOK/wT
FOJMuXKB0Qi7BryCxHOlPVlFB0C3ByokM1O/JcK8CU+pUQV9FEwvViX6KoaPrh2a
NoADkPF+6xVn85ERwUrEWgBPCOLNElpCZGiwmfyC/SegkebCCQ+7eFPDclq4Aiu6
xBrlKnXEIeeOlic7iZoH6bwCwI/cgUyPmXHv7nH/mOFLlRmja+k7K7tCWd4LBGZt
LFRNYSG/6gYzKXG2HnQ7zzlJf9nlj/XUMO8fJODZePYk0vx6Rpqe0LF0pbW0PMCA
CNTVBW32tJUPJaqXH3kgsjta8IStVQ3ygp/xfCNT3g7ZEzubORLArLdiskqCXbUL
ZuH0w+h8jtjGVg4CKm0FV3ms7Mhtrlh/eJiC+ckC+UFkJIDLhQYeZKdgr0HAMpFM
d8XqVA9a9KQm7OEAMrFCv4pgCoUezd5Za0aI7DKMSfO9G08MtVru6QZiALX2L8Lv
6+bqQf0POIhygJ1zSYrKAdSbMV2KNG8Cwmt3lp7RyJW8NKfaPC3A5Y65foqg1deQ
BsbJsTwGVXlUdLALOAyGNe/eRS7cAaErN0+9EPC1tpy6f4SPn2RdXT/2+MSwAFt8
cvX46btpuUdYQy2NxtQ1mcSy0+sZMRozrri9GxZVVSR3eMSYBRjQmaTmL4EGliC7
/jpEeLjIX8Suwn0lwfWoRzKvAIR1dRmq9PvQ2TPUPsMRDXO6Q3BT5gtTb2uZG/r0
g6lX98r8pAswlKniBeT0WITfPeYqjtAFf6OqyzE8V5v4w9JIcyIZRTSjiiAOtNIX
l7Zc2DRBzxRMrvXFvh/WUAfrYyiHm9cDejm0aWO0xo+9Erk1d3hKbJ++Oj4c/9f6
bYP3U/VHZb5HbLC1qIgb6qj7RPvBhLVdcCYoZes1khCYj3EilmUg67gfNwBVmkaQ
n4dLJpRgfye+G5x3PiZEZtntYVaiovSugYlFa5mf0pWCbTum83M8Gdxh1PG2Xbwa
vkv/wrlDg2cGkkZt0MT0mBvMLEL9bu1uCQwgkIhnUoBXbQUGthao2eqcL2K6DZCu
nL5yewC9jAWxshPWtex11zqfy/4xM6ec86m8PIkBg/zurghrQYGMWYAe3nHLPmwK
kjyussDCKhaurpSuKjczLNzH1Uc5ujVdAzo7WRSeImgDA/Z0LwWLmdFOVyHUcQqi
WDntMm40wopNQuntYNtu0XnBQU+vqsf6Ixs+1N/UPJ/Ta7hZriuFOMMTHONExCsB
ahIzVBeOK7+gL/BTN3vE07RwCsQLC22ckQgOVUn1AAg/5UY9adKTDtyQHnfmnfLz
Wr2qoCufQU4ugX0wIfFswMXgAz2tVLKhv5bWcu/4wZo6ezUEFbi0sSG1GvSfdj6z
lH07dX7rdt8y+g0sXzQWKisFVMFNpKfdzZ6So7BXTF+DKJk/Tvgda3GE8oPHDm9n
shEwSBQKXBAd7Ervq8WFKbJUknJ+7iST6QxB5xh+WyB6ZGuLDqV91pgC5/fks/GN
quqEi2FxCBNZ9vT4cXoOockxkfO6gJkI14MVbBk1vsteWERLFfXtD/Xn+IJPtL4O
khPRhm2RiivAui9GuxPPjCZURmDre5js3iQlc9V6+Dp6g4nA7f0zzM2sq8Nuxmuc
kGUr2ixjhsorqJQKZSdqPDKiuTm1QPfnOW3v5cxUzotGQTUK+cFwdM8slHx5t405
ggEtcnnd97OroTTjbRcKGkBu2boRPp3MwR7yoBlE3b6WLXlPB++3GlY0TjFeWfN9
SFdrejHEmrFNFcA9wRyGvvZ1QNNx0IDpFRxh5/DQmcbdjGAd61Tz3MCd0FwBL16F
zEb7WPthqA9UGTQR03Jha19ZkModJvtcmFbQZDmzm0ZFZ7ola2J78VRWzvR+tZIP
0sIQNyMCAel4rVjU0R9guV+dNnKLGU8l6ql3MpmMU86SGUO9+MM1iEzebkqA4tqG
/NL8/pVRA+TR0jye/wTidNtFlbZp0lO5yhxt4mU9aN+A30PONoIuWIaVrrz9V8Qt
EyyqWr+2UGE8yRu8EThunSNKlSEjRRKEdb3n/O6zEl7iSBYNfpsvp9WjxVJXUli3
97zDRxvgMtY4bInMf5e7nGYsbWoUDmH1abZak6QTNzehSuibWc6o9x4M1pEqIUzs
HvjuCgYPTRNAft1luWSldxPIc9LNs1udkCnRZg1wZtNW1STX5W272MqYzS801/3U
83s1dGm84RuEaMOjfUlzcQYaq04Rr+lIpFqpbWiXfNjlH0zsez5lwiJkSpDCvNvM
wHHJL1psGZ9MDUzTK/HPP+mO/tcJ1+t17EaPve57m8XAAaMVzc+OxiCdmZybWiXZ
EWnNB9nrA7aveZeQVnyRqdDba/ex2160BrpDd0jZShV0EK+38mdE105rUnpBNCcF
EoFjiawJWOlUbbuIchM4DH3d/XbGjQarzF3CZFHnMEEzxBMmbOJIsvWjUx/oVbNq
ZE9UrAwnkt2i3XaJ+ZweZKxtX+le0gNIGMWxTygFFn5PSeJ6u6j0czG7VQ2yX45W
fJG1ISd0pyChjEA+008hXpTbeh+l3g0mpsPDElIk+4ByUzDqhL4zHs1NlS3FCvsw
dl0p+xWsWpupPSm/M9iJAk5AYDr9iiI0/ZOFyTm/explIbRHqkjYt+0fSelXozB6
YfW73azSRMAzZS/7QhpVVYG48H6GcOqvfZVG7c8rKoXRjo2Xwg61VDbnCcRg9f7c
XttIdxpI6nTC273tWZTlGKQ9a95JBJkq09vH1f9egPvrkn5/ctBeEeM8BlFoFaNY
LipBzzTcJKSV0PXdgArw88vNIPXa1ANpDzQny265sjgda2uH26WjbI0TC7tAp/Rk
TEjbCUytQgiAZT9Blr6kbSmLuEGFX0lkzughgnpDG64KxEZuQ+vqv6IaBUHyz/Kp
5uR7nNHw6ve1w3u4ED+uRTbPt246boR387aO+MAllO/ndJCzeVp+32+Pp/qN60BM
eeFAV7b2nsCmqPqv7PuJ1Tc8tlvcTrGnmcaCmbPqDCBB19CWhtXRWu6ck+Pabzs3
JIT2HaWQRYhMbBvwhdKrKBkSqvIWybuag659wDn42gXYmibTsmmQlCbHE/4CNVJA
IrDgKydzDKQOvJqkPRDU/tVABpqZ5wUNlTUZhyPB2+t0l0nA55EHkLTcOACXSjS1
wqSYZFuHmcIS6qO7qAQsHVj2HZRZfjfYN/DiCUrAFVBk/yy1k6JbxcRjVaUD8NJU
DCHkps4DIV8pg5yOXs/BObBPpcfsprOCvLW4Rotxrq7TKAw+3Ky/7kdJH3CpbIU6
rrxycrQXDDYI0wAgY7CZ5byLMCnullZ4jU78dwbbsFy9mz0UBhdZJ4SA1PmilcFD
OQPgZOjXja6ODFUiIcABAp7z5xevGhXAy2vByxPYS78OdeATZTRsh7rBmeNukkpf
XNJMmKcnlIho+yWl/KWsuxyHbrcCgmFGfXvTABzVwrPmazY1kcVQyQgVmUB8Q6OZ
TRRx1bQ/YZr70fD6dEkCQqInQPmXQiq8BMechNEoMMc4JCqRkbj008uCAWng7Ie+
K8JHayFfZEEpY/XQMMG2zKaZHOsDTDqdR7jHypuIcLBYm9KcffiDEt52tWnvpSvs
Xwloz2CE/0fS/5RzgUoflhCA/Xpq8r4Y4QANoE3dOTU9Tr+PAn9cmPjKJnxufwFO
P+6w7Oe4/8VQubwgvWlBo1i2XAtm7W7givEXFjIokcC83XcuWKYKWVHLv9YujMpv
Q6Iyd7OTFpnhazX0VF9GGKumdBJYqlI/uUD31YNl9fA79GsMuRj4eQnWK+yYuKig
4QUxbpnpvlPVPeDxyF/McWU7rjuH9005TaxUH/8YeXBKpHDuKmfTic+VkReUSk2f
hg7Wharn7saqRf0TcHziQ0ae2JpnHRhGfOTUuD8JaFiZNiFUAnZhXcb598P110mA
9YRIq79NaDN/VUBOikZcni1oEqMc2ktL1WwLv5tej1c6ADMI8DZZiuHWsKaGg5aa
y9Nsew8Zey4+ez2LgtZSSNmRmxeqtzdvdhKwTCNd90kNIYv5J8TlWEj05PKXyMuX
1hmdA4LN4YRzIsBAchRO0GXzhfa0kEJZ3MwVWaii5fa23WDvvM8NQmpfM3KW6WNn
A3pkuSJ+NF7TI7ydsQUHTQR35hrqk19NhWNXWLzbzd+sfEA8PI6YQOwprCA3ffH7
WyIG7v5nVJSlCH5FytMi6zgItKQGFG5AfWhPAEQtXPP9ZNjCyUteR9CgT/M/Oens
kxIDF0dEagqcj9N7IdwkfXCoqCUMLHR9Pd9lKghSjzjCjDhT/l082HZ5Fa8VlulG
MmMxYtOFvC4FYAdvqV1Y/Dr5pVQQhhWD3GyrqJpqjwpk8bKcMzKhrhMSUkEdBLMG
YkhjpHWu7QYYzCCQQr6gnIZZhJCyFtfhpe6L7OR8ZwqfPQPTxhMode2M0hdIjG6b
ZZNIUR9gUyHxMMNZ+1pEtn7SKlMdPeiKcnZvtev1fRKqKiRcFuq9GycgfqPE/uym
BNUHp+UmX9VgC5Nl7zadTx34R5r4E4Wfqi0XImlMUE+5VdJ9GjlZ45LDc/IK3zYi
GczigU0E1UGgmRFsKUwTY0+5EYBOITU0/T4vw87ljiYlU1UkzssSA6vbwjkOtYC1
+W35rCb8u0mkfZgvL3Ce+WiShxPh/bl1BbLKkHoPQFkofbuiPc/9Qb1Tp6FujfSB
faXuVDCln8zNUhiHJmOP6wAbw5z5FU0P3jyxUn6Y81nVpZz9p8hmfDOjieTbOP/2
ake6Y/B/4/Rh23WwmMgtJdgX701qQ6LVVtWR9Xau81QRRk6I9Jw0Vj6WSJaqiXU0
gYUZrgUkeVH+oyk4R/vRTT3lbtG8wBDHmwVaaybrCqvNXUPPKcoI88bUGxTStkrd
SmRQFto+JrJSuujlRTYzEtxULMfPQaqwGNGWT2weN4JldneBau3Uk2cFC96M86Oa
ZBVh0pqgEZKR67WMyHkOrgO+0shD19QTf0XCjZ1ytdzz6qLs2VT9Qyd81XJOvv6v
ovP7hvolQ7GZUgEYWPYBPAt2N+dMssZoV388zKCTiTex9Zhd2CKh09z7ADlg0ced
/oa+h2aaAGTQXcyRoE6VOI1JOvdgi/VEILkSIMBaAZMd6y3Xve/ExSCkEGMLvaye
brJPrXqXCW1QfgSEHjLH/JC3M7TsRcTf9qPv+vu8b3afS9D+HGbbgvYgdfTrh85x
1e1tF87LydLk8F1bjRLUY1FXNVyuXxNdH/Nwi7P2xwBzPkEb2qzSQC8tP27O7pvL
pZLxMiuTPT9DA5d0oY/EXpMwU8ZbOhXQIQxIm0BemkkAm8ooc8Jw4x2Dle0m2lMk
YhYNvcB87Xy000Fma57zPCvzEwG04ty25gIEENV1UTxlo/mQUeth2/IBBNHcJcdg
X7t1TPFhV+HCRWTnUvd+XXm7Md4f7IbOOHqmuznuKEn6A6QbH/7Uzup6ZETMmnOu
yH3dmxaDbU0EbDvjL5iMDtUoKumvaSs36/rnD2elxN63eSkILeNrctNxIEvfirpW
VBLH05RbyjpvpBc6GyhitSAlPsbiprlhn+iqdeMJqriQBT9XcWVsxPzEM/Mwghhq
/7r/QON/E9rNuS8MVI0TRY7RvHhJXBd3ZhLfpwgPBBpZ1YiyctwNDuaj3GKxjJoi
kYEZo/I6Bdlce8pAOjEygv6/S7aZZhCLK3e5/5svWGHSVhSy/6MIGu2e9TIq5j1r
Cg0ab/YQCzpMMcTmHgfjyV5/1yVhFdmcbspHTD9T9Jp8xcxTY7x/aUGMH4lvBFCp
CftlmIgXbqZ0FDOhTrgx4mcFEdUoUSlsAE4ruA2ii/s0nhOk2wlbPsHh0hiemKOv
YNReKvoVQwc7eCObR8+lktxw69WM5t8PKV5vPAXlHrDgVRu8hMKBYstnwMzs6Q9M
IhATjPPIryNQmbZUWTAjoOcjgHMR86IaDumjThuh3TGYauqIK4Xg6OJ5LO7LlnkV
zKCQIydk0UOXAEUZIwOu7srJAueNBDQ4LQggdF5o7xPNZ4tIqzeU6Ylvd/+7KE3Z
VTqryDEBNbXVFVAmnGSUiUXzykKsH9rPsTc2XNfvk3zXJ3nKeftjTzNbW4pxuwfE
ij9JIAxVYFOt+QYBEA7XWdsVrSCLWQ33UnmhXh6Y68IRxARehWcQxZ2JeNFNWgaW
hX6wfMEn0nqwAUOQYxBJxIezYZHdJHw4fQ69jLuRWhGa9Dr8tV1AhH1aoq+YwrSL
k1g0kIRtFje6tdqMjWTEtQbYYs9DQsarewjhW5NLWETqJvkXOFAmJ64+7zy4soIK
7pnpUZ+AC0P04jES9ZM0VWiozjbHLXkQRPM5DobN6DQVxtyOFLlwzwQpaaUkZ4F1
Xt6c15yc+cD7oNMxcmoy4mqa0mb280VTX/p2tQT5+/3YQUa4mq3TkurQ0k/XMZcO
DZ675B0oiOhNcYI5WlmnNd5ci+UQqfZj2G64ytDmGvpTdobCMEiikuVPnNIpdNQS
1qrCCdf7Or7nY3MmzBVWFd1tPgYs9EirvIAYSfEF1o8JDl3f5p39UqSsUels13WC
WEvC01gk8sMpFTVJq+lWJwTuhQ2rCzPkTDAMPjubKI3qP/zxdy2HHS6ocTF2Kwsw
r6ylebUbPzpxQTmQIOCgBxALkf1VdgFipsqB/EoaPusmFR8o1jy6eqoKzd4Tpw3U
djsUzg25q0Ud9JBrPnnFWqPTyGCqYyHcWX1YKdIk+iYGCDDdQD3dpNpuKAYTvxjp
IpiQOY9QFqPvON4hr/ZG1739c6gphnGB7DxlcqTy5dhxXDhXKnoSBK0u4hsK7aRT
oO+kWM1107I0kepXhVHdGqw62u3G4qN3NO2nY+AzPmcoowDCqcjkAr5rTzLfUPvw
jNAW20Q3WRxtxPxB4L/vLQZql/gbHJauWjAUp+W2nlOW5TwF53nBhCDJMJzInGB0
V2saqExlOfMXyp4R4dsilmEsnJ0gX7Sf/oCMh36VDZoc7Wbl+ldOXje5EiwjWQWH
/RqsLSaslXtDFwWVuOEWJGSAnmzh3q/vWWbPUwsYkGTaKy6P+EySkVeVKr7ex8fU
5EtBwklWFtHq8SeSTiue7xM9ciuqvXJqrp0M+8t2IKevYnx2VqDYoN8rHCwP22Vc
Bbf+T2FWeeYjXclDyVEgZKGpEzKgl0IDhtmBMD1ffJ2PWOZgSCQHJN6cRRm8BoUU
s93b/sQwnM5/cJSaFCxQSStFoXko0m1TlzPAV0LMbbTMpyvh8rSi3ykhGvMgWsaK
Agd1e6vXIu1MmSLAD0gJ1Gud3HGQJcVw9IyNEELdbzlWjidT/EeESiA6X2CnyoFL
HDIZaqt/6cXiQQdEoPg+161TT4l5c8VTbrMkshN3dpmXjSqFwCX9VpuO5sXd8fVA
ua3AHsd1UNvbU3DfwDRT35W+wWGcK9X8KE3fuh4la8zQK2DuKMjFL/rG9Iiz0+jp
vJPxj5tEphB5cOzgUoTORF6qoQ0HVvjnvnbhh4E6MMiKUCNM5t/r8RSYQo7oGRIq
ohv2y6VKUK47kHOMshBVqDMQMIDqixakchxcGvJx6JLvtIIYKPLTuULA1rauvPfD
QcH+tHp5OPrK/mVsAcjsJ21NLFbVDVCe9KN/Ths2CGyE+IN/ocVf2kaTGMiTXYEh
kLzhAlKdMzRC8PUt8g9AQQ/xW1XN4RKO8+37ZZj/LIcq6puD+eOb/MBBg/TJutBk
rT+1ew0//IcPwcusHCUAwBbZSwWDhad+HHOAlg2GHzVZHzWxrNtRvdUcpp8Nf3ou
jZB5cvVnuqP4MHunTj9euUWwqI+7SfEpLa2MtS/Ool6ypyEsKFMMFAT56/sZ7EJC
obDfk4ADtQOwCLv20CmO6vQcdmz+GISc/z4kEFtKWzxYZ27P5X6kByzy/xog2lN6
gmB+Acd+OQ1khm10zRbOlqyr0acv5wcZGv5rnnj3bivymYgdNACVjH3lpTO4MJwc
OC/nkg10g/KZosJqZyy8yJTWRC8BZWnWXAxALOsjCmYWLRkFRDNBtr1hnX3KA92c
0Thf4V+uzdf60rDS27kPDxWTjfEYAIwkANq48oCCU25JiF5r63SOWb8k4FGim+/Y
mYbs7ec5jKJla9v9LFnqmk5Zmd6t5qx+98mHr/SIAxRWowa0hBGDeFATrNNWDEja
RK9eNqpV6Nm6cka9HmWF3KpHZjL73ejniEFcHkCwNo/CKuB3IykXhdZZRV/ZxIAa
1oQfVemeydTj5ES+SMd3XGpd3O+Y/u6QPv79GH3ohzhWIb9xYp3NLgZfljTZUvzl
/VPCoGDfFtSuOjrhSGU3hUqKNo8MykcH7lB/Dypk+laF1LaiADlngJ2hZvG+bfDA
z0ZTwQGRpV9RRiX3sIiJzyVnyorGlvSz0GSooXBucB06Iy+vvpB5bm1Gcn4mlM5D
Jux2xkMzTXMZRLvWDQGNtYe3G9WpZWo2NvP90OeTTTlIJy/cjhMPpt+I80vBOIzS
+vV1AmQiZ7d0vf5O3SYk41ErcoMrjgiFL/LZv0YHetBnAydys0zebo1p7l4K2Do4
Q98/p3LlDVtWm/h9rnmEzKcB8/Tpe5SaksGNTggZb/t6Kbrhur+V8d1kEEuED3Tr
Xzaw+uR+nk94aTOmQ9NSYZ1QCwQixe9B8f42/kx41kDCWNJ9bcjMu/ZAbGyOkLrn
SlfNkmFjbEAxRQUGkVW9RDoRe2Y8eXf4wf+W4BPl1WeS8Lk1Zq22bELtjdtaxRZ1
KLNM+vW6rwVvuePnweoyv5MqzteuJPHjEYfxk87Pw1pKi7l03upRfriG6rFYGAqj
BpXGwwSTIdH/1oBfklD03GDTru1lE9uUxMF+RMid5t+bBgctBc3nmEn7endaWITz
yUhZ+WOlRR+DBtPPoUb0GhqLDlr4hjYKXnatKwDAAZ2Op7326DHxV/dzhsoPYDyS
G/sNpvW0HH5rXeDIMwxeEolqORa8ySAX8ZKrcPBuFgXUZrcHL3Yz5hEn9dO00Oqc
S13L40HlBKiDR7pJIVQ/kdsLiWGbq8yMuZfSfaIMSn8IjwzpezgBXSP5Kyoubaaa
lfPN7+6zeQUt5jz185eOG/dfnwIfwMmiAyl9YYP0KnrWHCgpAqO1qzQX10OGuZpN
j0S327N8w13sVmV6LyGhA/HByi0KlBmJEhzhDdQo36jpLwkByH1d7kDugSvHFoIQ
EEY2mZ+FIuDMNuixK1PISAjpQLvbGQiJZQOCcbxtOc5ds10hHeVEpNQFLlMKFMNE
cTGEbEH/PxxtdpM19h5aFxAi26krXkFKZLbtZvnmDooIBwsJrXWwT1oDcpBedj7Q
l2uIPp+gDyr3cg3rGsDgAkBX1S/DWTnSbaC2PBC3+CoD/h3d2qgK0IjZRQx4oCT1
LYU4qQEymSTaIayGIGx7TftwbbK1xv13KUhQf1NcVk0zrZ6tnR52cYS8sYOKCNv5
L8/HKEclnGxfxvUEf8UmwQXNtghn6yb0G2P565cho4Fj4u3hGXFn4Q4/dIQ0PVw8
s6CO4/OXRMKUTVA5vrnsUwm3OkbKh8OHdniipF6KagUXzeFUGZL+gOhq/pGSU6pE
YTxwQ844L5ld9tqorm25DrOQim7HNgT2OHlub44POMRDDCazwW75HAgv7OIPqWlZ
jB4xZBksR/yd6rBcRlid0IC5t2BYbf6dscpWUJn9vf7ndR9CR1CN+rs/5YfW2hS9
7skFKe36chYNnvx1EYK6vqEr3i0JZQL/7yPZX+DIzPRgFOYkQ7xfGkz86kI07ufN
HnEiO6Mq4/F2CsKk9KaksraYN7vDELbRScAr/GV4/YoZ4uORTtxkcQdj1iNbEHLz
eW7he4mD+WtIL1aJO4wtD4lOPxSlAAekXTHzyzNzXOOiZRuSF8hnjNRJV0yi9Fzw
Xn82ya27A2Gkkk10QeVj6jWOPCd9M/54W/99I/X/dHiDrprOlHrdLQfGVql/74bn
qhjY2TjGnQJ8JpjQWGAzq9LyoFCMYLO10VWM/pvjlKNqQ0X2H9PpPjWkhSWV6Wgs
onf1pWSXGg6GqtGWm1NQm41p6+OosKOZXS+TsuIazbY/g0yna+5v2j7tvh/hbgGg
xY830RbKQys/Gp1cW3ZVt6plud7DQV3NXrO/xKq36jYzDFDwgJpsx8k/+IR+O/X+
HPNH6m6BpK8LZZwfeaOeG7hb3RhkdzMAs9Kq+K4XVenBayoOHQEF0kCtOqkyv7hL
Yf2Qr4m41vVh2w3sltMwGtKatw+yDwSPQWHjQEAyli5L95eD4v+V+avknidf7eKc
NTaafvw1Gq/fIPrg0sYa5eXx1JczrC2BtBY35etjb4yaGbBuSXZLA5WfWhoxrsRE
XXVuMzRYSy8J3sJMp+wOJjqCZv7B1kWsbHECU44Bcx/yUVNdYVs6M/e6qBWUKWZR
/oCUALEG29kN6W8yFjZFTbGtAJSYhgTkmevhi79/yxhp8Txzp5IaYYzXvndSxnHM
ZfRBaPqh+1eRBbMzjQqzjA1xCDHx9YbCphjYS470pRKrVxx+hruBRBIUQWjwS0Ey
RWdpqGpRBAs3MhguaiNPgayAhEo75hAj1eD4zCQSrN2Cb+zgawBv8v1E32KDiLPl
nm9jNTWsva6HacPKxhfGu5HsdJbELR4XSARXnxmfJJbmMVsBAyXsrxctSWAiia7L
ESCqClhT2NF8+FQBU1avlV5cCJ4SA0UrKcBm9f0RtIOLQm6uD20CrJ7y3CoQP/3x
ffG27I+GelnyoHJFnApu2ZYDke8qJzyiyf89a/7CwnspasqKan8tM2fqtpKhLZ8P
jcLWZIE1WfnuLRvPZDe7TdRzoS0fjPw+PEd/BFy6ySshtRWD5YgwhR9d8nNn6X/N
FcRX3ovcI3ybjQVjQbxUaUzcDfWRH+5H5NmkGNcUh9qUw8DzdE2nWwexQ7KwluiZ
vtm8sFQMhWf/TIIiThqqGhNx6L9ArUFZ5ppsojdTA3VsWelQECEfN1gxUmElgmah
CQggQMr0+XSzTpC0D/n4uny6Hub4Wsnm5doB/Pr2DsiLptASkXAmwdLBak3Zx0ye
GK6/fXGc8nXFItb1ezWBJoQN13Z1SItE9SFn5FqGKiiyE9tL0dYnu6VRJSwW9nyn
e2KMig25P3r9tYsHIjmQn25NAG1TKZZRHQww2U4wsMzmYjWYP7/6h8xm29dWJYcC
qgmohVvC+gg7K190j++lh/Vdcdy3xcZ0wBq1OUuXaZiYMMVFYgU7Nit8qqDnrBI8
tawIqwhWyZio92OHtcxhzL8wgCIl/FcErHTC8RYWt/dDNnGcZZ98w2gfDhdklcNN
M8ofAOqalwKJai4fd32NVpdYjj/8am8V26AGcS+gW90uNfM/kHL9VyJuiCMh0opq
wDbIe9dSr030PcNsRdK4qq6jYA0+qd1pR1gdR7aFdtcVDbyjnmty9i/JfYDY2+1Y
VuYt+UVIV4s0vG1wBfKwmShMZNBdwD2ydAQ11JpIQwjM3nZPMEAoGuiwov+usZuN
Rn94XPorEO+SoBoeWl6yASYY0uBBGuYK8oDq0qnICNL7kiMctwrLeuuRph0m5h4o
TE0HkW9XW7/hMhQXuKAiQqsQMzcKlr0K+cf3eOIoU5vfxWeEQNm80iZGFMiq9aPu
kdLOznSEvfN+1X3hvxoU6y+2HvMTWXHKwcRvygzpZ0kbnXeKm8kUArQ4FkIqoX4K
vJdgXV8MwO2VBkUnbgpKj61uKBlZPEvxsuoBWA/h0Rz0ybiiA9+tlWPTyf8Ka08D
7ImEn8Qc1vTskb16oR9N7gNAAIMYQKF8FErJ0ShZqm1ESjNexHG1RMIhTBeGK4AG
w7f9nQlSdkLCgI1eB7igX2zKEq7FaJ6ZkpIW/HUztNRQcqwFV4osRGEIXUYMHcH8
DYYvFkuQUKifthmWEkJYCVhfN1Qp7UgtuPLb4JWzYVAIwDrmHAAYkUo7szdZRKfg
FPjlDVsXCUBC+5Ukx8EhRLpJfE88/2oTQ/8nZsk/9QnqsKK10BmlQdJaOJ4yiKXu
wXnbBwAl2wNe5diFBZwFZot/ApV5625AwSb7GvP2qG1X15dXxk/FTOQOhZXAYPJO
iGhMQ+NTPfII5w3fgeG45m8y77wdvmx5aPkWLTsmJNwkh1nJbSCXVCrFBKQuwFwc
KAUum3+NqS7/V9z6L4vCWSVuaZRrEO0df1C6vCb7AZ3vi9svrHlQxLlMt1e3JFOi
rJMUXTAT+AWkCdaE1CH2YnS8wWTrYagYYXU70VEnMSJ/Is/+UpXOuUsZx9E5QLUi
u68r7kE7qEwC1wMeh9D86yQnt5CpaNhnDwRI8a8vt29wwN+FOrXHvy9+s/nSwGTf
rAY10+c1A6mNzHf+6+Bh3URz5KYHMJ5S7cexs1vIWf4lLmvzQlD1Kg8fGDKwSumq
XVmcprM/mgJwXjiMIKT84SwkZL35Hjop6FVUtdzPQotiG9CAm9KEC4ZiKev0cPoD
oBXVsbYLLPaau714J67mRJwVEe9P4/HFWHM1FMtbJg5F81X3YgytpMJDnaxHjQ19
WFFLIL+UvPqXZCYOIdUVyHeGsW/FGvAgqdJqps72TWzyHWxgvyxnAnYjikJbp1ze
QZwtlit2wmqQjYPJTb1GwkmbPvrAqFgQW0NJMGQ+3B9/M0s5Pw4ZA6t4X2ZEVKnd
rPogvca6/DNKfYpiJzohaqEm5XBqph+QFuJVJah0ixBEVZZ2TCojc5Y5AEGFxMaf
lzemVImYVwDpCrrR0oGg8pbEy4oZzokJGIDxeX1Mdgyd3+n1M7J+Icqjx2+B4Xag
cQAe8u1k48cQoZexvFVnEXkMx1SGFgHxHldaF8xbi1/9V+sCpHPjymkRClmtLMgu
1TL8JceK6W9oPFOi8kgadkZtBSekLPgMSKOPcwLsakE99LWXwT5oPm7ssz/HM569
Pj3kvxQsDjJA/EQ0VDCIrq2yn3oRy+xhg1PjcbVOhjyZsL9tl2IT20UH1tZh2uFs
XwICDdu1PqSoNb8B/zttaL/IRI7IFC6SJCHUKTvAoOPg+/Ekcs6Pr60jYOm0i3iz
OlLJWiaVi562pYJ/OXUFpCBNCfDWo+p1GmPDoEv1Lw9YAoA2mj3tldz/IGpMn0Zq
avfOBfsgJQN+S39YEWDuzvmGdZoUl3mb40KcxWPFADWAJLdZJfpt+qpWvBtpZIHO
2aLINTkLxOUUfn1Dg6Zj5Hqt7erpZKaI2iX5Q0qFaikOaOQ8X67r9f0WR33QzcQf
zTGozBCB+kI4KaanLR70s7WDpYkd9xsYusT+D9lm7yjEpA7dljC6Ei2vw9NVCyXL
XjfF2Qtn9Zcnk1r3QFhaCXT9MQLKNr8yHJhUJL6hKBw5HeaDbUd7F9ffwqDwk4DQ
FCj5nrdI7sRIDVGMFvfUSOTKxnJx8zekhGB+PdNXNr7V4qYmr68dguHwm9sBsuol
ovl8btLAoWnIkht4PrguNdZyjr9xB6sI1muhuqzEXWKkQdUoGoTeWpMhymsPo58O
whyJ+HTG84aLf3UtfIXFaI2cH2a3to44ex9SimiV9qhxziQAYZQBEYMPJvm/KueN
o9FTSeV2qxULr0191GYAag3UHEyPdlelheOwW/GHUT8NO6US9M/bSTD0fb47o9hv
BAZbJo6lYpdJq485DVY1GSLdxg28o9vVo/1rRFwj3Au6bmNvgZmiQaizGur/36xa
LwlsvrYAz1woVhDoidykfovO7QVaO5zszglFkD6bXRBVu97CNMUQ1AtFPFB2eI6e
DDx16iQzZCiG/r8FpqiZp1xSnhXocBUY7xPeTSG1PAAmDCmCixqF162jMKcqFakE
A7t66v6ZE95lSayFICrQggESeeyXkHaciEFPEyRQBeZ1znX8RXkDXJoQ2MySfdHP
+Dq9ID8gEeAFvK2eqrJT14fTlktBuMPVixXZIcAFkgYKgN/4+dxBT3Uz/YqiXpJL
7DpVNZ14jaWQmeNpW2hjEtOS5eZQzUUjSiscwpprtO5UKgSj35R9YVL7AuGDMICy
PvKre0t0xEnPFM6kKyhtwleIsyKX79R5bV/4CK/F9/ThHYj5MBvpcq3QYn6o99PO
YbcCQl8g5Asd6XtkbEoFKFGhu5KPMFNuttX2uq956DW9sZv2IQkiNf7cLHBoIi+b
8A4Qea7MU+hG96vHNHctJJ0V0G9P1m1AU9m0JK29A+9ACG6z8wt62Gj3ddb5mp3x
u+wauaFmAXvwOxrAnrGW0YkC5vtZpnIUIW9hbqBG3b9IIS/Ba4+lS3T8cZJpFPpN
QBYJPbzUcSDojrF7h3M1VmYHYH3NjmNsTjMl9nDyXLJvJcs4T94f2oR7Y2r/myNb
d1SVXbTgUCr7Wi64AcAiQXC12doXMQjeoVRIGsvd4+2OWX6xHWty3d2QK+IAwPAg
WnFpJ1EogxwiGrX8+bAF9KIjsg+cDJNK3noRjL2rTMVBnOKwlDeT9YjkYlVLOSAJ
tPXLROkc7yReQHjNnh+6IF+dYSgGXkSzy+LqJOFjqJ+R+5wt+uhtSMYm9gFDdSbA
KqD+rhWLiPDWuwSdxvOKoTCY1pVOaM+41tGoFV+HFW/WZRLhXDF6P0A4xmByIQe3
jNgkSymjkV629g1y6ZovikJUl3vG77ov++ftQuze/3ypyFSHL+mnnGh5J6NkDzdw
4nQanSMoCuqrljwCHyZU0q9K5U5HMIOgE4el8y6jVeRrgozy2Kb2fuN/LRTyGTZw
cI4Dv/2kBDfg/MrT+x6/dy3mQ5AqD177+46th9zlc4xAPpo9w8XM0GFNy20SokTl
hAqsVWxCFFfMuqlkVHYZaPR1kXkwe/RzLXn7wXUrhKpqq9fzaLL5WvYEdEVF3L0m
hFcDdGf8vnH1NHM+6vrFsXpPzhp3OxiOpQGONGYfqD/CCyRvoK3NCK70e6+AbDvA
Fg4ITBYyor6ZqH/GZ44IPm3BT3IvMJ0Na4Kix7qL1u85jw9LHHllq4/zJoYxQzu1
I4NrAYGstwrfxqUMq/ngl9DvNM32VTeC9BnCLXSfybZ4gmMY4DPJ2FmhhT4c2N5Y
gaXZNZQck/ZRrCH3G0EpHQ4g4OHNkZ93R+i3zfJFyb81F7u0cr9bRoaSe9ETcpgB
nDGOpqNv5Ve79NtMw2GIYrW0+oTMeNtk/iAhjnkrDCdqUruyF+b6cWLnzHfsECL5
hDwvN/UHDeAVg2AISaiUo4iEHGTUD73/K6WCYEf7QDjirwX598F8F9kcU+wuAOZb
FaqpLFpHCBh7qKWQwkNnVqMBLT9dC7PQX47qo7kTl5zKzeY0VEXXKf28ZAUUJfFS
jl2EfyDZv9YKr4M63XJowKZ0KVP9JtNr3+UK27689rFvbjJxYn0GaoVk4l3KM/+t
GQT4UMNNu15Df8KyIKc5zwsBeHpjzg1McfOeoN4g2JVhNDLV/Pd3Z+mZhb0ZK4HN
VnEbdZtdWKJMTLJw2shTS8h82zPifdTHQL1coLFh1pnlEaUxhWFncBC55k/lM/Ov
DEouCGR8rJyJaYhgaRo6wAAAHqaVoG9Wl0C+Je2psICGieN8v/tbynfnBSsoo4mZ
AYXPF8h0bKfZ4ZviLDhRu1JJgHi9jKOuXyXep/X6g2x6OCXV0KO4YH+C9wPV7k4p
Q5s5JL9080lXUfB987fEi/Sodg+X1WgVPFlQz6DuUjMXXaunk1TAWTxmXBbYz6MI
T3KaQa0VFtnIeWBymzCla2W0EI4LkuJ9hjd7nlwPiAuv8XDV8miptXTDHdn7CU8p
kHxaa8Wzcoa6CYH22W6ugjRkvJVQfGnrI5cXGxQBr63qdkDuiZlie53Rwnh4na4V
UBSkoXJNIU9FiG0XNGcKOsI3PjwOWarIr2GMt3zwQK1inSm8i83bEE1DSrV5JN3U
190dDb/3va2Ik4pq5RqVkEzK0o8Ge4EzdGT9QdKBKSFf8fK5cRqQJJzBvolr+dCL
Frp4cx7wEVXUoVxE2njNopmBCSeCy/GTSK7UWVjeDmz8zYrnTe8N4hv1N7s2IsWw
XefjIupy6+cfWpzZmY9SqpP5uUMBWyYbaHTYwjC2Y/yCIQxSRF6owQQ751q+cHKU
3/Isg9I4supzuoGCSUTMtAim3Z7Mc5UgHeUtVGQGbnMirAANdcj/SHp74lDzfW34
lCuMUKNGlibXUTC345b/LCse0aw+VzvfCNag8hN+8+RpcJp4NfbEb8Lzss6cZODm
jJwm08OqB7j05HqF7Dj5rRwTr/TQGifPwCEeuey/FyFMxL1gTXmSw1FgTNh1eqsV
iFNVDogVLVuNA6NlJ1RqCo/UsyJf6yxtDqE98TVQa6KB3Ii9V+iZfpYikbCw8vl0
y2aNAnwLBzX9Qgaf/8JdhzwiTdx9LCqgQgsKWNKagcWA1nNspIauh+StMHcX53kS
S79lW2v870uX07gfYVIaMN/kS8wJ247iiaEFrRufAdkKmDgoNrF8SGvNWRLg6uWW
RinQhYfddhI6WU17cRBXStEulvG6VaU+gRpjHTTj8LUHk4jMQXJUSzDb5vbNOhjE
Q5X3qwgvmdnGD4qk9A/2pXbJHdy6hUpqk0BJw2dsYEUd913ZO99GZHkP3MUpHGQ2
6e+K/UtDsaS5YoKL/b5S+T+NDngfzfujMR54sVdQxcV+5+OUl8cmVAeAbmu6jhfr
9zfPtrxYvrlk1eTC/N/RakmcIArqTirUlvMOI9xb+ZhSYyQ4y0BHqJgsYmEeMhH1
0Yw73oMUrKHKoBXotef+MUt4fMD7dtPWT3VIkk//CzQ410yoTIt/M5vXYj/PCHqp
Hz2jvqoKdbpxEpANNz78Qvqlc0QO0CcB1mUUoiuXtnUZCWfqPj8tHxLZ1vzDyODT
YQ9I61/xPcbChEbiCLkAtU5qd//Nm5GtfOFHkXVa6GwDpW5u5GSn/SBpt4VOWDu4
+4eM4WfBRgtimzLUnc/5JTdxC2iPMoG4G6RTMQniARj5rG0T9HI4iKprK0D8XZgL
RosYDfkE+Ke56rHtExuF6gq6+hIStFgX7gze24bHInXdQYLSeVcGgtrpdrjrxZaE
M4jMHftynmigXmL8ljPMRxvl8QzWSATJK80uaDZ/CJJw+DhNG8Qce2zerlhNeHtG
0sbT4fciOWBERhub8fvNgVuDCXgpvX7gIg2PlwgaKdDxo3omBt5EeehOxI+33VKZ
3WtT3vxNqSeTx22MeVArZbgUD2+LZ7Tkn1FCTn8NVQx9ka1YceMl5QD6jAlnBjXV
2SGYLjNJzoeneKGUke/usJgLMLhhAKaISszs5N2paHspNiBCThRE7o0I7un5wzFx
wxyWy9yT1rovH/BrcaX2QyvtEkXxBEX6wTUNiSmnDZewpNVXBRCyBKkJK/TwTz6r
TRqW0WifEmNUBnnvMviNjPNe3jfs6CF+DToXWCflL+Ryf8fxNIpDK8HantRvpmeW
wtH+bw9FqRQJ9Mg7Sv8VdPNEhQSURjBHBjM7ocZKEniSUgL40+VumJwahwCTidcs
eypEAyUudTV3QE+P8pO1yOVYsvd52fB0V+R0ETowSySRf8EsTfKDbLAOg5mypdyo
EtEDNaeHULr3ZMer0KjSacqcZpmNnGq8fwBh7wi5kaP5If9yO3LzN49/veBohPrg
tl3rRJYgZnGMZcSvHTbESzRXPzO2rkVODqzgBS8KEfzTC647DSqELtC6j8tpoXQS
G0tKZEElo2zirs9Qzw/8H21egGXn3rpYf/5d2CFH191tChN1F64ZjNIteyvKm4vQ
RNfouYnoF0dQETRyy7ngspgBfF9E9FuqUlg++Qr3rbU6b8aN1t33j8X2ekSMuzfC
ffTcf6qlma679Z4mXIQ0AnpB8ChGOAsRw02l7B/SK9ubU7PpqcMfRfCLhGRK2upc
173UIzNWn0fKLN+1xMUV17afMCmGFyuLXL67nd6d2naibGFoN52RfdOflQzdyolm
1hnXQYRLEEc6FsH8p7LLSx6vTr17nkF5WxA4bi2NfEWdAnO0t2wRT35GJzZkhmLJ
a3UK7UpBCCZs/yTB27A3Qo4INRkM/61p9X5seDok663ZDNWrXq/OkYXAMe1bLBKe
DGE7w2RSRptuev8PXPXv/232+7m5h6axskSy7pg7P3K68QuyGNABrlLFkrB6ppaI
tfch9D8i6SDej6+9m8ZZFo5yVzgL500nX8cF+XB7aIBS6gIP0K310ROQFa1iVh9f
p5OHsAU+VkA6Pa3mF4USp9gJJjvsyf5H21sYI1G8flaTaEhPqP8wYLTyBWJ2OYsx
eW3w6rBYiBtVxpLeES5w7ctCrtiPeYh4poIFVH1lVcxbDlU2mb+Y6VzyQ3Q2vVUM
ieNakWB0Lqw5Q2gs2s5ACHcDPcrS9arTZcX4JU0IsSEC8fQ3UlS33x9YLoUQMqsw
vurAdI2R5Od/51w7AreA2fAJEZdHHkzFSq/cBK+LOhDv7Yr63fAfledyFHSylllH
k61O9wsDZmgGxUFFqrPQAhUKYH4JJ3ahWQ8geze7NFoAsw1hWV4FF5KRDyEGAFvv
9d78avofxi6O817NjPbAizChKykdhl6yMAlIq5kfcLen+bNKWqlWsrVgwzqEsENt
ZV/QWmwXLv95GKJqjWkD+Py/ILnSHgb/I/FJS448p/1W+/ash67nVVaALSc01UHC
DWCxzFy/akvIRbUTtWILzsLRuTYU0OvG+IrxEUlU1qQd09IWAf0c3ahPjZeTsZ/y
pOh5JQAYTbVed4gDJDsb+LGOkqAWQwYzl8i/MEp0x3O/hoRm3+0Li1RdcSOPWj2x
i8IQ5zyFGqIgCdy+8MrhlbpvbVhyYvIFw7/+FdEDx5qT3p2V+qR461ps27klfZC5
Hkv4ksbJaV29Yyj/OR/26ttmvz1v8JNreI2eTwFaD8961re15/miPKJaZmH6mt9e
xPJc+BGg6wIVnDnabNfB6dUsONIRrb4KMfv6OnpPl5N4K5oapCKlBDfc9F/DebEm
kvm2rnxN0rm/2ZHgWWHLAsPs286qe3PjiHtcWMKkXb4mOFqRvRTvZxaa+0uHOFAy
crq+avRPEmIuGcI4AoqmKxsgIWY8jrWE17r4340nuRjYubrN5fl3+rKKKyDas3nv
9WLFPTj/IC71pioZoAjCXBbQJxIGaZ4/Nt7c3xns2fZsF/3O96WS41+LBmCR+ZEH
5DhOFD35YxyxyxOyYQHd8NjVwMwyRydzeQtzwhmKeMyoPSkM0H35MEAkpZVykgVJ
8Rn+fVtRoSDiJf+026MoMOulWd9lGT6LJlchXpC7BjldZJtpnh3mxrZLJ6BzLxGm
8xwFze6BeVAF9DEwxLwsBmAboPrkfZgiM65cO6ZsQsMsW5GYikjudegBxVYWM6fn
MORiP2GhnSiiB9LgBx0D+c2/t8/d1qRXAvPm3+czzGJgMB0JSajqs6Ocq2k7BvZ7
jLoqPJCiLDSor4sMQokaQ+cgDT6ItoiGtO+2tu2wirXhf6eXeOXIWpKtYQdPhVhD
aW6ZXBJgpYSh4v3/8nB6MTRSIL4k8UqpHP9zh4J/KOShh1mWytiTNOp6lhRLxgv+
W165d5STfOA6GgbxL2ZlsudZMAiHulTW2n0cZ4t+6r2fUL3ippawvN7LkQIkp6S4
nd6kSXG3V8BqdU2EqSz4+395EROAwlOZwQh3lAR/b6ZiaJpTdbumMwJZnLvtpccz
iR/VjEivtuZfTx4CjS91tro1tBoMOULIJPpYpj7xCHV6GGqdwCvtgHGr8XZGAiXD
Vh8dHa9dyXw3bWEQ453fj+mwX15Ta5IImDREr2cTmn1pv57xM7T9w47RRul6fmHg
JgHOAn076YeVAQoMr0uaACsl329NdF2s8PWB3dmMQpWev7Q3k9dHZcoXmBU5bZUZ
vOvhJH8Lzskico2PH8z00trhBMZaOZHxaaGhdp8pGiDfwe75IJNfkX3Tkyr0qc47
xaCKw3cAmL0xeE0Edc6rZG46vDtm+HWMOalWQe+zkno10Ym+i6B22oon8NuQaBwU
VENnjAsNriox/LnufozG35paoESfPKWFhv33wvTAPbDmwu06vJNlihylRqadaGXo
t6nveLrBGw5qQGOkMNit3+KKgi6UL5Y49cgh3QLdJJbMg7Pv9qEaR/G9horIvMOi
cc+OhzA5rZRe9VanonkUALCkTSsmUuHQKRqXzkpI+cHXZ91od6lEhGBSMDqghIig
7Y6LajufB0QFyMo/Makdb0n9YKGqBuRzbWOB4HPwsp7pIyywbOoB/Bvj44S/Fanu
bGl7v+Zsm/z4a4Dq65zaymgfq++NMZszKurt7l/aCi4Vb9Rn6wiANaahOFyY2PK9
IAwyBKtB8FL0LZ78/ECOblZWEKGcoDzLLInw4j8UsynuVUf+SXDQTxxb9oaNZwMa
cuYbMmzmAwqnZzyME6aaR0xfpSizrg/6HDqTtvSV5vHd1dOvJ4fKKzURZuobIvnd
yi8XtpiC7sR0WgOUloVOe7REu+Bz0M47LYj1hQe6Ynfs731yYW+7U4YJkDghN5QD
l2x9bjSPyc+EAlDvgVkP9S7Ltx4NmMszM2kH4qSacvDDXAI4MZE2NJ/JftrjiEmP
EuNGoS8FC9mbs9roVAhi3c8AP6CNVNhA5wdnrhPnDUkwUcbsjtUGS3bQI81K+/5e
1GeS9lIJTwRAzjlC0dAeZ9TGgQqIoqWA434j6p8NGj0lp5OA1/LgHCe0N/lyOcsj
v2Jin6PEbGoj/SYaCpom1yL4kWZ9ViOkf3JNEC8El3ETlfhxe69Qhw0+ucw132u6
1h9VRCVVlxVKPDUnNmdBbp5gJmIn4D/1oNbgqnKNCpXgNulvrfm9/rOo6NWvswtM
AOcOr3lxdsfxDtriIx7+GCPz8tUsQZU2RUX3N47NIaP4e56j5vlLHskY2UMwXbEM
Zn4/ZGzFvfx3PN/DTHjcqUUXIzE56daZwjF2ITESJ4Nr11Gr+zLj0xSq339spyrm
u9aP/uQAye/X6U+eRikmYXK3/1AdPjQCj34l1lcisFZ0V/8Pn00jEaFydWnVqRIS
oJZbcTyxvFkihV/P9nRWxu2mJcXia86ZLIxnaev9i4bu3B5XFKAf5Bs0yrSw8ryt
hCUDFS8H95CKajDJlNNQ0Bwz3w5cvMWg5OfsS8iDDa0+fyM+mnousWHhxmvez+O3
PCRe3EEyC/jMuvfnaWIGBegJrzIsmsQHdtfA3pgBcHefeEqqdxNcvuzkf6fOEy+P
V4VaYfZB732pHylcY2Igola+gFs/SrebfRGv3bgptawiDQqbXXY8N193PJd98qDe
ShMq+xJVpDd27ohzKzV+lnvLO7meXC9Ss/NyCDEIHz1fD4Dbqh10CehN0m+lJjUM
dJoExSqhYxJHmWxeeXz8SSyskVeny4H2EgXCzhANMf0IIUX3Lf7JcYSW7MB8Ax4R
ktMTDQDzAEvrJ2UwxLc7L7dCSgaXN3W0+lC6zbKyScA8tpt1uVYYsT+M1GZ6p8U/
ZyBGi+Y7vvv0J+ySBK/oITdPlvOPz5kLp7rQr39Hjqc/ofn0Kfn6Dw9hIbE+K0As
wkKk04wiHOlH6Jzbj7ZZVv1DQ+vMytx/oQgJKUJh2NoMf9Si9I+yTODF4hh+9sZ4
lKpHuKMfTz3DBv/H77REj1xzHdotK81dxoJiFcEnc+6Wvj4TR+h42JugExE7wyxm
9k7lGz5xinmZR202O+xmTurKYXGYQuedtHXctDMZpLx/7gbdYySL00BpQyCNvlHW
NlUpc8HsE6fbo6yR4Kx5ulRlDOKWTG0bFPhza972Q4LcBcnYNqFKrSpXEjiLYTM3
WavHNpYk5wuAzdEgq9ItPE/9C/zBUhu528Cw824HeyDgJLF7ZDZLPtlchq73JyDV
rPnU30361YVCFOGNduVzrv41xKnfNCG+E020gEZHYBG+RnuFzJTH9veyCj2PmleJ
zIwBSAKmkohid3cEVHvatRTSF0lXFzHc2+bTZmNPYwDABWCh3eoiDO8nOboWFskh
11baXOcSj0tO9zsDfgzEcnBfnZDhUyS7/YtKLZMkGP9LHu/eF8EnTCQxhXDs+b/n
T3PzcHRQGSt2GWQMLC9EXNpsf211A2+uvO6eBkDy3m8dQZp1in2nMcQCfbZI20IV
7CVAQVdMEMZ9EXT0kSdeKKUazq7Z2aTUH8Wx/Jn7u7BfocAPtG4l2rt4vhi66jHc
KxaaF9N5wmtYkfJtN2l2ij/o2fiUUpkMsk/JXm3WFkPQuuksjbS8k7xrbvzecGH2
5REPqM/EPa+JqFoBgt1l+Qn/qnost5zZeKFvoDxIb8Wxe+PwLomEpiz0WztGWdKk
pKJFcTW5p9KoctMB+f8FnMf+q2YgaKsgRia3TWRjXD+Qn+YEC8zvfBMr2V498t26
bRQ+rhuPrEHstCdMtT6c53kwktgbFsH/RYHzn2/Ox4ry+GGagkHW7P/ftCPgAcQy
QGbJwXIf7FvRVVou8r6vaRI1KTeSB+2z991cKHNWje+Z61Cn/ZkI8Apr3JiRHAq0
jG/jD9S2oKe73aVDVn64bpwuWhQjlw/oFnIVr7hIHPaZN7S4/tjEPImUNBdFLLRx
c/JWuM/MQfgdSpjPSPYbtu5FDW5iWa4Hmtt8MXmOa88tyhPNxR/QFTMXkgJdKYlg
ytSbUHVq481vKOV5JgnROXEzfklOw9VWvh3Fd5UT2N82TXSE8gS8+2N9TmG4GUan
ENd3FzFVMgIttYOuIBViMt8psAXg/Ko/0m8GVQTfbZjWM6UOES8pWmUOvn/j7Sqz
mB0eSpdFPAXnEQay4lEkNU7FzdLHe/VAR6AxhfAqugCIhZ83/sYUIuuz/lUK5ARp
7IfF9UoQr2pn3FSmzBTodF/o9yaAXUXZMW3Qa6Rnroq/b/u/iBo8NpzBzDzbBYMQ
FjfSP5+ILJMNE4MJ6y4ZrI85Oa0aQpLL0xuL6W9YA2T5G6KRuKvt2Y1Nkuv6Urq3
ix70kD39zmAMi0dVfwAwUrptYdphWZcFBCuCGeHiH3efFKpH5XlxtHhONQGkUyy1
3wUl4brrmJ22ftrTeyMkj1MTxygVMHi3h/hUlNox99AGHqXaeZiUONqn9RjGPWEF
QsWcGDQofmWhhemlbqv26n7PycaP1ps+I7MTe2X8bsQ7N6a1pxAHLO3wjjsgwNLW
PgDoT8hJORW1wPWqegNXdii0FrDMHJqNGZgIfa1h0F/WtzAOyLl0DFfO6PYjDrl8
6oK2zy6NpnWSETngv6AuraPT+Zi4a5dCdQSOqoYb8P/Em5qMJ/X1xSYgFnh/P9T7
QZD2BOQyYNYDv9ZDQHkICUe2Xcx60F8exKKSM5NjXPPDIAHvAEifhQKOc5cqXtbC
mffSF7y4ifTg3ohUvh8PCKbjhTkgSDTJCm0D7NXdSF1m+lDWNGlXFOsdNTYS3GK9
NXk0s0/kp+mXkeeIfOxkttRHI2hb3SvXwUE8XEMPJ5Fw9Oheuzj2NZlJeEsGM7yP
P4i2G06CQiU04cdmXDSNjgU2zj9qg2yORsO4WsAlEQ3pXrlZSKXW8Y7JbamO+ufD
GbXM1F2fZ9K9jrAbKE0EhrBOPNduun55p2x/offYhruGXn7Jf5/Jp61t1a6+KceQ
pN+BfWpiG2n5WqRm7FxpH/zR25YVZZ77iagsLcieFOP6dw7vrNvMXrRafOfX1k4c
0QcviZzXBwbsO2srgL500IgXerQh2GsPkyfg7XNgeK4VJnxeDhFcWA+R7az4jd9Z
iGw/xgjspDmoMJoLLsGB4KrP1B5uajCyxGLm4bohV2rcua/FCbJV2umnz/zJZ/Ck
pmNHIWqDxT6v06AveuIk7g3avZ20iK1pkR8FcSmXaw0tKR6PssAvwcpM+GswEbV/
EiQqBGkxJXa42wfGDWIPHoJSCFFHhXPKAdUJKTFEMrINIeY9jUkPp0m6QA6NDR+Y
hXaX8YGrnp6usnSHFfHhTKGWOLT2YTc33duZ0D3cxrwKIJjlxTyetahKiGLSoLVt
dvKV11/DtVE3xxGDBh9WizIOjdxcphUh9+cXivd3JHPQjvrDlZnZLaIGQYNlWdLa
yV7V46fAasbLyYop/WBnEfllSZ38TChEcRXyqXrju/VEX7xz9ca3HTYFEcPQwJJN
76qNpUN4rDcsE//+SUU6yC2lL27DxtPPEUJHcGDZYt6HSzHDhcu8DLTcvG2WyfW/
4QhQ+G3SwrmW3AuDQnmKuYfftrwwG8Kr6egonjyXx6vVKGQG71KpenuCjK1B/P80
2u88UR6OUD/2MBC5ksZIyJbIlKiZusZL4gmqLWRKOLb6abSWxvtBkBoqaTq2tc95
jh3//6Y6awLx6zxr01qfAw2jEcWZQpt6Jw1E4I98EOjI0nhUidArcH0s6F/+G97x
tOQPpT9MeP0D6t7pl3k2od63ai5rhJzF3bQ275VJgQ20LX08rmShnvcYME6HQKOt
ufl841MPKE1LYqMQM+hZ0Gzm5D6TIJwVCt/DX78KT3oVCb0MrmVQ6aeqM17gJpPL
VHo2OnRn9oseINAsNTqq6OXR9PmB1P7x5pT00T/0jtc+lNyj640QmCUGQBSLIAva
jFRGxL68IV9Bc9VQSapqBWFe4dFYqNIV5imfa3pje74mG7CoCGcCFO1X3czU6K0X
3mn5EQavD1G9XRTg2yeXB9F0XbGYdSwgJPyrZf9GqZny4TQEnjFoyVW2Y0cZaQ5y
CpQ0x0/V/EzF7BM35xsOGONqAuNsY+g0Q7SBlpI/wYHgLGu0frXVKjjaP3X1bEFq
kQsOe55ItGyybBaZTdxV7DrW9PKpqUs56el/1AeKEPMw/PBaqk4N6rwXeray02Ri
zo1JN7Ot/g5OQyUoToOBe7XrOKrc6qpjX5oXVInngFS2xfwP8GjQ22R2mihrDXaz
plEFaang8UvinuhgU2Ob5cH+4/FTOiihqnPkL/zW+tQjQp+jWU4+n0BsaCAIZxWg
R7AQcy7Ki5iJCfD04aVrmDdSGyrMIEZGtFODDlfp2AADnX0Xnl6PLDeLuIJCP/8g
si1W2sSZNLzNSgOzpHuhvIJt4bQ5NTrZq26B1bu1dhyWsvYDyBDaiiP+ve+6iN2G
U9Zv/QTD2mgBaQ54s8IK2468ih3fUtl8DzPMi4+0F+Z52OBUwh2/vJ0rEXS20kGN
kL9Bk3R75e1hTFSd8jyjWqCvvm2/hQxVBA6rATvgwaDj0+yvHv4ByLriTZP8FT6O
PvKU+4DTorfIpYu0ktC6zqQC5sNKNufvATwkSDqzV/0nXO+Es7HZ6FNLLiMtLKni
AHUbDv4nu/M8C+PQfnJHhfJzXxcQiFMx23zjcvYv16GTH0Ykrciot9SnvwL2vQmj
cGZyuIaQy6cK25l1bwWdzzAiCEprwAGk6WVKl0EV0A5NCR5+9P31qmxALsm/Uo9+
z6zuy23WhrSm3IEone11/pDhrwbbbpoytyRmQpzP75ICNUHgpAeAr71t5b0tZZbY
P/nOSjWYicPGzCVz1Wbaqf9TmdcCkaoaaWq4q2xi14bh1Gifl+q8EC6g4Xj1wLmf
595vjhwlXcxfYgrzUCiItMtHvxGt/S/0d1BZjjIQPoahzVx1DuNgKpXFsHVqcUC0
sXbYKOOMZIvm7FWBBoFbTs2jyoiIiJJoUD0jvqS38C8lL0DyApNm+WnhWJb2t54y
FCN85u0g9h/NBCKdrdNwVEF5UfZp6sQGjrtpNZ1UJgBdTsvjJiqZSqhMM52kP/KV
EgspqPDqTHyJUCpuiXqMfNCS26t15vGXReuJBeMfIbB/IW3cWPEqKad9Gu+j+OSW
gxEL1tuj+XvU0KNyz+oV2aaXOnBjiI9zV+62vS2rYbiI4smy1aKqtO4uEQkZtnG8
KQA5KtuFHkGR3YPHt4q40ZW3dh+AsPt57t+b8o/mNFcI5ssYKLxzCG4pxa++VYDW
zrNzIdCSRHnTPc6KxUFDkE0eowXagkOM6LOpvQH68m3JmSJmXwRHP/tXb61LnPgs
xzrzau3CvJPaNGKfbzCRE1YdAo0YnunQsCsjnVEHnBNNfylmqZaMdvG5/t+8xgq4
NY4GUUfDD8js1x23qaV405JuAFCM0pAdXSJmB6OqZsHbfWwwiOKueKVfyGx/89Y2
r4nY/Oc66TF32D5NhDJIuYlI65QiLATBq9sFNzca0ZJ0om3Iqq2OShL4m6S96hgR
V/eksDkSLhmkJxMmB4oj4RuFdQ8aSeOl6Edn+DKagn3C5863Xxy/WeYP3MHvmcTc
fo869RlIO/fz6d1UQJUAQIUchLsVkJV1sSkIQWnGFKGhDzZBKc6PVWrpgXO11Kve
ciI4TcnIG70BMq2bwi3m7GjbI+bqLCPokfj/BwMqyB66hQ9KW/sX1Izt7fXT5P5y
Sm2qgWfFvi0xy/cHtRtQDIQ/NTRbce78MxGrSNAcQ58yGzX3nf++SuyfO8XAgfaO
V41yz2w6eFvtEF3ADCqQsGt/fo+JnKRuRn1mfJQjCo0Nb1k65F9f2WNuRHb9+rGj
mHsCcmJDuIZeVZPijIPkGouacHlFXjh5ljfmFtwLjedtC9SN/PH4Q2w1yv8fhJla
C9xbdabhaO3xDVHhzGNSodOj4rUMo/NhRzZqkVM4CRGH3M2Sxf412TVo4J9aE5rN
BSD/3xlKhkkJtPVDvqnRTrmKwpmZt2887BWM8328a1lQZEu6ypRKXrEsSZ8oLuNc
hxWz4v5fdpBPynjydJMyfYGevaEtlpBPVK7nymgMcL40/pAOxZIwcIZSxXJwYVWN
feAFthOuK395G6B0ufp3YQJzs8NTOSvrXwH167eW9xPZnoTzIajGRy77r0QTWE/0
QDzZblLmRBX8Hd/T1lRgaDXwejh3ccP7O9tUjbr5TR0JWIk23GFoWRfHb7sexrwb
2fDs1GHYHeDnSzjSwwS1LabwI1JTtpS170rw4XO2UkgGl5WlyAVRBIIgkvGqZD8S
XUzRiBqyuq/6PRPe15aADmjxD3VMBTfCBS/qlENp/rhcPILTY1HzHxCruuxKW3zh
YY4Txsamc+xxN4ZZSNjB8lkUgjM2xF1WzG8s5J5qNs6mR62walEoWEnSGQswmfQa
reQeZpu4f8yvZAGRN6gN4hVU35YpMKHAu1VxaCqoMfRNvkyxH5lt3BMKa1YMsBml
Wyiawf6VR6GeA4jcUhjmww9pN1Vyt8UnSVcrGI9Fx+JaBrjsx8qpMbwm0pTYicIs
rGcZQcV90ImwtCBRRgSrstHC5DMsvp5SkulU3DYjb4e13MwAbxUG59AfWpr7z0/V
oD601Tar0NTL4JNVLowPOHAL9OY402ohehO2c/IzpNv9wHRy+2b9zrQyXaKvCu8N
6EaubQQiIP+15jnNyWNMsPPHF1FDjHMoTx+qQlmL7Ml5LvnpXl9Q3q04SXUG/WAE
mWWlHl6VurNMvYW4xtubwZZJ4CYsWtfm19h0aZkYdFLEPZ7K8jp2y+Q7k9akLJsd
2kr51VrGdYTFyDFnrNbAILTSB4yKxreQfQf7zbHH24+UAKEk0mNZD4GcrNoIpjb+
7MF/VVeVv0UBHmzTwZVwWLdrb/sgX15AIgJGK0cLnTJF0vBc6BLPAO7MkWK/B5Ql
FDaLQ15h7xV4oQ66WmkFnDgnQWPDWoMTu4aBe2ffHrC00Q3wr/aRdZd+j6O84lXC
Pc6BGSYGl9cXgJUghS2W+nJSZHjHWS66KZLjmw1viMI86Thd0DJAZmspkVlPAPgB
UOd8Wgr8tSZWXjvEpT1qqoo0Ma2gZirTqqOpMofcicjD5YrHBlkDtblpNra9nJ/W
Whvg2UlXVghzVcxOBNITUMH1yB9rUkMd9d1epsjixHSpf+QakEIQDwcBZ1B+gNyV
d7ZIiEvyZWokawpcgRNLOpGAxu5qzILJD9VM+b9Mkg/bcfFjZMSIwZBvbpUTzSbB
V4XrMLNs87UzJ0JgpIj+M1xXHMTwFwLF/0YjYNiV1bRBzt+6Fx6bjBNn01rUDZDY
t5U+plJtWw764VbgDa88W+4zeBVvbjc+NwZ8GZ2oiXgiB1JGJdRvYlaM9XZzBtQh
5pvJuZG70cfImzsHmx/5sMq40fjulSUHP9fkHsM/RsTYjgpJ0F2WqO5w80elrufx
rCcuv3Rh7AAQ9fuUhuCcdbHhOQ2fg+zKL9y/YH89vVakSw7pJkv8JKY3vANy47Gm
kIXBis6Sg5NkTF/U6Cgzpz0TusDbFo0Zt/5NjsgHuvVaJTU7ytqPyj33L28XBCqa
gJnzcnpbO8Tx6wfX19jCyDvSsK86sodlA6pGQvsIluCT4zRnIqL0Jf284njDjGAB
AN8i31e93Wklmr5AURL34OJ78sT69SuhrM9fC9ZWR1ZDNWhaTDnea/oroUIK88h9
BaUUwSCP1AGQlTNUgG3zbEoMTU0fWiZod8N93WfuWjiW7FyX6OJBhWBpcG2siMMe
jnetoYwzILFpF8PHnLqmpFfpj0GCstuT8kw1uvKZEweTfaJD3F6oNa9m8uPGJFs/
KQSb2don95lHZbmpfhWm8A6SQCP1pnLVVnLB0fsSsFPgn+A+U22muRC7jRQltLdO
us0eLU+e1eo9ArWrZwUzdYfAxxz1r04s+r6p8PUPTPlSGFdxehOv92ZQzBFQ+KIQ
7N2Rr9Aw4nLcSXzgJGoIPPVQbVmy2y3NLVN75c6/5chCay2OsyGK1Xtkc92pWOQD
tRJB51qhvClamhxtqst6DR9f8UAe8QUzzQBzwyDC3r9aByEb5iEkHkkceHZDPVnV
dfFZX8X/Pc6p7qRISmB19BcjUiJzHKd0y3VhMBPZaoJqVDky+HObdUbNu8CO0kHI
Lf1VyTtKJ+cYtQ+b9Vjlu1R7G7jQGmVjqAXzY925VgCW7bkb1W2x5pso9WkS/emd
Ol9yAlDRJripgA6Gj6tF54It9yAioddxHpiXMgyMUk0gHQvO4thuI5iHjRoCaqLb
diMTDRNYbhhyqe0n4MBjAqhGWPis4lqIV7NpX9xufCZ8e+ZnFaZjO+AS/6KbVKkq
9PK5COwcdZREWhLxQEVY9+Mh6oSf1plUt/OXeeUa+IaIRkyHzRzRaagQK+Vqef6N
j5+6gYrCEkKZsi6aCjqBKma/+I9R01ximGL8HiJhC+5P8a2+ow8ujKdx1tuiHzcD
AxqINE32y2Uis5yesfrqlj9QcWAW/y7l7T0UI6+s+YyI02O7I7nIX/eCWznnU9Qq
Bhoapwf2hwJPbgfPnlbYu7IdKA9tSecas/6o8W/55Vru9fxnsWrVShntOE3QfulL
jDlUARVWLwci075RQQAAPHsK4Hog8MGd8KJA1G3lx7iv8jTAzpXUqr2aWBRfYLzN
fpQZaU2iXiav5qs0THfLnbTXcK/EsntwJ3/6LrpY7DyCoPxzJx3f0+gQiFw7qPL/
zT72BcelIU6eBW4WMyMGHxF9Tcb1E217tCzqAhxQfV5TSNIszTs/Ed+NQkMgvuuo
ZvjZGpXwWRhFBJKzfmM7TNDJtiEVeeWC1/pq3CofbDcw7suJEUyTKx9nIfDEqABY
SZx4BI16LisSbUC8FHWYspgnWQBk5r5M/NmT6tAFKbTZeOiH/dwCFOLi4BHf/4gu
XYKrlbCkZAzAxkyoYKJh6cE/azHk+3SpHjR5uLjaXgUM9clLmI4qTdb3+bvtXe5X
MkrZATOyy37CINy3hOrsARO3CG0D+5gi8kyI/j50TJfLwWKbZn5lgI0Cxffbn/7R
ebY5kyldR9lXktzQ+YMvzmlPVSoYc+vqM3ejctYxPtTvNF6c4pySJVTVwJvJm3Un
AY8TElHDXjTi0PZs9rEf31Uei16mFiKDp15xDldvUdOz3C9KKsjV5tayrVuqcoXQ
OOYKt6aoDXwQDiC6Cykd3yuxbK2aEa67a+ukKLd4BrrWfYrzwkyxkYXkgE9mnvn9
1oybwdbjfj39k+qFFYKuQx+Wip+CnN4lqjfu2RlWXsewWNxGLxK4zjjGOtgVLD2h
G1lJe+yMyZ4IgUj8fpFodcPJ+UEP9Ya5+TC4eZeNz5E3pWkbxZY117v1qOEPGtAG
4qqJoP5vXqH7MbgeROz89p4pNK6DuaWw/bbDNrH9frKaWAfgvII4JKY65Q6xDe5K
uXB9yxQMzxlCqUpxfQhLjy0ZVDTBWK4Aoj3py30WZfqjq3eqQI92sAOlciEB6IPZ
TX/4ETZfw1IfHHdpGSjpOedNakOh04Udu8hJ7EbBsAZhAbBJKItl3SXOaWmuOhy/
RYGqLO0QyFz2mQkXdrYJHB3y1IxmVFheiZl+BInNYH5ObBkeoqOgUicVfv2uYCBk
8kchUkx1rZcnrrd4UqhqwuoEfHnZ0x/PFxQRZkimfIZ6ed1zeTb2LhkB0iXi2anv
UfZ5OjX+7No6ZlxalmCCOQh6GbzkFu5h0+1VLQ1Du37cUp1X7ojtbRi0Lm4kN3Ei
lNIVaTA4E68wSj4JA79IdcETSVSlcKvu1HP6229R8kraL6QZ3jp7Uv/+/bCBa3Oq
81RK+IeLHFxTPxr+zLNQsofC1RnLme7kN0VcOSRHqHUoCGUmBoiagoUi1l4iQ4Q2
sYe8Gt9LAhzraZqj2675G8B52FNqMzWjnCZFw82gfsvfoGCaB3hQtZzsFNFLY7MX
4KB4ZnWNaUb9Z9tVwZs4kBnXL5T4SxhvbFyUt5/DqaFTPlSEUh/0VE33jU4DBEjI
ZqqiuHzwfSeUDmggUYwg/nE2afJ8TcM7hW4RtQzZx9fLT3hyWTzjWInu8CSLdXRe
x0evhnmLNbtwbB9ihk3c9wguLxYVpRLr3lQjI3d5juvIdlGJ0jngp4AfWYCYDmVL
7UsaGrBgmlplmcfUT2pUFKgJVcpb7S+KzNWPcOjyymIJOD/hWxMiE4FiALPw2RtT
Ghg2rOEgTEpK+shLlimRZaQqkKEYQCpkiPtL8ShdK3I0CS1E8Z8++J5CWEkgdq/H
dVVrKDU/hiumcRGW2bnvRST+6+9RGi52dp9gnNUawLuEcbrhsEIiit15V/zSoOKU
IsreNVvYfWRN29zcy3Vn+rFwLSCuCKs7o1U1Dwg7SDAs9O69xUBNKwNzbps2GOq+
wVgtSNnI353sK79E86nf/25tNirmCVlAmxS9dVq27aLMyeilXVoScH3zSWRCbWGI
Ed34V32lS9NjBLi2X1iEy0n9iyUfz5nGL7nWa5RKzfMAVb7tEzWYSe57CK9O1MZd
st/cBOQNFWZBCO0msbO1vjADi6ooGSkEtgrJvAGBcVOE/eoZCMtDA9By3HL/Dphf
6OKDCGPHeF49OXWPMU8LGhVpof39iQCbwCsDkQFGzsvd5XD7ZWmiP1Tm7Vv1hTbO
oXuDLBaeyJxjK4tN9fKJ2t3I9Lik3MVYjkOMyitI/SWV/TUYzi31jVElrlsn6xJj
KFdOc2VdgX/iJpbOhRdwKzbmXz46USGkldmuUAyPAKdJY19Ry37xnGESr5E7PAfR
CSt5d7sZwOFHnqa0uOEHSTUsbLdgRdsC21FSMBb1NLJzrNZ1VRjIYR2e+bKmslMa
oXabL9AcaK8A5rySVA2lxZMuWmUaAos2J5emliwmwJiY4lq2PdC6X5RUQHflMzte
5eFtl1PeUJne2QoS62P78CbBCAKaKPxGjLjHMjhi+rVJAJnyovZnCu6IG0AWyisL
nSle8ppnbUh5OB8Pg+tWGVpbNnaJH8j3HuLgp/ZUJcloO2cQfneujqKeNqKyJCHr
BQTGuuCWxKm2HDbFiclI7l4qe3v7OdrOoZoCVTc3YsrBRe/5pJfBt7CQR4iSTb/2
aHZWJthROnMdrV5oqymDeCXdLIagpGCzqcOL6j4/abMRCY63IW3nkilKFJ4rcO6W
p4Zk6ggV7Vu/Qv+Nmno+5fgDJt2O2HzoPveBVfWVqzFvsJgNR/pKfOUkCMNQQaEq
G4UCaSMnH6FZdtyV2zCIsYaH9BWc7gS8xl5wvLUvl6G4zbwGm6e21jVATLk3EM6r
+CjrVAQ+nmnLVdvWnpWmLaEhSVepiy3L+ZPPEBrCeQ8Vovxs2M8OPUcbIwl6yOZI
8mi6bR5W+c02EoadIgQDNqxh9gsW8jl8KgX/HiVt0cScA19tMp00myIuXNHMNeQ2
fpDjbrQNege4dMn5NGTeovFThvPw1SBj7MEwRh4GoJCnoyJaxS3wEXya2M2ts+ZK
V0+SQaUgJqy5E7dH5kuTo3SuxSOb1SM4Ht51yv4r64Q0MMbDzYpA8yKDZ6qAunLq
c/ZZGFTXnq3Q+doSa0tIFH6UPFbw/JJSdI8Zm4HJMcSq6soXk5kO4X+m5+uutn+x
kdwqCEawa78k0CnY0EAEdf68vtMkHaj+KSeB/rUROPbCGVNKjV1JITANZflZYkXG
PgFnP3NQUKSfO2etf4F9BCzU2FI9FGpRZHM6Ubt5hpQ3c9vHbwg/a9NhqQajCihB
N9HezaZttYuZX6DWII0U6jz0DMcZ2I6cIk9p3lBnjrLs6geYBmRxhq76HCNBvwzT
uNsQfLmuEVTeq8mbZt0bKpK0DzhmQLpBk0QbdiY/o8wB2Vg6bt4wlq6RnEWR9yH0
K2FEZpixKxWub2uN+SQ206EvpgniVkhOvRINf0FsSB1bJjvNL/NBmBMsuKZKptO8
S+2FSOg4pgfbNHDxb6y0tm4DjzvGvFm4AizncLIo1+nPzejz8CqIuzH8rJq1D9n4
kWtkamTOt7PEl+VYBqM1kYhBTmlITxBavntwaMd5qhlM7ShlO55rdAiaKq2nhCXM
5qksln87u10MfFqB7+9FzKKoGUToK2jWT+WKbcv8OSvRE7vvkLJcDJfDUgDwvb7W
xbQZ+f04aQwZCQiV9kadAnJrvbpidFeJXCjjdv/6O3NfSEsEeXYuvscSZWuzH5tI
wp6K6eJG2VMhl0O/yGG/XmgBoX/BfIixfkVOXnJBcty/rGQq58zgjVHV7s5ool9y
sCf3ynNkZmrHqKleU/jO6nZqxuBnE0nLBTUpJEC+HvNPz6gdIonEMcD7qhZjTXNt
LPIaubxJnKFfPKdMCx4ctxpaYMLXIH6kQA9ENDLm+rkByITWAseA1Qa1WwzkQLSp
L9oHFbjoFj9i2ajPjzNVUhVm9xR4Xlc9k0Ky4ZRklTwVdEOq7fr07kVo9ZArzf0o
e46Ne8JW2TA+9Om9fdMa627IOf2bF34GI2YrvSWSr9eFNSbf7LRhiWLqO6y+LATJ
w2LZ7Dqsf9LNhoxaQfPXkkeniLacE2BUXMR7qwNtXq55v1s7HX0X1wv2JWcvGT0m
UnEhN0M3sSBR9yAOT9wDFOkMQNcdAZ0E8+2bDGzbS2jX1z/nLOnBr/9/XJpVxf2b
HoP+jsb2h0++ixPND7LoUnzcLrCEG4642TkB8NP9POE+k1rVzS2HTEOYTCaYHy3w
ls3Mjv31Kf8L4ehLt226PfKKo6Ly8jADsgnuTc+KxD1zOOfEotG6Boq6usd0y7Le
jEENplxaFfMS4gyQsTxQPFn87Syj5s76z5saPi9jo+/ooJvI8QRidHZ7oZUViWDD
tDvLGWTjk/Mc+u+SSPTi4Fu5n5Epa8BjW4yFciLC75QaMBH0pDPqqWDArieRsmFi
Y7YUA4sqzwVBmhBH8937VIw91q5YrYyAdlIZqU/BE/BqgGrl3QNQMwX6wxzRsE+P
MDK2GZy8fxVJOCREtsEDtZNkH1hz27/rtg2VgNozzAM7LoO8pw7OZrk3jJvTZ037
9V7WG6dwfhhePNe0uADSfAsKe53MXjY8d3K+JpltPtv59DfMM7+9tAB/LIQjEN9p
boB6VKlwXZM2a3jP2XiRnRk9I4eOk14YU10fhwxvI5DAoVUnT9OItPvU78IcgpVG
EubwBgdKF6Qmmd4ho3S6oCwN3ZooVnihntxXAdsobplDvlQg1gzxP6GaviF+Ta/r
JY2vO3hMxqkTmHiGKqc9UKNaRIukaGgVE98QCsmUe255iqYM4MIliXKgazcdZAYQ
Rl9JLHU6W7Vj2qrF3/jiliaXytlWrvQROS9JxLN+U8N/puPUtVnLr6W2S2OATHCG
zyM1HpYHcQsKhfwraK2U1LfsC+VvM/afPtN4wN29W3ADaSEUGlSLgX3avFpulfQt
eWb/LvshpIZnokbfl7DJLrQqUCkEXzWNdoo7O+60aGiO50iBei2tvXTXN5cx5//h
b0QUiJ31fV9/9RkDH898a57MEk6R/fDtjBvJlHrb/cmX0S1Imxb+OpRVc9sDLIYC
T3IEfAPkiXd2WFuZNkESAARPqFRc71KA4d3igGmSvBI0LkfDwA1zXM0kLpVtAIls
+oxN+6TSkHsBE49KsW/zbo8vKLrDHkxOsxaEV1qxOsFvypz0Y4yB6LkKlQAvL7bD
VlxiQoh6Gk0g0iVXRoxpi36RA5clJ0KCGVy3pltBTlVZO0yfkOfEsfjrbtr/7C0I
65mNmvSmI8oyo6UD9BtgVfXkeCAw/km+ATxOq4cmL2w8aQ6jRdjL1X4zB3wvM492
poQ9WAwosSzkRM3w074vOC1YTMfMoTA+hSWSE/tY5PUoIoZMPm9RDlaDy0nG9UnU
F3mrLCGS8UAxsfrkZO6o5Et8u1oU6IaSvDFUDhtZI68rzSIZ4+alOBooxcogFNbm
A4coPov37+1CpyEaf1HmrdStxg9HRFla0/76S41QBEqtvZyXcqt90bA0RVEPRGa+
XpxHILedX431OscdKk9JnCWxumGqZEf2ZZ5I/+RPWhBbWB5xYU+bP+SUf7zd9lAC
xSFIk8vm/fJGzNPIwLpQ5GeiXcACMB8oF1lJMrknv5zvGYq0//6esjvZrWgUIfIg
A6CcUgIP0NqS/GLfn1wCS4VidUloZq3jONO9z7BBWQB6tRUodPuDS3363+xdY7mu
JmwbVfBxrnMLj4g7fz5dEw/tmtoLJ2KNv26/yFY2c/6HSpNCeu3zJPTdGDdcIDGp
tFXvttbuPqUldCrHuN7xUBKFyD+DqFREm0nigRg52k0h+cRCEmd7B+mNbB/OhL51
NP93M0XAIxkpdSIO0V6V8bQo7Bxs4n3ZWfaVw5i/2L3C/gHrPkGChS1FfHL+GfIn
UCOh+g2Ge9VsfFkmGWv6904pyL2P3WjzhcSa75aMslVj6VWqAQ74cO6zu+he0j7W
0YNV5Lt4uOGPcsDvp8ne41hNSxazrR0U+0Rkafqw6N1/CczNR5m8WVEuG7tTPz1w
9g2Aoqqo6Fq1bbI5HxafuuQJd0AfYxtR1MvnKKVIuvA7pbvv0Y4ke3sVcAmHkS2F
KrsfDdyl6JNd78EL4chUrPaH1Dh/HTH2xHTOSewx5ggbWto816txoyf5Rzr9HJNs
tVoITxHNA3P7WddBAe7KBGVjgF/3Jq+FejDqgVI22TUEp69NjFcJTWRii+w+fiLF
EvqwrOFSwwlURbEFQj3Peicv09hCc2ZOvGE+x5kVo+Tdrz8roecugBchLUpIZRqp
iU51f7wbsFAWym+TrYwQqDcL+VwfE2nUfoe/nYb+UjVoCuGhTdxniHuLTIGYi5FP
JR7HKNiO2mAHN/akG3MCWPTIVXQp6kIZ90f1+bJQn4ByoY0oow+rIugI4RbHc3zx
ZV3K8MX6mL19C5fmc7V8SUYBGY0Dwi4poEyiQQlcYoEFOSNbiDsYnuaLIEScQcEi
geKKkoFxop029tzOTprqDhDfg1AiIeJrTc5rXtLGIoFh4++Al8ACs2cp+hssS2J8
TEj+50EzczVRV06ZEp++Aij9YMrujmaSC36LMiX8StvRFvtf7Kp25xlhOTaLfP1E
P1/rQcKVWdzbIRIrbXXeS9WtSWJrroWlrGQ4rnyYyJJVIi1SO6D3VXh3Z4GDJ56k
oyixY2KvXR2HvLPdPgan4qRDrFWa/IZzgvk2bvrMKOaVF+wCaglNhWIliPi1ctht
ARPjmWlEPmjZJ0PAf0MTYbvKloy4kkaAMjxsl7XSQjv308nGGsxYKkJbomhWDRWi
zz90RgD6oo5v5auv6sZCNrPWsYWHFWcANCcN8aTkd8+sdB7bSf2Pm3n/JEMpJl9w
uekhnfJUDhXofIzQGdn6qqPQl6Su3NDcYFvcEQV6IUWTGIjsgsufzRs0EeB9znpc
nJ1jCzknsZR7fI/C8VZn/4v8ukK5FO/nLox5KgNcjTneERsQARtpGLhSoppf4w7A
4sPCzOyff4wVw6EsJwir1m2I+pzqJN4xI0v/aXsZ8FTyv1YHbqYdqUROf69PrVdi
pBIhpo4tN6DtL9lfkHEdH1YkLHcEvKOBu3tvWIZPic6M3deTSQZKUY/HUbeYwTOs
NW5Gc6H0un9Mw8599x66vSiBaKZVDWWoAAPbDuRfEaXjiGcHOdhEwbNCfwcnoxaK
4h5+JB5u3o1VfctMp6RfyI2MUTDX3fcCkamhEANtI4eiEZFFcbTjhCfoyY/WxYzT
Dvn0fzwz1utbML/hsTbhezujyGKAgFCqPpwQahVjVsqeSdr0OlUkya+NpYVjjAJ+
8YTN73DW2ywegYt3Uw76BZVaL5aI2wnKywTHpraXyZIggpuAA6X5sTCOKJbIYUSU
7cReUNsP4dERii4M8owco+sc017z8GGed9R90Ake8ldntTbf9ySjG5zWxEqoFmVT
8TcW/lPAfC2OMe9JgT6MSR7wSbAVTzG52/9Jpsh0W66Oi1rA4PgVQy4EfL7nh9Dt
v6OVSNg0D96ElEUwdqzo4crh2uDiwKwQXQL/TSCl9jxAmkJujISq0/MdzWAByaDt
jk5zyVCYCnsnytrIZ75rB+Xz//IvVvl8H2R1hAvsJH1TZx4fTT+f5IgdRTRXhG7U
X8fZ5Co5rVEhkjhCss5fJH/66IwTqsTomXqhrApuCwOfvH8NPN9/f8Pd0YXMKfiS
CqbclUSXn3ieJXgPBhLBVm/8AC5iQypQPGiWrHVHa2fNkydtq5CKa4t6o3bY1ndm
1Xq3qB/lMQWtQQh5IpRd+JRr2tMQg6cUeenca/rai8eJt+4QGA0s3iaMB4A5fc2H
WYYKIUKZGSI7Tl4GkBoVh8BheL8mP3CymF5qjlIfBrojqPqccvKGuS9ZLg8h1AVw
gdNWhqlVFAZIbVDNEQa6Ob3kkrk0uwmbA8tBgCKZJwjNc2DF7+Sd+36f69LFQMJx
8DYRuqKm99swNfAfwHisqeR62vMa4gm96tiujmd6724Uo8LWXutlKfqxHogx/2sc
Fyxi3PbSivkxdt221ri0Dg66v3SAMs+tjXhCcY7L8+xEU5UZ6oRveP8BYRjpSanJ
Za25dUjJYGn9JTDH9JwavuYysQgVhvXmit8EG8N/g84rLwZTQuChDf2p+nwvv+1Z
BzH6xGY+X8w96qF0pyR81HiDnnJRhJNPWc/32EujyCMhEJnCH4ibJEvjYf9MlGNz
8/EXQIzulYjst9aL9HQHPct6PwVXvk3hv2bbPwVHeNCQSOGv0wbfcwggjFl9YqSY
0cGz+ttKnbwGIJ85ZU44Qjvi8057KnpFLh7AccntXh9kfVwrIbVjNVM1IY39VOys
5VnyvdoJX+1jDtYfddmwbH6ux0nXP5Iq6aVMxgxBk9tNx1u1aZoZVSYH7t6oqNgy
AZbxEe3iME9RJVXt+VlzvodmWH9VAjJgpji7TluWVAqY8M76GJEAj5Pcqws3xTh6
SE7h3/PLkJuJ0q0LCVC9xxkQUVrhmQx2gbEPl0qBd0Izt2nqq8zEYcxTgCIdpX1o
tgz804nx4f1JExWX0HTB1fIWdPsgEBkHc5ksWTVfEkc0RNC3Ylr6eXRJqHtsHBT8
PO1vrHDWkaMyrsvDrhByCVrXFp3+ebZg60kCnR6C+EjXLxEzUtXBwceAnIztcpYq
jOEeFaDMtENk8Z9uP4pmq/Qfh7ez8QbEEFHmAweLqWKRI/O0VZlPU9qh/ZELP/98
PPwGsP+tCaT7NemXobB5KW+qpf80lg5JMe9xF51Lnske66VcL2KqFsYRZ7Wmc6Gf
eykrQgHPtMhiA1ZQV56QRxl9gbLG6WW+QF6GzPrCAj/zvaIIIKz/T4Ms2h2VdQYe
HkqScHW8G2HSDyevPvRSOL0ljQ/EfXje00J8mpVy7fTXeeCnoPOds5EXAQFKjrg4
HNrpsOrC0eGq6FtPcn4MTLWDw0JqJBSW+fFzVudVPSUdL2RWPKArZoUCkrLOg052
TS84HK9b39Fszl5ZTl2SBm1029k67+2ov0pnsUbb1UGIb2DNRhgbP7qbcmGy2Is7
6a32GJvs11V3cTyKJ/WEgOG4m8l9uP2/303jfJinpvIBnYZfLArHodB+7IRSsdY4
O+bGZ1FJ3mndGnLSGYKnSRmj09mjTsHk1Unl6SFtS6lFPATFdbclDa1/YRCqh0fI
WG6fUuSOLTGadOQXUi7iOjucCY2e+kkyPjRPhNjh47Jg2BlJI7xKC4jF3V5IQpfC
BSl4GTa8APQ1xyLDBQP3AtgJeYnYU6YxQNLxKKAY8CPo1augZiv5MXVrRCZeXuvm
9og22TjmVnFak0xtizrouPp4OK9wTLXUlPiibwwtzu80OVz1iw7H06SbhLadMZS9
aaKUhQ1zqlbg7WQQMN9eeq/o7YU4NbYhAVCV1nXAdEX+gzMTG9HDYlo33zCENW25
77viV40Ib99gwNEJUPHYh7JiEarT+RW5huHC9zHxWMvKJ+N2ymeqTqmVjSxxIp5G
plVEah8QK59Rl/mLELVvX82tH0fl86JXvsrdqDDxmFTVV5GTAFuX3IZHAP76nnj0
0TGw9EsH4e1SyNVADf4AIrIqd96bpAvvBEoyhfEVtjqFZppIhR44i4QzxlA4DIyt
CGi+OoPa/xYuv9drk/fw/wut0c6yo4Xn0C5rrnlCggHJWwCxwBJS2CSrwRzPHCCH
aJUJjYdOT2vmbr+EwUDC9QHFeU/Jz/qJqgE2j2ew1N4CavHRs/cRBKeDD7s0l8Yp
q2hIlfjXVSfdUk1zjPAU6f1+PYEgWdCeJlojveGhOs+hsO5bvzzJkwt6s5RKrlZF
qu7QCWVIsV1AL+dQCvsfJk019TeOlZ07Q3jphI30IwyuxZJfPW+43TjuuYXf1DSx
R2dmv9TY13HHgCupKqAOkyRK59yGZR1AiFC6RtyrKEfwk6DyVpcYv/nxGVFeTX56
EuVyhBVFXUCfqM5kAtd8oQdtT2gvjvc3VFpxKQLTvcs1Lu7rPZS5adyi1EPuR6hY
MYx1sJdrGrzPXv+7g9gbH5HAO8I34kUlSZrEpzpHrRLKlrVgtYO/hjJD6prD4tMl
XcTdi+SHNWcbL6jVncm+lWA4NmtPU6uB75LnwdETjXHvsPFGHyUibtWiVgXKOiZe
HuTNbdUFujpcrh9GctyW2xSIxc34l7naloYLMFsvkLr4g3lkAufOQol5HCxwMeM3
FWGDhvbDzcZQGrDBhjNYSi91lMroJ8cUSgsmzQrh0HF5Lk8IDWHcVIwjJIyfydH8
Z+M3MLUDkdVzrhp6D21sx1MhiwvLaEseaXemreVtS23Qz4L0XRw+53ywk+arkToY
7bbGtcD3h8fdnYiiD+CLc0pzpIc3s7O5UaY5IM5vu0cg8BvvHJl/evNDEFghfSGW
9Wb0WWrlcyhgKDqj85IQM8YJtGDa4mNRrl26emWfZkvPCiYG5Pv3QqYied6rfNoq
3mcumSA2h2WsVAOk8P08X0nqwzblTzDWMFW/9WnP0JjC9THDPFP4mMliT97knvf8
N5kLff3bCQfA4WnlxG01vDDAqxNkOStVG1X/UOFEJ6hMmoSJunBT3DTOc1xoyfsn
L3xfmWARJNXnAtbtfB7S2hmm3GDgjz/CDMtjPxdm5IpG3ma9RnTa7UvJi2yJGhZT
2b8lLmsUmDC9Rhc0SSE2ST0R5dklN0Q5M9YxRnxh/aWheYo50bpJ2ixI3d1I0w+K
l7nlBEgSy4OTsv+AA8FyVAqDpwnRJ8ahZQrtwtS5clV1gSvFTUPEx+Whyfm4Snki
q+0qegkpWUnoZPCCWMkpvzVIm/KIL5bXGMrMT2+VvR+K0E7xPzx2cC6HkksnyLp6
ZobCX1x8kFytOoBCPOfCyeIudrXqVk6zWpxtrUC9hKyIEdD2SmI5D/yCqUdw8N/6
6PchdcXLyolav6oZcizx64S15zur7tZBnoQGmUwiN5ZmPlxdtI4x2/JjcxzkaxRZ
KHvOBFrrcp1EIyB9SOmXYJqEYK9+u0jBKwAlcMdIWHwqukCtLPgm3UWMU0Yt1Ff3
OImdY1JUTpoj8IhYVDxtld90oO/AvWj6bbUEOUC5n/iaSmmKi4ckDUWsc4hl7F2L
qZ6AQtDqM0zhLKQY5GnLjR6G+O2OKHncekW7jigZ8zKLQAvzw4pp7fkDW6V3TYMh
kkkgv7KUxbV0O/EFbJGbcGhZmUTlGdrAG5pBTOl4XSkyXN+xqYnihTAYp4LlgF0J
8GMpj8DZP+yKOKhRRGNM/n2fMjJtDZRVgSJ9Om4zuEdCWTrWEkjuMYlZeol4UnHG
aC0EUNgBB9zibqDub8g8z4tX/sZv/dyc8ONikIVo9S/jrtINtk8iRBzTt4SEE7N6
5FgrdzYvzbn3O5f/4/ztwgH+rJN8MkXd62IhYtuYkGWCzkhxP0k6sTu/QnWPVgpZ
uwfhlMCFbKPgBG1n1VNWDXsxAoKWaFtqHpui40kxMTG+HsfBJmYzekVy5GTPEALe
z3YD4em0B25Di67JlKrTGTSvbmHpjm6XPuNYae1mHyXxTNdLxAQQj5x0F407XeS5
spco0pFsoxTpORmTWSeibOacNQvTwWr+4UxMBB8pYSIsA/utXagWWJOo8QUqEu+g
re746R6iWwUAbj5u/I9oSm+3vueEPx/6HCi0upxCKi68CJt1cKt5Cx62kIlWpc6I
iCQ4JJaW+iMagEoZKrwJxhqxrxp9BT17Dd7LBhKOm6bDStUast3/19yDmwHgd8t/
iNvDps8UI0fmaIyEHcDgiZBpdbCprhCYKBVwcCbLyzT7hW9J/EOep4dLEGfYmRga
2OtWhFxZVgUptjmJE3boKDZWKKLRyrfFvyFbx8JGeK5OmTEgEiupNEkihB40T4sb
LEhA++gg5QTzf7jV712DRec4MuYrQq8LMJDrEM2SwkzifmjKusd+4zaj8qsV9k2Z
3sZ1W0+fuUnBSdBR5kSSzugYBSEVR3iJpjzWIBfSmdzxPovr3tUBWAcG315QjsLv
DlhTSMq6FtUWSHZnPp1hWysildbYO4CsTFopU5zEK6cjO2y/yUqFeekvA0tZNwcb
o1AVANfHObv/I3iITbE1LbamoDVcfbW6MGIZniGiOG/IKTPUgJtLNsMddtCq/tbh
J22w6y00J50PRlClEVvn/4aGEeC3+bsRfxTu9PKRh7mAVasylIuLlXVWWIRa5pXD
btniydCAfT4XzB5ZbRZIvmqHrywGi6oGQjhuQMbCGX0lsI0rcgLe+aHO8kdwrrXg
5s1n4cyapk0h6PWaNeFLeGK+2/owEMpX1LA2qKb5xDcKSUeTDuDFnVMuDz+6xyMq
IqlbfVZbxtWY1ejhrdqOpalw8Hbv0rg/RTJDO9auwgdAcMtY/Bo3UcridKo3+gAQ
xSF9Iyn4jGShhFyMm7Y/PuT3v6YM5uHATt8OU4Y9o1zq6/K0PK/tmIW4mSE8cyaV
qBylqpwLboakwXcq4GNG4IlMixk2oC4JhFn/5L32EY3haq4K3dw9ZPlL/q38QaLo
MuC42NSZUGul4B51Ke06yz22lWu1yhxoyCQ4XLX/U2efr1S33M1yas1IF5/ujKFY
zGFBJh035NkOS6vfXXA122hJ8eOwQEpnYJDeghyYFN9GFsayhLQmhORk83/+d/mg
jm4dcVXKvi04ixyja2DPWOqKmPgIAyRD9BxLIn1+qtTWG/pvNsxFiXBBNNYykE1e
/I5WU+RSuNU+eRAxKfXB1WUJNM3x7RFJIrPffjz4hai+QEWyXp+fUavlgg/Q8vW3
McwzuWa6z2ev5nnpZQVglzdGXArrN8jDQIBa/8IcV5CKWl3AKrO3DI7+cJ8Bx24D
Eobj5YkwqBgXATs33A7yDdx+kXylmPLDWFvnldFwNP3PbVw4f6TUpHau0nU9gDsh
3FS79vaVzc9Qj2prLh1OqnZLqiPKHmtChhwc+1pl+hmX/69T2eo5xWjqPHpbE6Ie
osmxpF3p50YARPOZiM6gZGhjsZvTKtyIcToAW5nLsWfb6cEPfZM5S74hj2XcC21k
+ixAkX1j+CFmThuPFVUNZUMmbnoNBx3/03YwG7IJ5HKc0aDJa4XKysfmEG5Fglzk
THXh7BeRvA0urgFhIP8pY2/rBVKNi+JlYJX/NT0a1U1lvuG3tnH6welRm8fbxqJ+
BYig94aYes4c/uet8Yqs9i1OhKtlWES6+p3YcQv/N1UWwbSqAabVxCh3Dfv8shFj
zPoNwPVTRc8pse32MbUr88aaxYqXNHhi/ayQQf43KpP/kqsYSEkiMPhONwbYsQX6
Wf0n3JrAIre2OtDR4X/iQ+uSbZ7/QydigMJ1tQ7/F0DqFEUfSd3EdpoNmC74YTXx
srG/Oj7Z9m+AFw4k0TSyHoQq+tlIwOjRh58RvfOYPtIlxLBHIp/UQ57YsOQ9KvKG
43XSr3T72tJnXnDf5wUOQ9QHsCMiMrbRi9ATOeq33lJGu3sFKgWXPZAJJEAbPEyP
GkvmDBRFcPr5mrewq7qp9AXQLeGp3nZfFuTIWgejaCTxrh7kApeTxXH+oa/2BRNi
Ik67PYhQw90OyabkjxDx1pyN/qMWJkOAAE6oU4DU64NZngSF/Brbcv9WWKSu2dsh
Ww7UuMTP+LbuCgitDscJUqB5ebdRSwAxaU4ZvM9mcwhHqofi4F1kFJ7AT3gT1ZxE
fRcuDUdfO1blDDK7zd/KXP+AwLhV+5P9zrSK4ox9E8ntFu69FNG8Q9cl7RB37HJJ
Q2HRagKGv8Sf0+ISth/RMIIzp6aL3YWlshaWn9FmlpFpegrMDfILNmZX1A5sz3TZ
ujSSavwF7YuN7sL9kZUx63CnLhTMcLaGF9wUqEJMSkPbhuSxYv914kgDojlXufTr
eUmFCbdCx5MoS60THHjJ5DRSo3MmWl5GNPPlID5HVn9EM77Attu2O85CJC5sRZ0W
p3l4n56Zs9YeyqrOovqDiKBICxlk5jY2YXYHzv1kBvhvtt8iVGegwPjZLx9j1/nn
UibcrXZhwXStT9deYM0+0noKlxQsnVEY9LrslmreNfYjEqId5i1Te8DNBbJgn733
P2+rjxROSEJIVg96dzUOoeBgRxs8e2z63GSAdueiJp82BJ22jwxojESUw4pCM5Lv
yfgGy1XVgwbeCtGcc/cz0xSxyl8KafmpTMbdBUHAf9DsaRA1J3mJgTfADfGowPQX
0XG29kkRNcxwcnBrV2vZj90MO+K23lmftcyDGnMZZ7O78BIug0etHJZXxIP8BwMB
mXYhFFRf93ry+zO3qmjrTyYSp7BxHUIccP0AIcPGi1C6Y1zAaCS1DQRnmDV3gzcb
ITUZ6vIitpn6DBEB9yZh8bICf4FOOrjJAMF/phbBhjbssIv4pduDBR42VdQH6mIf
pSFwAePnq8AwrzWbq5ptVYNYYyVYCphSs2Epgog1LOp+szjaJQNZCNbDEmgKKeKf
9m+lmUM2ahlFErSDpMnHg13R5xbcHgTzYzUZBbEO9hujJvInD5oyRlMP8pZb2XnD
sSatz4/gS/RuDDpsMXv1W/jZkuk4xR9N+TsfSle27vC1lguaSuago/uLazEN7bxj
GRiTy6dtRzASJ5pdMqNl25kNk0rDg6o0BbIMnIXy2sksozTcupfQzl8DLrEjAw13
8I0qyNhYx8l7ntne7pCFxYmyOZklaAhdN4uVQFGNpqHL9zeP5Ke4hlWPqvLbrosN
Yp+5/jxbTGCBEoL2+I/hqivXh7O5cLr377b817EVdKGAtt5tf5a1Bn7uMiTuvZ7o
bx1p/yLxYaRsvakiZqGEMZpIyBoJUHcPB5wmIBCe3T+HW1NXDNjMosvB983qan4S
9c+z1XgU65l23Hr76nGWLE7i0eKWBpr52V6cMmdS3/0AtZUStcdUhy/jks9K5Dx9
EwszzvPsLU1KyQylV7faixkbARv1QL9k69YUDzdlb5ERAwkY6FHqxtCBw2JjuZZj
2prqxmODSGoy6xfx5ocSGknFBIWACB9tAMn4DSoA/J+sneKksAAVOXcs582hWY/4
JEtsIOVPC2cXmVFREkcH5HKdXatJD+MnSDp0HIuTscYUEPJbXqkHgj7tlkZB71/p
EWpNgNTwKifZe8MaJxS3qDftlmRJjf4NJND9EClOqJW5IObiPzWflaO3VgyYoxrK
hHajRvdBh9QyFfw+e5ZmYYGY6W/T8bz/Z2eVVEB9OBf5UnGCowm6VcJsfFeARgS1
On+7Zthp1FKaXtyd6fGin6IDNqd++bLfsX4GjMvyV5trDIvUC2U0avAbiPPGqtJC
DZvMJauziCImHmj92E9aumVUMZ02cDrexZpAw/vWU+iV4Gt58OmcJwby8+vUPTPJ
GGNU92HgLg6bwPdQE4u8VAzJ7cVM2LT++e7NEBn0/ehuq5SBTnIuAi53NVY6hdPJ
XbDsLjkwqIZrbbon0ZV+pJN196X/NRQHDDQObnLtCihSa1xBCfnfXUTFMxJ06jQ8
ElnJB8tWyjhKat2DV42te+39Nt1qQIq5mzY6VhkOyP5o5EMg/PwoHZgNwYNkbnMG
NDdlpruNFbVHBuXUzKLJtegF+W3EJgASNppeX5eElkByPmzvAguew98dUTalr4Xs
UjtjqxwDlgxuw2a/bSTjIHoPeT7E8/4ZiFryKK5GNrosIBeH47fts5faACb1zE7B
x6lC/ClXk3GVgLa59MhRsvtNy6GoTbm96d+jHsK8ouofBK1EHgm9e3HGSttSmiSn
h362Cb+L92dQhot8cjCOcyeC/cykIBZR/i5yfsUj2XgRHc3mQpU7RCzi2vh6oCud
qYy/YYf+AQT9BTAynu40yUN/ttxIEBmtZSLkpyk/KVZC3HPdGMYH2q3FgqtXaGtL
+RRNOCg6A1v6DyBm+60xFvI9yiDrHOi9PfbDRz5DNJ4ipsp+PVOXbWgleUz9DLrN
U5BBLxv6n0U/3Y7w7u+42LzA+xpPxfNugGCSeEuRizZczGwppP0O3WjTxnAJ9wMI
iRgxHKzT3g1A5dU1v3ElaUxyDOPqgAU0Gm1TrZg11Q+Kteamm+j5bxc8qhUOn18g
sYtPixuGjl1Xj+3yRaK1g4Ndq/+I0pvS93QztI0uCJlGZdTwScYII8EspZhLui3x
FDPWz4NQjjJZDV3eAbSldAlfZsnWfeAHNINzAMAy2x4zRpEfAwzVxSnFqTYCv2WV
TnXztTn8McTbz/s+Ht7jjwwOFyKQuFvnRJcvAu+qgwGKzILnlpjvnbdNbEZLhkoB
ViRlMhglgQZuMdzkxBH06ku8KzzgdCZBGaC9iOW+tZYQ3hPuolP90OEUSpaAqHni
FmQxkoZCP23Uw4DfwWs/tumoPgUmeSgih8y54ucHtm9Q5yKicFfTp8NtPA+hWMvB
pYT7p+U5mINW8PBilyx/KTIU4lnvBMJBzPPvRoWuYWTWWwexWq9UqiNd5kiEVZOu
MhRco/XXtbhUKZUJu3Vy6mdLuoWMFwId8WbVQbUFzIVk0MLWMSxdaBbi/0vPDQwR
qme/7IrCvVnsf0DZQW/IViaZAo+yJq8mqX9wzdy9X7vkXciGnEGxzOBQ4/QfvwwA
s3WaePHfofQjSDeVQzlZYf06U69tAkVN5hJGBevyEacGKR3tDL8Wzso7+s3j3mip
b1p6SrHit9hiipPiCXjeN/c+O/fJrKkDeUhMqkBxzfipFUpCuaR0EiG9FOUSFbjD
IdYqxIl8G7Nb9XEVxSbp3b8o0WsVmDNQpCUxj0avSHBb1yp0d9j3Fvsd5QMOre2f
Nz5aNPrpYsS7ioSZBhCDfncyrFCyLeFTVek/H7ERU/SglgI2QXLJL/63st92d3SS
6IGcclsik77/SL5EEFZPhEGFA9KuqkOfIbMWdRC7iZOMiH6Hp763mAyv78PGZrsh
no2moWCr8g3/34Lf4swmnz6p2go6YrWqFa4ZvdGdSdfXAAn37aEA0ie6aJF5Y2Iu
YYzifs6ymSKxn4fVMTK1Y/a7BPurTkTUN66WViFxoeAYXP7sW/R9f0ZSPBTq8U5K
sXJbCK9cPnwTeKi7BDeZXADMWYQAkuMWHSrN3/exyGcMEsZBE408U0rMrHhAelmq
ftyHRYCzJZcax4KuvIEZAua66iMNO5er3PPIunKlWystEJs2myrpeXPF81PvOa/l
TppczbLeuu32E/fQ+utg9U06bTdorP94vquCrXkIRu61+gyz3ZocCpexcOactfjl
4OTwJNcGiH9UC9jzOTI9YDpadyljB1qq5Lbn0KgEc0TOeD+VTh6rdbhQA5syNc6A
c2jgnrPeu9KAqBQbPddRgtu1jX0OD1Db0fuxTrUlWiwHRy3xBjrHRfG2MjtiVqVV
+T31lFhlAy+QXyOq8Q7xx1rCBQUADF7tvH4LWysTRv/JkJfwP4L63mPrMUIS8gYK
Dpzk1dXmdSxj9vJ+azYcx0Cy2iL+EwbWDMZwMMUYyImJrv7UGiPAY4PkQ//3S3Zm
7cMNWfV7XBubX64tGg0XGriyjTArWyMeCoXVMP3XpoVxVvFN4PqD79cXym83bGqw
BMmQ0IhdhbRMxvj1o62jagQvTuN1NkN/aEJoqFSKRaRgzVIqt/v8shqJ4uI6GZWt
NSR/+1jtDAZcCp58MW+Ybb5ls1qkH+kFFtM9oRGarccUybozKJw97yoIwJlqTIIq
kiXwjPvCQcCum9RwK21K95WS/e8wWc/KZe/idK6u+qQUvBNquNBzi/+ou69JYoly
FjEEIakz3ekKjkgxy13F23xWXHYTgPqz657d944hCjcwlphW+Ex1TMT8YRqjGRnI
cPehzp80k6DoKW6ocvCR+6ZT4cnVae+G1IIL36g+HNBmoeku0ZCeomsl9IEmchH/
dNsBTy9yLM+441JBs0er7W6bK69qK/9YnaZTroyhRfqFj39r8S9OgHqgxuuHAZxy
fHbNPGKVYRrTjyNTZK1Cmv48TyVBC0ZCOkqOvUgVfbvx6jb2gO+kWknYHeW9yCQ1
tPiRvkfTLdxXVJm+XoI9VyBXMGFEdcOWKx/2dsHHQOPwWPV6oRqD/2OGNtLQ3Bve
v5dnJurM6kxGZtjSQQ0PGsiiDi/VfQ1Di0C2Uj+8GpUcrX3Eo6VcTmaEsuUhmQw4
9Er9qfXtV0n7Y7FTSZKpf9Jdxl5wyld4CrmSNPl7ZZqOdSCZQDeGkTKjDgAM0C32
poPpzfTOX5hkw1Tg/6e3wHNKNjybHnqNCgOV3jk8Sjs2aFMHe9XMtugcYBHutM+c
fpOh/wFW59NM1ctemUS1FotAgAcSlIlYqAoNdJ2bZ5Hi5NyBO+fm05wEuDhL35t8
UuHCrMmnCocayefpG8ml8TjOKc43yHsO7dUOLpDaG3+hiDNoMixRctiYsPMJzcEN
cdXaAfn11mBVw9czIbPNdnISvGNf/f3SBf17R06JeP9xvY5n2uHFZkaGbfi9pihD
dmsbIZGSIZ15IxYZauHp+cCaCIwOiWl+TN8TrP2A+GBaW7tBWS9e+HDrGMh2zX4b
YI2Ij0bMq2RCDR6rXAgvZq+RubhCmgCNfXzc3pRuRNM0ExMraAalFvwpJSmpfiQt
ys+/6eSYsHTtzaMLUsFlJYa7ifL1fc61RapXFU/KFy+kMpLbSrmw44rssFWljhm5
IytLTDcSwZULt23PD4oSIzkuWe0VYG30jBNuerJYLWu1GPrbnBi0F4OOLc22Eoxa
K3s5G2lthKnIE5vzSlrmfgzNwAJqGxP1VnjI29PIdWbu4byiu3Mfea2TWkCRkuG5
1UMQA/mdK3afcjde9AeHZIyWAJsu/HCNtO9TYTl98hmNWFWezA2X4VvyyuxAz581
KNpM2D3rha7wnp0jdD9pbY8IU4K/gBPAbT3UaKdWaAlHnPXaRr6elCQyBuAVPmgF
G3sXSAmuYyo468JS54NIkUqkU350S7JNfbqUcIqm8QxGvVDqVl/IA8jwzb3fkG7I
noRQ9biEPOFek78sLdRj0sq0xDkFzac5wmUajFtJYXsPbpbKo1NyhkJnmNvL0aSd
gv0kOeBpH1CGsVDBGwlay6WwmNfH4KvrQUiM/1lzQnCIM1Htcpt+F/lJ61IdsQPo
BS2iMFLKHwJ20pe8dOD7rl90O/vzD8eErArOV5nH02BycV57Gw/KoOXM+CFT6Ovg
2MQ8T/bAmRfXzfSTmFu3/24JiHsFoCFfzcolLTDn1hq3Ba30RG3/mXeUTnfc6rTU
hvdMWKnVUPJQIRkycOoig8d1/01b1B7tA7J6jm8UjEeYEti8gPfrIh2gcdRMLMhT
n93zxvH9EsUSqECJUIKkoqMAixIGVSnhOO/tdfVGmciJRna0PbcDKjT6zfsM2GFW
O2hT0yrG+pVhfAGekOnG9PpsXZuTVkjDWcWwTxgtMr6lshvOpiZObbsvq7+sf11s
ESh5MSHXd5Bvz4pav3iR8RnoIpVXgJwEmqY3geYjPRr60UDKHLJjbhnJ179VXSny
8WkahG0IuxU13jFtx2UUYq4el9f3mgfJcy8LGLWX2qgq6As6mo+Fm7d86vEeNBik
/HeAcF4behqKkcPXGdbx/rBjjXM8Bs551LYQWJPN7Zzyt1BuqrfNYlan2K+ghStm
aRLnHK5Dz2TnDQQomd2Qws6WNg4FD9Df52NKza8yCD319VcbobFNuEdGXj96L0Ln
y0Xv3II/qzlocamoRi9SXloF6wHnwIZek/hqksaqQQlTx8x4Zis3xyxZ9yz+66HX
m4P6E/I6mplNtvMzM9LWsndBfxcMT/ny+Jq/DqThErVy0GcWRuqmKPiYJNySwbmA
hmYt97pkeH4ltVhuNja824/BhzUWnnwm0M5RDPjh8WvMEq1csoTRWqdt+PiYy3Gg
9ej3QKfsmXZvAW4satfs4QVEXeUGM/d0LeliPs8x8utLq8ilbNPM09AVNtOOkS5X
zozHZIjv7UNWHr1pU3m5I/Bw+5haxC9c+8PfBbKrkUy+Lji2i/FFeMHsTM2UsA08
DyAaFRJx84RA/iA7EyCjNaQdrlrOsHkgp857hNVkP+F6JDwfh3RDOQ+lp+eaX5X4
gBNb0FIxc8+MJqyRiMFUhJ/bzvY6tcm1FbHM7wUbovzzBitFETvNBfmBnEa8l6Jq
iYRuqyiwGTw403KY/vxoU6+PEZuRXOxrzTUtXAYhzjVAyzmgTTocqKTxub7ZCsxn
Of4p4ANCpxJmKay9bwXQAJ+quBmVwmCQ5Rj+9NAK1zuB5XxGCabcLjliV1Mq/wUV
1540riLZIXMkC2IPmqJJxceCBPHn1zaNrTvbl6vetTpJ1cwCNWpSpjfd7JMmDUbH
oBqcNoylCZU0uf/zR1e+1C7kYR8ngtWaTw+RxhhnFzayvI97P9CCfiXFiNiN7TFs
zjuXDTmIJRlpssovCfxi+UvhANSgsjR5JUftlPLYIURx90H3yk04ziwGuLrE91ev
9+fm+U13qErSb9VZ4ge6MVI8IXIFViVAnmfnI04raQ7MTPWpqMdaN3LFvPuHyNq0
Rzd7Rpk/v/iT5Y8UYbTQRWcO/8vJUjMCdxHr6GeAAIFIjYPqPNY9VMEKr7TVOSqD
ynNadns7+HdhxraQFEeps1IdzgFLyZFzTPlVKYyeTD2NmtywpmxBWbb2I49ZKG/8
tXuYWBWgWEF60PWvy5ZB1aUcE/7aGWBHEWczyLlJOixf385ZOqP5Z8paQWTl23tf
sLxwh8EFddEE4FolRJADqB3b9BBpuDsrxO8dEpQgv9t1Fk91M7SLTIEKQHazNvoE
amVedN2i0TanX0BFr276Em8rURAbW/o6NdLIo+KEXxkTq+hI46DHwCnavqeNitym
HGPQx8my6cOxH/Fob9QUVaT9v4TiCBy5h11zR5viT5hRSLYIIUlThntalSsJ8aRF
84QTvNrHFUfokyRt8sJkrWXkyMhH4PPycuFkf0XYqnzIEVNq3ar2Pu6KOsdsHexW
y5WWlIwi87865I1Pz+0IsMhDSO2O30x+auUmBq+WO1j6x23+xS/XTBbcOzfi9RiG
Mlfxo5UMLCg0h/vMxmbKBPaV2vFpt92qkRFR+vknlaG7YaASjxnZyG7/gKuhjnEB
G3VICf4zy7y5lDJgTz1uIDAJrjtR49Jhr5UB/sUUqSjDC3Ey9qqrNd/yfIsRQdrm
vXvelZQXeyY4zK/kYCGM5LsI7ZD7QOPRP6NHrizzyuE89/ezwp5TVLC6Vf7yvfav
PM+Ur0ErWdBS2o7qklK2Fy/lLlURzPl1XTHZYrAENO+dKzhWDGR7oun8loR6MqY9
DY91FaivDDse3q4WQUoeWEUpbpYlSdugqlHduwoc7etBi2+Jly7fjSdTfjXPh2gM
Ayljm8cs8LBfvK1odab9Xu3Nbi+LK/PTlxm9tPXMJlgda+Ahzbqa/hcrv4I3jSI8
y0RVi6hmhaVzn4+Ds6aDCB53fGZXC9TabqWWEHyPD9zI8Myf75fs7dvqobK8MSoc
rQ7UKnnfsH0jH1MgQF1b5qsUtuZz8a84Ky0krLN9A3Euw8hnKMEUTG8xr/bTaqu5
A5VTbToybzGhjqAcvj/6lNCNitgHbP0LLWORhARv42tiykWvHaOH8G14JDebO++X
7MVWGn36Zpp9m30TL7Lc3Sm6Yj6Hu7lQx7/ZAWPf8wjaGFaXmBmatxxgj6a2xQZR
Hid+LsFZiHcC41x2eFpZWhvBaUh0X07pZG19sgSKVZCuNEGngW61qPYOw8e6QeVy
jq/r1wmAbyYfChnsICCLTV64BR0KaXavFNLdWB3C11FWWp8hdRwOdSRb6/zmND9B
K9ElKJHohCvxP0x6hb64TpqP0ui3/aP+mOQYGp8X65hYv0tYgBVQUlgu3nWAQSMs
LhEHU6PYoNdnVXITvavA7EZMiikTLWTICP6FKEYzgYRyvFl4QGEre9WAEdhoo7qR
47ZEihUcOCpbmEzBOrvFIV8FFDA6g2NsE1GRZe/d/nxVv0NPAPua3Fu89tksfWzT
YEpf2HPTqwjLa43bG/mq6pEUQaax2KqdBtvTG12Ml+WlT2ytnn0yr9TedkJTEWxT
ZdvHKrLecefVVlWzzq17NWOdkx6jXFUlvtljNsZxKFf33+DHpxDCVMxC2E/DbC8J
LQkANkQGkzctAfiNgV9egorLNu+o2JFDErQToIJ38im3FtgCaS75hQdhg4T+W8dc
yvHXcuqhZxfcDu+OzcG7Fn3P0U13irQ3+h8f6fKG2QawvVX6rO120DfTk2BRMtrD
qofxfKXF2WccoCB+y5yq2m1V8OP3V5LaQkct/S2C1djfY40uO5ztgPNV66435dxU
Ecf4Ri6TxAW3cxFBq/+FwQkp/5M1CBHIlN6HTOUPfNMCTXd+oa1ecVoMUPJOPmis
APMxearcw8P1R/L9F8EvcXahVUEGJz//98q6/ksQmabfCz5AM5g+0Nuti4DyEyOr
FoNHS2sWhV2Ki+9glG64yRhUAk6kGMpiECm4kV3c6GgfUzXo/a0AiUKK9Rm3Cpbp
g9m4OP082zFTYbBMahvQAbwgcVvM4JF/lqBxUqun/47264tnIJqZqCqcVkHjmIAm
GR1p+XALX/OHo/7JE9TRWZk1egEshnFae/zknX5F5gSV3SHAIZeZXu0rfLP3CS0K
Lgfmw23hwwZkqvcUI+nqj0UaGwrKoOeRwjz9y+9DAp7H0AqAbODE5Z2zj5f8NvSj
NZ1bVN4GLaVH10U6oqZdG/kABXwWR+wX92tE/McOsbk0pF7zfxeR6XV+UQiLN/Er
iLWnAMWT5LsJLzOU4GkxP/s3o7h0P22JobJ6O+1T2JzRO/325NbQrMwziaoIV1FA
FGzSSSzv/dniL2nXP7BHe1vqOwGcFWfpNcYN/muNOgd2WYV61DTE9JVBQOnQio/z
pm3aWFUYdDmnuRDaFSj47dtbObIgPJpn7vxZRVLSVo695RtviAb+Y692McWwvvKX
gvsqIHr7+HHUjFI9N3f/EYqZlXswiN85XOCaYH2G63vIOTUPXIxEOLc42giiPw9L
lEOXR8CEloJc8pOPDT2jHJAq+ickzKVYw0fQHqrv5lfksn1v2CctB5GPzRtH7Gvq
NKR7zrsWxGTqGTHa+/uV6mknSOkspw3NOM5WQM+raWr8r5md1HqZt8VQlZve97+8
vxh+oVKTXzJRak1UFNP0guCnPDSYPDll7xdyGmU0jXnbuXYKIYSC/bykRwQ8wr0O
3MHLYL/Wfagap216vVQ6uhcVgsVrchTf51Pd5hdwRhBSNqq4W4640Z1aaRAnCUTB
BhHNOVnhtMR6L/ktl1n9UgP1nK7/tAz3ySvUcwhYXlejaDY4Xr2VgLQB1Vdm5yHt
GlORU+R8oWd24rrwfjLkd1x0jIZHZjmMRm2hQG/i0RPhWak00Ty0GmEpasS1UumP
ZKVB1k0V9qIOWYJHu4oFxc1XSLXPdw7Khd67s8xZFgNnhahLr7Ss/pPMcH4BFsB7
t5k7/b9dJ5agaeF2ra00DTLFNWIuUx+p7WH2Lx+toREpuQ3fNSLKQZnN24IENEpl
KZ0shSstdDMRZNGej2hT16QJihrLYmjqgTFBlKmMbg1FiPRBwf0urz9J8XEvyEhA
Xh1XbvWqtblVntg+1mCSoN5XWwMVTwBC7HJMo467nw8mta6g1ngbV4Pu62P4M8ew
hNrtwDlAMAjFAoR44yyadDhZpi2EoDPOqNyB3l5ZLU5AbzTGTEN0kQFuecjwfxsV
vLMuX/K+TzgT6YmqZdOFZToEXpkjAP5HZZMr9teaqOvPqpYIe9rdjrWapRklW+8m
qfN/l755pX/rhMcaN4xkwksY+DijdF6QNlWNADwM6xiJryFql6Qcd5aWnYu6X+C9
i7flS4/PegmCr7zMGLJjYj12KR4RLcsb9OlbPwhm+lFjm2NDWoXU23G/sAKYFrdX
qJs4+SUChUgBFx/5rCzNhJ8/VjB/OS7G4J/A1gz4q/QufojbTC8CweoTQteWGEwy
q2lj5akZPdCSAPqmXutOsE0TyAaLFe8NI5NaeUJoEVOBXr+4LU7+XJGewQjHhfS+
f+2gn45u/No8OaG0gHiPwQ+mBWPlXaa3OdrjT3uyzgxjP6yD2EdmF2tnE1TMxVnj
pxdjPQgl8EXZ3GqXCoYdnYxWahM+GJvsol0OHA+0Wbp9qQN0p8etqZve0kQmYeOq
zSgXvJjD3p/LVU95LmBQVIacf7xiHQ8oue/W4jejLTe1rXcr5XU27lyVJHjE5vSs
o39TmQ2/ikIw0TehuPcEjLdzlaXgkceE/eVP+eohfp36jLpkAB+jC+Qzd/N5pDY3
djsrdo29TZNjp//F/sp2cD3zvqTjF9g8DjeYGuRXvCxiHXi6CzEYPHuKLM8A+E6R
WFi43qNMooTsElCH+VRq23dsGHSIDmvFmLNMiptToHLRyZ5XT2b7zuHqkoL7SG/B
8HEq55LLGlO2f+R9Z94xqTuY1X1T5apsRX3i6dFjdL6SSn+BiCllMxQaLHXggfHW
kPKVGsAWptljKYjYCLMTMWb4ynLAVL6Xe73uBKyWowX0iP5ALNrI0moIgixFqwf4
AAqzb7bmvXjG3lESz58QTR8ftiJnsXaZqthM2E/nVS3G9HICU8/Xq6ktyqjVIz+S
3NTG5K2bC3LCAK8Ve/TzIKL7nKw7KbmS3Y1vJR0uJ0UTciibt+fu6Fb5Z3CI8Hcv
qTc7HMio7RDAnXPBewZGFvbABAj7/61HTopmetavMVqpU2vxn1nVsqBnElJWojNf
EZ6zuKFN0uZG+LtKFb1FHNa+hekiEXUvw1OXbHr5mZujFH53p64IUBMb8cT6+kiH
UMl8B+0+Q1jvIXVyDHXjOVu4d40YSRWUsI7dC3rwXJT74fhUnqkPWz75qkVDWYK4
WpkW2eURLDllrFB5V11eZzpAOWGEhSLEQfmFxWG0EsC851yXJZss8aUfkOqEnLKB
ggc4o69zIjMNYClQiJMdZb3N5KORst3AL/elNlrp3DEkHmtklZVZegAj+ykRfeun
CxUMhXFJUjzUTd/np2fAFiFY5t6WAdaWapQ776wHXKWOMWDgyUm7rwYe217NNr3q
XQLaWJama2Oqy5v/4l6Vm+FeSCNAQ5tSZM3QbP/HKlS1ZbUQQoLldhDWUkiQXk7J
e0nNZupC32s1x2Jq4jYwjNbEkrW0AcMr9GH7eIDN+EGWbuSTrYg/hLRoYZVQevBU
sLJMJi2PZYrldwj7avFG0hZ2ZvOngxBuCZabUvUwlbgumxiMrvbTOVVTruZWsthz
bEAbQJ4TjP85Fm4VBVsgGqqEDBSWbWZ0WL4wyIxcK4TAVIO+kYDVuYDBdyhWsMBp
AW0QhatXVZw0p2XEZo7SQ9XUy8IAxQqTSmrUOFwzzpNXTDrCUOVThWAyYc+APq5z
MSOM6HHoDDv7Jgg0wWEcOY8N7xCX82mYkHc5Ptc0+3Q2Qh6tWjx0HAjCblIoXBAZ
NGAgT0Squw+xmXWdAPR1OFlLRoUV36uRXfq6Co2FlQalNeDkIxRjbVjQuiv78GA3
aIyD/rEVObwPUBE5aH4C9PTQHs02zVUTrD/ynph4T2d7htQ9Yzr40GFYvjxZEE9C
BXSGLUkhlHcFmbj+MvgI582mmMn6mtkBV/IQVCQW7HQwfMDyIWmRGVBQXnYEKNxP
UNYAkrjTaTU8PwDp8a4ovKTBUy4jdlWBbz2PlVoqqmhxkspe4q/7oT+7EMlQNKMQ
3woLXq3sfDhVQr1T3dtJurZ+hXFgidcKodeiBsrM5vbfLlJG6YpspAh0Vb89QH7q
e/HBpSrWLGSoH1QlZTdOw/ppfXZJDvgX2UWy/YoiJLHxQmhZF0f17aHb8urzQyOK
+t/KLHTTa/J9kXoQuJkBBM8x8q9M/aR0JGGTeqff7r77Ok6TG6xx1CVgzh8W77/O
VRRy7MD2v4kKD6dcwjZK86IzPGneMXdw2KEVtMVsaTyHjLibdHbaYET+EVLktDBa
JqYrlOkicvo9slsp6oprSrDDeuHrgZUkOHy6ltdzfe4eLBkz+qVo7XLDKDSyrIml
nU23FSjfAuuUzI2ye5RusVBWiu1p4LSzxUbFPQRzx9qaG7D43QQIuOh8vjk2l8FS
Fgd1Xjr6vH8Hnb6UFF/sisz6VGrr7T3KbHLskkj6CurPNBIBEMJyWuGDyleb9vRE
kciBjg99H5O8o1A66c3XSft1440ORot00+O+s/JGCvM/dXzQ20erNB036m312SXN
TPGL3SrJhV2y+MXxjoO6/HOR+CmiL6udyPt0lbwm1d9RmF9DREPb26K2dWAtDY8Y
UQpVPjbqEZvfy+/Dt2WxupgvyZh9hPP0w/FbEybEo9K2aBUZqLA06JTesSzNMyBy
wsLAL0KGlU7ncqBU64iFoC79Rj06ddSj99QzBN3jFBUe4NCHQswLUWQHVg65UQy7
N89Z265M2bfEAO7Og00eP/+tpvusvQiZ3Q43C5xhtDhWWya838BlQaejVW90zu2T
DaZzCorBzb2mWs5Zht9QhdIXYfHjx56nqTLdCZP0PbYR34h/81XIiRdFaWs4Rh+G
PZAjmyywM5kc6N2qi9QAAe1SQrcYpfqM9+ezNrc9sKS9OEsaqW9FC7Q298/vi5Ph
imuVmr8M0P5iihejM/v9ULDT6XbqeOTqbK5z6ZYnsypSRZtCuGyIRAUcNwHOPmU1
2YDmBdGPdDu62qEogk3FDMyIQFxWi3yJI6kj3p+7uBG3MrNktWcWko8E/soe8Npb
2ECXbUos1m1y0mreL3KTZw9N9s5Bml0yIr4l79TseXBIH3ipklHCIbTP6bHDsUDt
vN4fMyXwOj5LO/tuHeqmCT/3+CfCtPABeClSm/UAAQHALPhFfiHiHOvMzYWfcCm2
JE1oGc/YKH/igHcgxvzngCHcaD4VUQ3vS7vTBhK1GwnuZtXLd63IbnJV3C/7/615
qkdSHGRFp6aaw8O4SGs81BDSzp4dm+AYPlOSISXIHw2PSXUHz/mvZx1fDB5yiEM6
1bzAJLU+uzWjafISCV0+wrm/XMupq5IgQEmdRwWlPx6g4DQ6IFVRUzhaR87mAntY
jI+UWtCCfnxQK/NzWRCHRZK4M3fmqws7D2N8VZQFJi9Ba2fXFtJ+AX5zzZtOYV5y
UuJT9uMf0GfpNfJoItcaxz47+6usHhgDqtLXvJ1gZD45a92UyCZEJ2IWTjHfuB96
ibuCnT0P5Z98qlkXJlvnEmQLmMnujiefkeKesUwKfPNIZAJEF1ha6jwEwlGoy9SA
lrmcqThn+ekqcf/25XsyuiS9GtlEWyaiEbuk/WXc0TIGGSJ1vQFf+JeYAQGz+3ps
6G4BSKF9sfhSi7zzO2cV7GyiiUoiIE1LVQUeQC5A1rhrF+D2Lxsm2FGVYKLTjwU1
+euxkL7LlXNAFWGxTcyVrsE+j/CB10mN58rzabgrt4oojEsD2oAbh1oc9shhKPJc
89upWDp0p4iF4jsXDBozfCpzm95wnEtFY1XpuGcuEU6mvu0Jr31H8Bni1XpLnC/p
l6/KqvjeDpl8Znbk9p+l8rOTBmyB+fcvZqe9Rlb42gT3r33fYa87DIN1TtsHM2+F
Z2I1fEl/floxkn4O1Mvc0Ymw3B2se/kZXR9S8Wxc1puHpZFoBrafJly44++YKu4S
v2PLpVc4NcmYrBEN+RK75G6qxsgw0qh0DYKHa8ZfrTW9wfSxL7iEAuuAJrqZtQaM
ZaJN3tfSFqzt9AJ7a5bLekZ7Gywxt+H07NDojlRQ4xr1VEEW7n+RDEnr+FS2Y2eD
QqlE/3SFmXx5gzz4UyH75AUnR4Jwpux4Di58NGahw5+HJ67o6uqyqxBBFxK1VCc8
eZxQXP8su5N1iE/G9MKxfRcrEByigbj3KoRGVrQ4uT9GT6a7nP63LtqpQqfGiXSK
SuAktZOkghsG5oTA//cg/knpx7PrgbYKWImeJowM7rImzQ03NcnA/hhFJESH7PqE
uGK3+nYoJGtK9BS82/YgEDFdj57hOR0r5/z1duNw0tS8ccpgZedxuDfjOPC+qJ1Q
26sz/lGR193sVtJ4jHPUG1cjMJC0U5+xelCtHk2+MKn7HIkisYhJrsJAqvOV0Zra
TDTUgZaTgc4S+owtVOT5+XGK00rWI/0KkGmIWlt93u6a125WzbxLWUsrigeUAcGj
aloRoFEuKH4+xt8V/JJeS0JpG3bU2v2nKfOS/1sfyvWYE2DduwtyJKZBC14OkZZj
u8jxt6bPFahbcZv/zeKyCUOZs6gappeaavQdb7d1V5TJzqtErJa1flhgRXfa21C8
YOxPDJUrbiYTanlk7lQ4sDE53X70KvhloFXjZ2KYdjsGDt1wlJzAt8jTrfdDwyaL
MBVaJmVcxWa4oV6y7GSlIJX/oRzo8Zlyv/RmszljUb4i2dcvI7yTev/lc2jRKG7Y
xr+g3e/7Jmqi1d60ZEe7Z4bv5YGaPObX9uNPrzaUTAYlCqVPyv+zfVUBHG3yGQAM
loI0sl6WYyTp6bAU+0QuTCNTQ37HncLHAlw/uwZHoVcoYBglvfuERxVp68K1tbnW
RVVag8CxJ6jWocM04fWGeCuW6D3AH/zkt0YlxCLEi3kN7twrRfZB/1+KrATLoi91
tl6bv9JFsa2jU/uC2VjT0QfIe2kV5v2WwEs5TOjJY650X/cVuM5i9JKNc5o+aUcz
3nncg97eDwllOarThoNfCwB2sWsoiYlYNQirMrVjElsJByxvd7WC3MMpnwJay13d
ohilI+1ehDeiXJcUI1pxdyezqjv5Np+pbltp/CkVCTyoayU1QQ3ZkFJYlOmbNkHV
wyBlS1+qzT21zZ77WoSHAtbCsMYpe7c9WyB+o4dGJIyyDk5WS9GTtdhNxYRqsTIo
zqpoc833Vfgs05HscaUWOyqyGmCfOs1QJeTimKxa+tncWfjI4XHyRyuyZ+7gQQrn
i5TRVjTuOLtkXsbknEXLWmQL+IQfuTjntcDhxOx7Cnt1Ubt0Vqeu0TOMgplj51Io
OdrFoWXz/suH+ZYn6kYTOt3z7QZe205JI90XyGXqB/haD3aiw1yqXoDJwM6FV0s4
zHoY3IG5zMVAiheR618T2rOvvTIRL9BIxSeKnLGgKjw8QcjAhEpmxD+fJKOEU27x
rhiT3lMD6c7Nc3Z1Vx0GWdy3pvdnuAGrW4byWo30OXFfnPCoN+jLTWRknSQG7HAH
HK2UxwP0Chi/zaD76vByR0kolyuo2uHQnQpsN9mStSrm+Fb/58qQ2KsdTUGrrRHq
0pp2aZ08VPh4bGr91urLERlLbO9vyCQuPn7P19MbJElpEC/uMUFfimGSyKmIbSQn
Bb8SxPc1A2lDgJrwzcRl6QWTGR8hX2MKZVHy7MVIVnXaYO6XA2YcmSb5yByWR8Vl
nF2k/vSiz6NX5b5+oQFU7kKZmlOjPmYVPF/c5V/tLnmlmNpM5A8gz9aE5Gvuj4XZ
9LFMzh+Wg4h5h+2LdKr27+5z19o+8H9DK+xwlM9CWQQxeZSn82yxyDqtVj1ckUP2
YiwFGBGRPIkx5PsNhDVWMLeHjySHixIS3p/mfppuAaLPz4Cr2iJAH2bi/nkon7yz
ClTvSWlh3l6IqkA9en74Uhr7adpTTKywRQnUX4YwTqwv5NulnAtAPaDIn1lrSG3t
vYWS0xmiIiNQOFtuVICo2/u9A1KU+PVNR5hqWT6jRx4XRmIwyjOEexCGLLVjdQ7x
wVFxn5TT6I2IA5XeBFYdK/fKBWkhGPm3mdpfDfBQ8gcqcSkIJEtR8AF35Aoa50FN
35bTBO2W+fVPvyIlf1k39KRoG+y5pWkoZkXxl/2Uv0w1hHycvYIfOeNPlw76K8To
nnT3itU1aY8RIq9xcvuSdEJBCD3mF8S0BxrkgHoH38zqhnM5YOfzM/cegeMoEnQT
as2cVT4zY1M5tEd5vo+OvnG3qKQKc7zG8OnPbE7ug02JT0eO2kw4v+OmUqJ/Rgrm
ETYqKNanVl5JGm4OJ9lcbkaXM7uy8vANYrkasHh7DlB8cDJ+iIPTNCqSq9VIhFDx
deRcJT558hf+ZaaKRHeILVmdqxZlhoyBU4VLPRsU91dFsbyiE9D2VW5pmseaY3JJ
P48mudvLO4R4YR/Rot2yItkifCLrpIURdJDwfSHcBQiH/EAK4H+At+tKjXOWHy+S
y5JB3eMilK7PlEvX2Mf0ze7N/FFXE2qWDw8NNMqjLjVckI4w1363xaz3SoVVDks6
1CnbOtfSSJHV+XkMLVcDAXg3GWgkPLhx/vTicU2CcCVN9CJFK4I9SmK9ms0FgN/V
PV78b3p29plDHRgvSsUKFqjeohoJttbGcvxAVVWd7w5AOcdsB/+8fyQNLfSellDr
oRzbWE5qf9ODFf2cXGznEKSs1ZP0QeyiENN8dKHJ1ZR5fx1N65cPCZzzmbmU53K/
637gU9K7HCKN/RRLKyd/ItHLfeKsi8a8ryglttUZIBiTQhwh3h6pZ5kPeoqyqQjt
jR3gErALubKI1wTolotY5s7A4WepFO48aavGttJBlqaUd6msCB3IWijrt1b+VwEr
yrFA03sWLw3PL235lDW3NyK04n6NZ4scGQrjh8XT3fJPVUdBwH0XARuI+HSysj/L
OQR66754b5VHlaOxwIr/+aPdI4CLE8um2CUqr10CgygXFKvcV6DKCqXhZK34zXvK
AiIJJUkgn/VnMTesqFczfQpadYhbKtYyQKTatXJuz824hiRGnEfRl11+jMPmz0R8
FY0C5YzOnDFZdEZONLvAuXExtwPDapAgn6ReQJT5/Hp66RgVNG7FKR8DasD6Awy2
t3hvgj3wWAp0y8isBeBtDm1Tk4w9N85O6O8IdBBKNiPl7iveN/i2KhaM1jjfBhnx
l3mbUBV9ACTzsr7AK3hxlg83Xio8BBRNkxxhDvAEGSeN9LtDUn14mpCg4Hr2SRyE
babl4ZG8DCcJKVF88HWGA02riToGvfC7r+OISnak2XMEYKEv1SsJIcQdxX9n+5BC
J78kynIUfp9ZDSuIE++HL62E1YKSnxW02jRy7jE3bgp5qoNFeGpqqPQ0m3aND7RB
ZwmE0ekyxCUB2UcmioRpBm425RacDEDLir0cU0loUS6i8aiilS1v2VETC1vBr0Nt
JzRbOpp/D/bCA5x6VExUtbDTg8RyxA9VAMH2S1K2z0QdLGQvUSYxZO5AL2nkL6C/
N5J0fPj+KOvf8xEeuLVgAVLJoyon0UbCXaAokuyLZkThSHkGYgZWDCRewbzYQG01
xJZyEGRdu8CaGqav3PCH15PSIX8kd2Tqd1DjStPDMctF2b+7cl8rl1XeDUfQec9m
OOvsz1jlR0gKhcoKyIAEv55eJzw3MLFtTHK8hlSwpZTyOd/n/ms09ODGThzsZoLb
Dtw3/rl8Hijnfvfn4HkOqssxCIYcDiGWceETFtjUvDPv1DC2OpSPITJfpMLbtBR4
38+RwSfqoRQe1SR8i0W1VKdMbt/Ehel4MDBbp6E1vPyTKlsIymnvxpEftT8SAsLS
EiN9iMtVx+rezbWMn0bL3yenTPEBRyRFwHW01caM33ZwvY8XW96WLwT8/jefpgP3
+KaYlO7x+WOA41gVANR14jfxbt83/oFWycKsoapBD5Y7Gz3KSOGQi5oO6WaKBVkq
cZj3g1DCY+bCb1phRF6SzIO/3OHICjUCnmIkUFyu3unoD2PteJ1W9eTSo7xTP4s2
3bOolDjNgfBq6c7AnTii1uX9GA6FWeT+Irco+784DTDrY+lPps5pewSgWjVSOuqP
ozpjw8I+Nf1zKJSC3EMSHBGNWuMn/NNT7+rl1ed7yNqbeV+mTRVa5NIHSLCYnAhH
3WtcdSwlJY+Sbi0c3XPTXQsYnYBB7yql9UHQuHY9ilEJoFim1HQoHJdFwhX2wBfB
RbVHrwnWWS0UbjC2ehRZvX5giPXpwxy2QGzrVvF/WIWY9ueyOtxBHOQUEwA5kh7K
rKlPGaRO5JqHZahg0SUpL1NR62issq/Cr+3b1jeiN0mAQEX0VqAxBiC7UuD55t2N
IDWo23FzK2E/4WivyrKPYT6B0ZApJCSeQCrr+BcgMuOw79UsljRR359NIftc9FE9
MlZZfyY1iR1zC4HLV/irkzZA1uQ0jm24pjrhywnBaBgNTLX0iwK4j02iH43tKin7
p8mmNr32s63UE4gjzwp+KCy4exB7GtXcBZtSpJ02sF2eyPbol1Yx0EAOXAI+Vj5N
WGGZgnPMLViXsf1btdgsdL8ccebAiOC26VjPmjJI3P3HP8ZSt5AcMK32iYoFqKmF
VwtbgF1bEfL6cj1SnBYkn1IgMKrB1paxQw26OxauVFvCdrL8+9Pz/um4XKXOyk6I
tGtzMJLC18ujJxBwVUy2O7YhOJ0RtNbYcqn6yDRq9VMdzhWMAuBVFhmojWcwGbNx
1uCC5apzYQ4c8ZBTs3tffBjhMy6PrSMrAftRU5u0TG6sOGgK59Iu9tYdsiUVcdTl
1D9zLdg5WGFd97u3Rr4yFsgNEwut8dfHGBTd/clzzY7JUoJfdkCu9nSG69vE6qKY
qhdFhjUPgTjdXPH03Y2nAjYto4LOHqD0V3PkqzOlS6aclWAJonuPwRa4d/yIeb4w
Wp0cum/iZvi0mZ0fSbTiYTUpSuNzGWT3d7b8Nyl01aLPS1UqwD/uRDhsrhKj3rGC
igiQAW8UY/l9ZK05aZWlJlOrlLID44Q3MA8hLnEJuDlZ+Yb3+NkLdj7tQdWuvzVN
9A9sDUvRTWpsqh7+aAu6e1b6sIhzgmPH7Wwd/BhqpHgZEvVE6dKFVODh317AMD/y
s4FqtHTX4ydm98XLwjzA1Js/L1eVt6oSrHrBK3gDpYV/IiEVjCy/7OYkHr+jnZMD
L6kgqM0K7x7MhzLbvzfB3SUBTqP3RlIvgXfPOi9qHqZm45iwG7I7oqrFbGuKS/aO
n4UXJKGzwS6IAlcTS8nW2rjLqfEYBfpQ0gD81B8CLqnf00ecxDePt9uVSXMGjuDh
vnUWpsWDFT1kWdAefRwljPFMEzkXEaEEbtbssYFdanuz1ZQxJ+BW7AZ+B5VMsbSK
Js6UuliIK3id0zi4l9Hx4M2fmotcpnNy88wRooA85ya25W3i1xWcUdheTa+iATdR
EdwC1bIyqUh80R1CJfa8IgDqoS4ZrcEAaCJJo8FdjaBjl1j93OniQj5pWfaenCR8
9YEMAWN3vqyvus6EW/6UazGkCzrYhhZ2pqjD85ltpDb1PMAPwYgcim3fzSqWZGaX
4TrR01dJUwAmgqmbDrj09eN5TOnu/y5oZ1204AiQ+UbeIjd6E3SYjtJ1sXB6JkeT
CxMcJo+nynx9Y3Q9bHQNB23uTSRvp86x71V/8fbj5/MCVX5gD3YaxYR3jK6XDPxK
Y0X4L1koVrDllDOphAcF/KfpjeW0gbrDRUZLxksovTMxU/8LmTRi+SgPr0AMtATn
mCaB3NX3TFYT/RF0vZ6rEvw/8JILCqNcDDPykK5z00bTH7xuSrDtbF3XbMufVGz5
qdph57Wtv/gtAeOCg5Z3xNCIS2CIFlEQCSZfHvzlVZ1bmSUzgLzFLYRZOwh/UNkb
bj4m1tZUZY0YjxqsW77hkddtrVlROBCzvv1JvOzbcQUvi1XfIHdvJ1hMWreykncG
YKvpE2UBDdJTOitamB2aaXPTJp3FRhp2cw3kvS5EPHbWsl9oX9wyY8Wvs5KMmUv9
sYWO+yOYuK2sx4W5+vrUUaqEEpN/8V0KNiqJH7mHe1CuxkDZZM7K4I2VGvtACbGp
4DwxToHVTYhKTpTSM++RQtjKvyIAsBI9ewiOs2tNplMZgokLmUCTZQrJ0oM11BVP
0Idt8iegaoxOuZHZYxwhpVTmo8khN7WZAhGpOGC8TrlrPZ1CXthEMMIK4YyPRLG3
B7NbRBXX/4ucfyD7YzlsQhX/ZumpT2srYrcwQP+DgX3NQVWj78OoUV63bzh3zvKR
PF9jFpuho29JGf1071ySWUtOmRo6WFKIxS4QOTDcXMlx7hmY+wRXsRZy/rC2hT3z
ChIxwP2sv4Lx+SMublUpdFMvJdpzWVgJQJ4qGM33HBPsDVieME0A9R+ysxGyt/Rt
V8iwgfTdxiozjiSJzSC0I8ipKZDuEcitQj5qfMwECLoT1BMLOcYxRHpWCIJTPmyT
6kSIhJTTmlVx5e0T4lYSAPdR1Vu+DLnUL1YztXCb2IjVfrjrvU9MlQdgKu/CTF5U
CE7j2lazZ0hlwhCf1TrchYc/y1zcVXM5J/RNIVzEZ47nLXXHkFxaAgPKapblbCi5
dk0qH6YLPTxn5TTW9CKAonijH0UAvYH/nlk8ocjFtbrtgXAZqvclys6wKdhxRPlv
1F4wwarvh64JeWHxugZkDEVN3j+L50yHfnuvwwJibDtSW9qIVujO6cwSDb7FRL4V
BTeRH5cdwT0wWXDnqd9B8f7PoQYrwZzZL3tDqkpoBo33tGHz9cJJiISqzpFzSQ0i
XXLCEqavGgtPnzHwoNgnL/qepV3kmDOuUgD13JV92AgKMePCWWgqPz+yiKF2JyXd
Zco0QSE7w/p5W+W67GX7FAig9t8yPrkgQ/5qwNp+n0/HIiSY+KXHzDjx8iPaXn6k
uBDNJ0tYhfLvLXJk/OA0QInj8n/xvOVy0QMqAG75fy8JqF2JN1Qko3UdkLA2zgVb
PxipCE0gE4KqnGpCxF0KIIRvXa5rDugZe4TF+iiCccmp+tl6TRCqdWIBjrK9wdPA
8iVhU0/9ry4Fw+JsFR/zLa15hIJb8h3SLWgXbw/Xtn64Qznm7msZy2IID1gTtS9V
9ivH3Kg9rG3F7LefvNiPPJ7sPwLsqNWLFMXk4ZByUs2VP7kmRHdJhOuSLd3tAi+J
tWlYOot5y3ok2s0bjZdjps0fDHnbwxsIK3igbnjyvcYGqjayCLLzhfTyQ4ZS95rn
eSAliR5RAq7ed7dqLsuVlDNLpmW/xQuwraDwpAX7HlFjH+soScMPpcBS1E7vxZoS
nRP2Y55S2vwqrr5rfOGSz97kDboO2xZ+S43zMFo1ViuwQo3q7CXWk8X11b/bgMY3
hVLt3XeKA0Y6iniqqTq/DNDp9759MDYm1SbeiggaTVcrfKoUFpHfvn9L0Bs1RjaT
jj+JYgmvFmGwdJlnMDrTgFTfABLohjDV4ncBBwIRyM8UNqiiMV0K3B1hMk7OJikB
vKZNI1exdmRv7Uc695FjSaJCSNqiZrvkh1Ua8aEw8tY/j4aZMQ4MtuM69tQW0mjh
ah51xKpOSihKybabJd2rcaeuVIpp7ik44n6r1JIrnstRKTzMFlrMFCcG/DRoCDR9
opYaA7XXAHI9u7GLbrMFl/nuyS4qefnNydhhIC0nQbVejthChTXM34B5/bFDsjjm
MiMohIm6dbm7USuDAhhFTvucRzkTRyv0RMelnQiwFwNXhO36Pg+qzQrGShGCcqHk
/QoqWQWiEHj+9PzkeK8tKvDjmzq4X4s4KFV9F1AVDBLeNx9bM4aJCM767JIH9V86
97i50f1JXqwHVudLal4ewPGu1yF7++c6wgWzPmrZbE7lpVi8tUOfRb6YOncRedJT
qp7P+B2MoDYs+Q9EehzaP+e5mj5iGUmvcQmFcKc0pmpjdRtzgDMRtqcipOgtDfZO
rKMWuxJlXkhD20ZnFYLCSuz+IaW+YAINPNmLlwI+9N1gHZx05jCL2hvFEY12vaH5
wEGzJoS5a8lPLS83qF/Dk6k+vNMUhE2nQQ8EMR1lqeWQmOkEoBfSn4jgcryUvizu
osHG00ukQI2hoytuEs01RsosztLRGkxBHvusLbNdA4BC19fwwiLfSvfj0M+1CJc7
ku35i3HyYt4AeLJgdsInVIPDFF0rB3SwlWSPNI8jkiVwflZAsn0NB+k7QH4jCO7w
h0Lvhh6BBZkKxl3ZzrHYDwkqu4f8J/LRueLBu9vp6HWEMkiSHSZ4V3/sDM/C5K8u
IsLFLs93q1i8j/ek9DpmpO1arnfox3Uk4b7B2E/+xd/0bW12EPDZEKnUmZZP0Ltw
Mj2iQcjrPL3KEfvEN1n3OrJFyBXOPejAuCQyDiRnRG+Nhfz8Xj2aNLtth5Sm8HIK
yUOMYsONqFzNwr5q5IA46Rk53fPBa5uQA5g+TOfh//1ZM8WFf5HeQmSDPAALCBDU
28JWz4S+toY7qH0qbw82Mb7TgjQRYrBazO0vBTiYCdW7DsiIp2I3PDLLhjt8dzG+
J+dwzC3iSP8bzkvq99NpKgGEiEo4d7p8B2eTuCpfYKfnZSi0NTkWNpmWXY2Iod4W
ag0YXFLW+JNnWbj+P1FYy98ELu7YOEwfr6ya9crS+y4heCD3zc8JBsGaJ+srcWG+
SZBrud+p2jJDo+0reQ+okEhkO2WiFflLeqHOtcux79BZXaB9q/+jv5HIwsrQyArc
LA0sSTyvrRt5U/9U9TNozYbmqLWMKZzTyVdsKdHutqrVfzX+fcZc8XDe7TYknhI4
FvUOyC6P7h5XOIqiYs9+dR3uK4u1BsfJnYjJ+9tjuxu8WU4gQYdbqc8+IGkjdLU5
z7Ka0V+Na5kr4/hosspVuD2BxJ0Lpr3VyDR5Nqv09t+3m7IBrGThidFeM+CaDyh4
KjFPOMiihkG3CGox0CG8+su61F7D0g1QKw2yCL1soCOWqeoK/vxrYB5BonkAso9q
cuvt877eJQ3H8pIyeMvoQ9JYAZkKICcaanTxxGD4fvqsNd+zsm868Lq5gaTMosns
EtxVjE8mn/5K+C+tmv0Vr2MQsUA4iZS+1EqcWOExsjXhsHlMp3+9766jrII9MKUX
AujHGsQrK91K7+qVsbV0b8MBTls0vrZdl/q3yGmNxw9GI+ZnQ5nxk35RNKu+xwS/
DvKxIyKmZOgPNisONy0Ux/MajGgLx2Vw5CAiWjDuuczEsN8m+5yr1JH7KjA14FQc
kZ8uKWko98iZJMsIHnsuJBph4dtTsByNFZ7afTC0k86C6vCKrlEdq0kmXhYCckyW
a5/JgWmJ/LRFj1OvyqPuovTZc4teHurJeKdMYsjJHHeJPo5YBeW/kt5l0rEnuBxQ
hVQPuRUWCgPM6Cf9lL6MafQElFI1OBMkTSvkAxujJD8N2zXp2zXP0Ur5ovpxsZ65
juGVl/uc/uqszWdvD99h9W3ksn8/mF8DdMBga8tkpIAO7GxsniIxTYLPhSCquWji
Tw+WDL/9DfwN8AY/hNebLeN5SwO1dOW0qdSdPCpZh+Dur7RuONkxqPSWTMR+X7bN
tLdbjG8WthDSERLnUA19mKUUPIPiw4WyiNdso4kCLb7ogotflEJPl6pCO4tf16dJ
szoythzEU830uC0GIErXhM4IBzKKRmeC0lds2KC7OcrAQkuW9TyuofUPnyQrNYe9
WwSxrfWkYUCOkUUbGJjFz9VYFoR6X9zihDjllPE2fejW1tVE26uYtuvrNzisHjwc
Knr4OLmcO1HyLDKdXSlisP/k8Jl/b6yj72H0awkuizfsGXlca05rMYOsCp5JN/Ir
idnkg+7Hbi+FU5uJ7MGJ5xbwQrB9Z4pIQX15jLnRsxSaGw2ptdoPjOWxAhgNU0a1
4UbeXwHCPKbnO0sYJ8aTFKV1FetOXbHaHGmyWXPrgS8dYg/TNeaJj9ltrSbMx+Gs
c8r7gzIg+AlPIFAX7VULYUpS9EgZsvjzmlC0sqtvlCg+zQJbfrLihEoslVla6YnL
COAzozzYaLss+VuMsqUM2ThDWcD8/vVKAJLUsR5L8rqRjVo1x5H5M3xm9h6ujzBo
GjocWJ+N8jn8pigrCG8cRMJ1/9px+n/b/zVmPEIzYOa+z1IFgK87JWBB9X8bFOwd
pqlIeRNaW274w+9vgAaH5wCyP94r1xdQiufzYp7xs5y6NoBap5ngDrSP+UJo/DA5
oE/vrwz9Y1gz4OWM1sWLfemkT5V0I7bqZLKoa08E0ke29GZkeTsX80ei8Bsiekb8
dq+Yaw5NxsKTHuHOEXyEfA72xt0CfaSC+raSxoHva/xdW5IuSzw3YwoMaj/Nmski
LtxQz/ooSZ8p0Ud6zY1cpaDl11oZhMfm6JRhzcXCDoEEd/DBbvU2ffZzG4PzADnx
LbTnGocPHkKSZAn1GDH46IR9d3BK8cTWOvWjykC1tyvvmxN9RHJO9yBC+976L2eJ
9EitEsFzuJ1wVVqWZqY/YYENRUvtinGZK7KfLmQdvQU6w2vS+AY1oRp0HKFAgQf4
2REKSv8q4anRzOhYgdMM/+faYpBwPaUwtGI0lhdNNI41aMnRs/chhtB6sl1J1lm5
TD50Osw2rhoCimG4Hit6o1Y8UUiEw2eHxE8psJ7zMrf4VhqtXiSZSXtfLP8Y9+kF
wbeKK3CQSDdQ3rdxLOg6hMfgiYIje0bvmy6Rrpfg3kLVuKLwsbcwQKtickb2j8Zf
bimhUB/vKO76mNtG4WY7Ns9U3R+7GUP9LOkvzowgmMBrjkrzPgFRxFElpanzX0it
WIeEdZ5lnYQeRm+Ni3fDc+99kaifEMwD1pFkHP94gbFteef5m0D7x3o/sMV92uOp
MjRNzDnR6DFTNTFd/v3txvs7kXpxuoaygw0uAibJpvaqs9GRD6ATIC0xdfdihm9m
zwgw1Sn0aiL/dYSjCp7iQ93JnoblAzfRZzHfwzIxWTqeiNua9J0NE6wsSp43wCU2
Tig6wxRwcDxVPW5StxfXEtQlJEK9dxbSr+Svl784cqyrMZGSHLjgQLSo4q5iWp16
uLcuqnwahyQJTe0cA10T9pWH4kM8bKtzmXmxQ7aZpPErL3JS8o9gdFSxYAhBS7Kr
nMRG3oGQcldU0emKS/m2SaZFcvj2tdFgDV72qivM6gVHkyaj87lgmelvDlmYne4O
7UFaR/WRa8KoAFXfORxzxalOIn/qVdvctuRU70DrV1ONVyWJrXifnRG96GfimOlG
xLgUytxjpeb5J9/pgLIIWz+jBfTh7lXBpH3UitLoceR1kCBF0YZY8eJF3wrJgtZY
KLoAn+B+tcDQ+v3ladmyX+DNaCv7NUgo6plr/1pEdwduznmcqDE6zod0GLtTXZug
9dtEDLFg9g8jM3t/84vVeQG2282tTErrPngIYOAG8oeaXO0CTwlZKGnep8BHXSF0
rAVI0rMTW3RHuQrJ0hdo3tzgVvOmmeknlWSDMdb/uh3hGB0iNdryqzfnzmO5wXyc
LUAe5f/KDNLj/lTJaE3HsXofpXIzWif+hnhQ/IZYD6z+27ASlsI9orHP6FTVOPV8
xtI/xZyyRgnWN3KgmOwQIWv4PmOb0cp9WhroRy83g5N4MFWGrlWSLu7vP0YLlepI
GF8TxJwz4UHqCJW1uW/0jK5LrTHpmMnlUYRnp3LivMCAvvbA2MtfEZc8TyighHkI
NTUVeuWBioaJFi7khfVGZBzI2GsIZMffjSe7ilktVC5wow8+YJG7mCgBssWgMbMO
f2hDWwZgjZZzRFobB4nVmAB+TPpy/1NTvpBkRHH6SIGwxybeeSFFGGb70fCSb5BO
SMZa+h1S2aVsTPbwcVZUFLD/7SQF3kREEqM5zy0egAEHEWwbuWTPk4DUEI0KE/4d
nWE20qYH0m2yLGY9NWHXTpGmhYoqdOmor/uVe1STGZWjAWTBAPyYBZhQUk/umvxQ
Y1gjv/xnVBQ1+EJA+TYiNooUbqh95hXK6fn1XWmuy9j+bkGcLSvKc9h2WqCCicbA
v1Q/JYFYi1vgqKn4Qc/8X+U3oClteNSgGDV3dlWHPopptmikUdSrQR29KrXAMUli
+cZeTIFtEjWbNoNYFeaH69EeJcIvOV0jjO3RIYp12ywMlqZVt8mbBzuHOFiLIIxx
wJ5pW4MVaOaSNN2mENthF/v307h9MiY/UBxRbXYDSZJbej3ge0DgZkgNBYJbHEA5
mANNLlJxsqnV/EFcsJ5RpVaHsIzvPlyQIMUAUf/Nejl4re0YuxAGbbcSLSPpK+2Q
u2hPWzNNwk30LsTGNLk/2/Qv2dMgld2vmJ6k/qgBTOd7TcKRRaCiSCY8AvFzxFtO
PxSsUuIQfjBSwwC/FR9mzRHSGtHtzJYikfDaeu9hlSQfBb7kGhRUF4pWem8L2n1Z
v0LUbsauQZlVc1TqkDYF8n9S/YjMf/YQ9hRah7c53s/2mJSLJCZJZ7bm2IQZfLxC
ojabmJu7TMdm1DiXKTE+bCNoGoayz1BdjrrT7xBbHP/xJGLYLdcGaT7mtscXbtVK
CcjdUZiGcN5XJfbytndVse6A1Skwz5OC2v/GFxQtBOEibh+NimbYSSmbnA19IF8V
zCZ0eUwErjnZj4qHen06qhxaRqbsnTpK4c+P22XifX+Z6XyoxAoYp7bWudidtynQ
fRKEZl6Z9OnRRC8uQH3kfRbS//994rDyUidARz/X/q21OvSY/IC98tOIYYmCNViX
m68aoJjMoAsUh36PgJYJJF5+Jnn3kPHdWwyEI8pKuJjkN+/J3DFYyAX1v9n7EWzp
kUETypDKseGX36FuhIAEP2I15NwwfE/N7b1LK2TNPeOEH9w548m9ERgQQ0ghcl74
QNmqlHqaI+Mh5ffkG5Sgsauu5z3KHhnyc9TpB60HgOZu3IqNairJRs+LqaYYLpqi
EA2ilLSBqgjKGC9SaGjhjv2d3UbxLnn/vJPWi9niPSwsCyN1CeG4hoSLDyKKiDgl
u2ChrNDNuFKd6tNW+NC0pJpLlNN6ma2HV+RiLrFyxEDD2/EhT7q7VUGohJymH4dh
+M7WosBulf3z8I/ggVJWe0aQrxPqIBr9v2eStxP4oV5HB0+trEAVcjdqZ1LgpHcb
aREPH7QHhvvGeIych9U8FPJ2hEa9GmB0V1ftMiJ8f4XOZJK8zWU/Ncx8cmHt1TWD
F0nPcGLC+h7aVEIN2efl9DJFlXVgxTNIJ7UQdIo6rLhXH+5C/+etXYNv7ZaccsAb
fG5H6VF4cLV5QOvtxme6egyUJPCBNV0uYpkFNPNy5KETlovQubP/63JaOYsKRALZ
xsB4DLb6yRDYaDxQOABYFFnvsroxt2rDW+HHbGdUtqRgjKR4GT1P5821o0lut3pd
hgBIFRDotzhGDl8bvHTZ3y8AlsmctCNZgCksAEEziBihDlhnUZrRU3v3XzddJ4aO
X0eoVF+/dnlcGpmLmUAyBBoLvl9GvASXCb9bNJXsGtEwmPssJ69kpdLQJ3MnS/to
FWElthokV0tZYNsZ84S2L0F2QoF5wrXDZBlSRhkAuj0CdTFVRv8VhMkq9V8aSMY6
2TC7CyHRgehsIUhw/Sxy95NDuVOhL8Ncz/9BJDPrWjBZZMZPJNiKm8HtQJs2dn45
tlwAdWvWLQ8V1bscW1zJajYb6JGySGmSdrATinTIhskOVkoKp1DZ5fPFjESWTWo3
ZNc6FWmUI49FW7vP5a2c1W7UNLQbx7IUWh2JcGXS+UIT4VFwrVWWM/v0ablKXxAQ
e15q9JJgtW2SO2q+TjbrpfoQ6idHkombT2vU0qt4hpkKNbYyBtpDruI/VwDblpft
qeHpFyQ8C7PjPZ1EDnWC8uzu4mJ7wJZDkpFsm6rsSG78S1J8pLyKFOIC9XCvZCq/
O/aFMIGqUiNev1k1g1WVRDAwtAzHYkGCrECeeEAnbAQVrVYcyOAtTlCFFfbEZCQx
i8HuM04O1uQaCT/COLiPP03atQrgO4Wr/vi6DbSg/evIE2wiavyI35IYObUrp4v7
F7JGCEYL4ik6eiBsInMORNsrsQs75LdXCTXSwbtDp0LZK6UHxItxEGTXlhY69dFQ
y8yDhrY17Bxm/Zv4Ei4zybiEL6OUv1l8J4OCZKB0+Szi1F71mTxXLjtTxnZjxECM
cyfRYgCUU2cnYlSF9PAIlSX0IsSJsYG/sEtjU4INSB3FDppxHsnQrqo/I3bXalm5
ZmDoPNOxWpl1qtUejHwVgaCjJhWTy1JJUzuVmAGeSj38kxW1jFGGQHVc620TJUNV
kNPDvlmZEhsb8tZrdinFgI5emNNkTJmi+9YGUgOoZJTxV02XaRlZt4b89UCHU4jv
OuTQOLxe0Dk8/6yRWBAKOjVFZI1bLOGAu9zicFk0BlgCgjQxqUh7tyGYS9tlPG7e
zp546QgqIPxJPqvvnxZo3XPX38QY6R9d6VBCi5MKX5MxSLW7X5cxgPFK6B3SiAa7
TauSiMkn/7aJIliSat0FH4mN8euyl7WIFTYqQj/SCUpzDyJzn+SnHmlgKyIKoiDn
0EDhuV9sLJZBJBxirTSkN83Iji5ZM15PvtZaE1t/M0kF2u9yvtZaTY2wqTBLZJ4N
c2Ifm8R7t/AaP1NsNJ1iehRXdejjnQVuywa9BbsA5furNRsgH5jUmDIY0J1aGHdl
G9aC1/fi56sIuz6W8s5gjgzFtpHnAbwsFGBiQ8yzYcMVN8XiCklsoeFOG1PjiNcw
BUa9YguR60RoDPRu/c3wTXf8qPTHzHpfjW8it4OzRZ+kVos44tyBW+Xydvw0OgbF
yPaIQonLbxuc3zHVdHWpIlrhmcPlS9Oxe3gU2Z43cMoWSPXA8HrrrvPAIhzNqbVX
CyyqbPX47cma4r0yzWiSha74hxA2OB6puctzt6fyohB08ehmhlL7GyWsSqaFOh/y
bTYE+o6uFIjItl1pA3nBAh0oEeEg13iE1b4DnW5O/KCV3aoDroo+ya06DG67RF5t
rns4n+7FPMywjx1/4IyPOQ1ztzll0Y1xdfQuM1kO8msqjbWdXD15cC1J0XbwgLzZ
honvRRZ1C+ZU+XBfNDHGCWPtoUV48hjFtoFvw0vtZmSueU7piA0Abq6E5IjlrAiZ
rsv9g6Po7ZHLQrAjr1RATvxDZ1FjNTLeBqwsBSDNVFmzKg7JmbrDOpmzpntDqZ8X
pbYBlzrR7/HyEo3lOPoTgpc1OFa7OIGL9kdHIdLp6kyNK9E+yng+dHQYRLJQTchJ
cRmqh2C4YQr9rfHGavznnk00dPM5kz1uV3LORPU0SJb4mYs07B/a8BJ37zmXAPHS
7Ohvs44WokiaG050gFDoKsSEprCge1L4sPqdohz/U24WARYTWGOtwdRt2V+QIvqo
4Ti5CUUHZaniMtip8SAETZbDfv0f0Y68EUDKREUmYsNY/lfdRhL/FP0gcOtUJ+9X
Ksk06oD4idMBQWTjffs3O9N+EFTZS0EgVYUgUf0dhWCul0JG5RCUreaaBKmeX+xU
k7cOJGCOh5SprakItvBotox/CD2pIs6AljnYh99fkuVjZi62mVXKEWtCei+sDqUN
Ki+22pXhDqsFkir40U5Xh3U+l37ikcAtQMXKfNwTAClj9t/c91IH1bPtI/A/op5D
yt5ewzi61HvW4LK2w2g/hZ2NNcObXm40KZJZUTHTZaJiU3iomoqnwp3rZUvSpTr3
N/gWvnLBShns05DsWIrxvh4B9zICHAk1698KRWilGkfHqOMipfHEQeoDMrns9WAC
FCZXykISs9KU31sz227bUkFplyPVsk/85tXFaBwYtWpxQU6yGBds2Vllq/p7O3yn
lRAQKcpG1P9bjuJ/Xe+A1fXbb1IeIJUw+vgR93Y6uo63svdVoFKjYgdWYnzxvJpu
gquQ4lndSmBRPX6rmbZHy5d1l3ihRCG2dmYfvQE//q00+qc8vRE/w/3Ebp3UJJgc
ZwFLxzjKWgTEgTBA2rIaiBOeabtkewKol0b2cKeP+9dy0hX5cFOPUoQa7RKY8wuk
RS1pqSGj73+YylEoCdDxIMg+r7NhdxbCIoCOXUvycAdkjyGG3KSZWp7WF5sRkWJH
817i+FiYLwlNs9w3GhtIV0AKMSkPyICp/iUIhlmKhrnJZDuoXxJ131SHnY+EO3yK
+ecL/J5+i3J4TkaTlnOOGsa1Ba+5PcUOFeVbTOKNHllVXpv7KrzwhfhL6M3bDikk
QsnjTk7Gj59TAl0bU0ay2tSxnnA05f+5+mONh77KHww1adrPiiRsW3VhemUzUuh9
MPC8H+hjBKPPlwKb0lr5Z1FoL8UqiTZbi9qY+y/4QhZKwuEO2133j/tJ+m6sRLN9
KbkUA4zSydzyoPSDhjlayQGLWDxDPwqPQ5TTsibq7GTGGI7tRv+VLsNx7THE22bJ
ykEVOvrvu86zvYeSuG36BZDxhYBvZpCgqUGqUBCS6l2V6TNZwUYXyAznduE8B2zw
jf0EcIRb3LEfObf3IpUS5h/yCSrsA30NgzVZP+iAhlNx6C6pPJEFQH1H+Lztdbbx
FdEHhSoVPi/R8u99DQ7cfNBUGvCOW8V1TqQ59Z118K+FDLhV/mCN8CDPEDotT4pr
SHPJRH1vGpeUtZNMHp48F1gMb0M1ErJICV/MhCSXCSUGFL++j6WTG1MWIup+E5En
cbkP8TRTmVYqxqukUr7T6Weifg/JI3jMsijfFATLNP6zsQMuU9E2myZ7eYs3KRD0
W02woiylI7DKAEDFUXfvUHEZEyJeDgSRQEnWc7NzHBgRDjKtS5lXAPPHb/MLm3n9
Dv9QGz0wzjI5XbbKLmdkH18fRY/3I2nJGHkYKMiayrS2tc6dOSKId1d8PJPNG18D
Q3vWWV0k3kgH5SMxvtT6lb7cr8kh1CBtxTWgzc7AXWQ2IA1wdMnn/jjMhjA1txfT
iFlcHPiVc9Z6IIX4r4ntbex71HlfzbTqUarO01RDI8VsqXOHhUOb0a9eIvEiBPjd
jevHWHx1iUqqR11LdT4GCmlgWt6Iz5eIxB0o2whbjicggcU11g9D0sNp+XtjIP/C
FqQtlhFgH7q1rgZbdCUsNg+kjuJa14oqMDLjGPDdNrP54ZyRDeBzy28edpo7L3TL
utSBMEHRzIPakyv3h0YcCJ0T08CrFdDXfcJ+3hb6lTN+47mHz7HyKmKdxk6jiJal
00ulERXDzQm5A5eMsCCRsdLBuZ4ln+spQ2+cXtZRMQoRL2OEX98L7pFOrhuTar7+
1w7N1lvl7uYz1/neDXOzovAQj4A3fY+ndrrtKcV6rnnGU0NhB0UisRyg0HxoJJl+
c6qTvm7bYV3X1QbT4hhrrBFzJgsty+uG3vpXj+m72Q7paxF2/oa439DTAqH/yTpt
xw+YWxAFW+T2E+NnHgrWfFUiifXhrqFZuaYq7sIkXlQIOJO1/I+3IntFvpc/M4C8
d2cQROdFrlQZyAgI03dzbdp1Rh/xWfOKw4guyjfFOK7NjuFkg5XWfgK7sS/4YsFF
QJ3BgnsHk9N0lecB13wvtQN/akP+cg/KRVikxueFB/EjeDn/wZVskk3PlfRcOeCQ
X/4vhGTjFahheijjKF9NYGhpcU8mDk/ycT1v7w8JnJsTtLN4pn5tsDAyaW+4dMev
NfaIC+hm0dRPx8ebjggxOpL+h5E5CQojsELlpQKSNrc0siiBWzaItN/3FG41IonU
FqquPwKLoKCijo/6y1xuoqWuxsyczcEqVw4WDffCHZ583YwPxAF6vvbh4aUgSXYc
q7cKeYDPf/cVkwVT30sUkpow/BpfvCiVa0ww6yTJMInr3OBvM9EoxkqdQbqIu/bG
+kbu+71bGIFXZHTmiPjm/UzChdYHmYo8rZhZ0d0OhhCsaWpGg8CuHhks3C+qXxHm
KKN0qBzMf6cjMWKMehiugXyJV7rxCIntwwApgP+b3em9Uf8MQdNTnKwp0JJlzQoL
FC3GHVI2YDc6xsDBx8jJpS2wbOX8pQPiHdFoFT2V9wU10sysqNGcIdXDX5zgiRy6
VQHV+AWciC2JbeWQ8F8DuVrlGZxUxIfGHo3q2KtuD2B3KCgs57Rdz3MfNL+81rtM
YVbZd3h5OhzJemtqz7QAHpNN6/KPxdUHGUvLfVMh3WVgHaE1K4iGiovOppyqp/VL
MHHkP7cZTyQOGeaeYmF8R7rEGD4k3Z8prx6gzuWdSyfpFwTwrwiV8fHR7uGdYrDj
fvISWhDFhs5t4ZTPuV0kM/bVzKXT0Y88tMUjvGYY5xz3QCyWofUu+58b5t50j+OS
Ns3QXX+/VVzoTk3FYOiRqva33sEQs4uHKjwVBG+1VB1tTDNBoEAer7moSyUkeRio
focH6MO2Ea2tT3mREw0MANx7Qaq9OuWi98TDnv/uk/Bmwn6YPfOj7pUufayIUPY3
m3h5spI/KaC+12luK0MWz85EEMwAsco1HN3223S5HFeT8LmKSjjKCkA5V4lb/Jz5
9PqZZDhnvs/Q1n+h9wXEmsYmFSzqPwgh6xtw8b0z4/kmWnCQoLDaYYzmuyUF7KAY
MDF7Bdzc7Sm9iesjdcrqbIja+7j2sjRs4nVfuZYm/XrG21tiKKX2xMHbxxNp5fEn
3b4dYd8HiKXQ0YAXNUNkXKFaLBFXjcKeISYAiIbq4Q+FFltngvyNqumubZvC5rs4
09N7qLucNXDqrsWUp8ZsYOjBFanm7iqJVmNXKl9HjjpRNzHpEOn9bfAYD0P0vaXf
enS36EVGxVJwQwp4zv5Z/v+k/mQIxKG6f5Z4h4/C3o4oasG8iLZjaK8Cvd5KKqGU
uHvBTtNmybhIIuN651dhvA9TgsAvm+BlTvdJj4VloFhk5mNY866ayHd7Vbz+bo2j
zv7gauZGfZTie4VHs/ClHKhMbIxx6lfQhLbU2DXx44cbG9kK1w7pinsQp84OKz8F
vkwLN+Gt+lPZSoN+vOMEmPf9bbPtnIsvtV8/8jiHbU5Fs3gQB2K8YCnxd/IxHonE
mace9S5Czq9mQA60fFUI+65+qt6JC5L9l6LQVSryvUk8DnqdI9Gtk1PxxmfNEl5B
BtKR+PbY8M71h1isgHnuIVfXzUf+VVf5iN2dZkBVD7G7zAd9/Ul12ossl98kLChz
lXrZHvbTZdRQg5rp7ilfRfRuzUD+DdnmKsKVU1yPvDC0efpGz9lNPU0ijAg7vXmL
ywKWgxn1USS7sg1V5W916DfO1iNKU8E+ym84zbMn9t6boigd5Gd1PEQH6hgiPX8q
f5w8EWuQPr6jnst1xikEvGzPnklok3jSx7vZZa3J1ep+wAJrwjO53jwVbqi7WV0b
0risKAbRIxuCLsx6CbUtfHyuELRZYln5Q5/t950VoI5TyA8se2KHPF75B1TKtv07
bpcAAq3a/H/6FBj8/OHzhZoW6oktmmw3bDAaW6NKLxopxP0K02qkIEn2tC6E5aOh
E5qfqVu0WIWxHsa6jPzC2evrNVe5ywLjMlLlc0VkYiFBJbZFeqVO6Qf2sgLLquwH
rhrC9XtT+MAQZa46IKZ+DZ0Ep0qN9nVA94V1TrBaYxMrNBTilRKD/lRwGgVMVoTc
LgVfSfIMbQldPy+KB/Dv44a86NqtH1SwMsBwH1zrtV7XUzkSgb8uKESqtQ7HUdjr
3ZRCnfk0G3PaoIcjWH2yVUPr5reWZYt0W7Fxg0/zfrMtl5DZ5oObfm+0M3czgyuQ
NOnK5jKIGXNrfome+4Z1DrcC49xw01LBeW81jKBtdLI4iiYVVWWeWh+mHux8vFFK
BvHS8xC+ZA5YXU/slAU9asPiE0EmqvjS82+1YtVay1H55shZadjn6XpSdztAQSmA
ntkYO5wgEjqJhqPY9G77MEOjXcLYQh8tMWoD8U5enUIEpL/J/FgwRM9SuwGUMfAr
+IIzIjR0FCOFHx6fUCyVPHL61mXxqVy+lQ3byBGy8jn/WZ8WmaB5rbdc4LidJ7II
/mu96RPfZzw0kb6AE0OMBJfHQSgRvcbPzO19BpigWeVpVT3LeZsm4ieMetAV4FOX
qg8E2uvXC1EUnsfm7d/V7B7r2V/HLxmQKMsixp9UA2oF3lowkdpz/RJbUx1rKWzQ
R3/huEiI/nd1ocqIBoWHoLc8lQPKLdCyMpqntpL1pmcA/tqEnG2i6GbSRTzieNX4
sTCR+Nf0IkLssVLeJ+8spsMmvP5KmvbiNusgdu/Wvd1P1cZbbbWv0R4eSeYbV8vc
gi8rVrKvQhpitkL9j1eYRVaGSTkzttGGXNQD9YhfeUTFi/E2lPwwJwqtZnIiu1j0
0/4WwClofTxGpbiuZczkfqPh3PQiJSC5+usMCZDZWfu7E+VOwo/gDGCssvMb7rx+
z1Qrntx29Seo62zHZXgvzHTxKBNAnm4td3GRXkLgluyX3Sr4HIrAI8ba8E4cehFM
fzuYsYlhwpz0tMTefiwTKCyVqhN4Xn0vkTLksCLQ8N+UuPUC5IVZUE841gbi3XYu
B4YGdLStEV4B8lWxTKdo6TwTcXj0Sex7lOo1KkYHpdxo59a4bU27fp/pHipWIgWX
cH4t/+BkDs6pwP6UOMM2ChU2GGMAjpKgmTriqUKJO+dcWsibO58y+OoQs9uou3Nv
LIG6vGSUp2DfteZ6uMWuSkd6vt2iKquZYc+5atN+WNsIXw1K17Sw2fysAV4+EpXX
uFUFgtIdkIvANQ6dhwkdpAQT2OU/nHugjIf+MXuBhh/QsaWp2clDSmPzBbYMZj4g
/yuSVFJ8IgsrI/IDepwwwnYBRgQINbYujPUyMkY5Tc4dJohgRdCXY04GTrs1Kxwz
Xv9JWoKcHtpNR3Xv1MyQ7bXT3qlKnSzniTau78+m2APKXXBqhQzN5RUIJW0Ib0Ti
95IXZEAvD1Bcd45Cw+rbSSjVSMbE0rokLgdT04JpnQSEuIl1cfTC7zUg6BVNb2Bc
bh3hYNAg2Dro3Mcjh4+v9qWI3TjEHgWxK365/U7VH2jstMA14uKNDkENbANyQEiN
SeZ+z2tNj/5TGH5FmjvjE/HWGucjtJ4IRKAz3FLmnEnygaT9cYusr9ULhNiz28dN
0XIWvNC/yX7smbaIYFrllH8jqXLtzWvqWoRq+6g+ScHwO1gC+XL51zZdCZ1kBcyS
6beUL4PHmE2nEY76iivJcy/0PQln8Mfx9LVLSEu7u1Oy1HmnnE5MN8KxwVBE8H8Y
tXAIOSwJuaz90NhoPQrxoHzYil4LQ4pd+bRKj+A7Lycsvb3n2KUy3DCt5J718IiL
wBbHIyeROJnjMLEouWQj2ZZw/FTGQ8U82iXQE+chjyBuUxhmb6FoeoIhgt6NE/aI
zh0h1JgKSlFPIr5gq7lhh+xrPQzxPXhJfHGnRRzDOYIY+2SrGqEM8xp9hu8d5WEv
aJ7UzfpOdL6tiBwK994fBArfiQI+iZVjw+NPPmMUjgAN81YNSG4MwMeMcJUy9mvT
WM35LGbPq9Dx3d1fgh6LUK3RHAcmAB1Zk+EPFIDCttEE4yNO3UdcNxSFahWDAVkB
i7s1IGcFlDlRBXP802CtgTrUpf0oAr97/WlPErS/P/Zwx7Z8rIJihrMf/JLle7DY
q8cgC3AjxCws1om73xTIXtcjpzfja8jL7rC1F3+Pbt5IJMljVQBU3Ohhoq7+FGhl
m303+7SdiasG61QVIe15HTdu3388Wh869H36bKth7mDr2Ku0KW0YudRdo0lXl9yY
ynRZfYX9d4OSfv9oSTZrlSdG3ARFD11fSiJ/ZV0Ft06MijA8HBGgju+YddaUAWQ+
eXVpOjJ7ZKLjlB7t4mJ6x/hZc+xvzAVk0ubpysuurGrOE297s0yodDOhY4XQdVD/
TueRBdlo1H/6L7DBTe0ZpK3CyRMcHU4ufd9nn2eiteJmRkN7ENegQgrEmusPQ4/D
G0bf1hORe9tVKa7b0xuQ/uGuQWGZar8nFUSShM4Wfe3NI165vmqbkqF4edKwKRHv
GV6EmHnZE7+MsQ/Z/adw87WDOcnKRhLPW3yBREsxynm7k9u47LR+AuQ8YDqBjIaa
vHt1G16E26ZW4ZKtbfXb+YzYHPiuhj9IHeun0YpbIJ+d1iAbfKpQvR9grfGufJFV
tUUB9sQIDgn3tsjohTOOGVCzNmobjk0EqfNKy10KDKqL+mc/WOyRpz/y2Hhi+Bf9
huGeXoWiSPKuLFEE84F9KFzRooy99kLJEHCvE9mR1IXKi6VqIrMLS9Y7b4mKwqF2
orfP/2Nww2g9RLSJNAfjojb1cy9bLvnn5lRIGGtVqdRbJD24NHOkMmnl+1fAI3vc
WgiwVi5YjPD44pTmcewwxlx2k1qomnFbjVKTipKud67fOoQqPC+iqVhnCY09YiHv
/My2bqDbGKhnXJ5pnsUjfJ6kUo/tgQCEE9BkiQfeu6u4pRvTt+61zSl6zBR+HHHe
SRERhxfX5Fndyhw6VZ9j+Ocz5Tq88rMRGXnKTCFcDzXN3Vw2ekz0DPUacGHyOWmC
+ngD5hn95TWX6toFz/bBMmam5UgDIPwVZDO2gpusNG8WL5UHqfjwuEdzq5Wwq2MZ
ShRY9WhKyUXACDhPkJMQmKE2gaFwPTYy6yde8IpG1WyLfIgfh2fnLuOy5SpMKWhx
VPhYHqdkJVnEmoDNtu74UZlmj2uHXTDP1UnwFEPSrVEngC8aR+skZ4fAvgpJf3EY
diTTCnQ0q2OZJukoF21J9bye5LmAiikfQ3Q0zwVxaCRCychf9lRilPkJc4nVA5OD
S/MJYUBCSyHbbRXSIScFfWkFyTinjcCxPZzCwK5B4Y4QnSc8MogGjG6LFWqXpi27
SMnKLciWaSJ5OojaQiXth12EwN5LCns3Ow7o8jw02FnrixKn6S33K03Aomlf1O2o
UsvDsGctKNl1zcc3J45OiwmqUHhS3dJT/732HFoIAmkP5FyRIMlDIGlveHjfUNrF
JU6dKT8/Eeg2mVn2QCzlsFeJUlq+OT8sJhhjrsHhPuv3b5m7mrZ+2meJx51fCVXi
iEjEB++nIbTTacTHNs1UNyPpfORIOVU0fGv00LUUYEHD8ooDPBZp+NoPGuz2c+68
M/Azaa2QMHTlc1XY7ma+PGm3NzkEFPMauensAa+9rCYyN2FFGTk0YO21ONZ0hX4h
Ih2pyNThrr5brlumaXVMXm6UpoPR3ly2aySJNXPuNw9LbPO4GbqozuOXiXwc8tJH
3i1iBsKlzpvOEq1uThyO9WffDeZWwTvNxxYUHRztPrpg9IEDf/BqEfxnQocFpei2
7gUWnQ5q1BLMoFNoar9QJ/0NA9YA2APqpXLPD/2230V/zhV8b7fz0+3XajAm+Ue0
MeBZFCodYp1iyh5Lqjcs1AWhLmenbDfxjhJxTptv7jy4oeEZVoeN+uao7k/c21dt
H9qHZbbXnTJCxBrw4wQ71cnCpjtqb9Gxf7/VuEL6zneXQDgAJ96ndmyRLP95xaAD
srUiHpycndVuVmJDBXTEizWHnG5LWGHqxnNu+oIsaJ9ErJst/SDM4LYfKokxDmH0
0SCtYpdVw527az5vlwed40rnJ0pZlEVBUvwOVaKJOJB/Oc9Q0InhmYQGd5+mktSC
NOu8ZXFguUUbvZd0GW2jQucsHOijKO9IEMPzey3LGHmObtpjc1oydVLvGa0DgdEK
7e9J5O/1h85lUn91gLRGr1wMdpT9f3lUvlY41YueHpf6Moyqel1pwkbRqTUsWKQN
KUUTwhFWje8ClKk5Z1aXvEr/RTut8nBllC0Zg/aHQ9fNtYMy7gBOloOxn9snz/RQ
Gj6mJUpdt24WBCD6WGz2Nn1MGPNHVbpwBUc2qK4nb9lJxmkmIbnhIlFqUDroj2Mh
mz/2aXSAfnRb9kgfobBToGkpzFdMSyqMbCqE7t+ceWX7i1bTtYo2eDxoNoe/jAYe
PFcoeEf0Pm6AWVl2DsT+qF957eNLlbM8E4T7xt1dr6sgCT4nA6lHUjEy5ThUR7A5
whpaLnDC7LIZ66r2plmOsT2u5xI7iVs5vyNUbGqd+MjRiR2NR6EEgVycPYPlPlXT
E8jCTkv7TybfsyZRFKj/JQ7l6COpMiG1yw99+5wBhAHzie7MULwKCokInGpvCmtg
d7zAUwMK6PgVdNbugy/CkuvTIh6bdoRONBbKcMbDznjUmZX/YxUGuXml5YwwM4AX
OEOvGbyvjCtfba8CjjmGcsT4H3WF32qE+C+jQZku5wGd7PmO39L6ECmP3w5849PO
xjVdK6QkbtgMZ8hmtSAonWIOHCfeKu3fGAoJhlh0WakZMNC1hD7Fk0zofAz+LGYV
2hGPxhsGW5hvCsi2nMckPRP0iliNyLHuqkLFPxRM0eGAwxgJqPwzmsoTLhbNFKr/
8tPxdVMUO8q9ho9aVwIaMPJJ43PqcBcX8UTDbsqEgtrGwMSNg3BGpg9nyMffbxef
ogh+2FOM/bcC6+iNbHWtrpsw0HezU0EGURzbNa0UvGyDAYEAwraSgqoUM6kt5qTB
YU/AjqwpjxdRlWoHKQs88cDVk+xD3d4TSvmrrZFVUsoPPLPTqxh2o4+d9UQouS4u
Y8gz2nG/UPMmgGq7wsKy26zTeCRbooE3DhrznvmFMxIKmefyuIiOKK5tR5xNm2Tf
xz2zq7fu1hzASjQHuygLoDT6RHIvwN4aaLNglpysPyfYvinBo2Zh+iCtM6LwdE3B
PThcWRGMFIXWVsQwo+jcSzmb1mdlujFbPyPNeYvjScn04nhTbGTk04DomncvqSVs
8ztrl5iZcqmDuWpKMgYkqK/+ZW6Y8NFkz8f1btXIkP0pnefxXa0C55ZYw4HbRvWF
ZiPTL7VELY80xh7p38IwPjPSQlmOB2wC9zbjtRKxYaVI/32quHV5G2BW5zxUG+YT
y2l8BdHZFO0x/HmYcyE0MxU2M3Mv7G4rwNb2WOzyjIocAzHlKpF2cn8yO0GosWf/
MT+gNd8eItX50k5odD0FI+Q6Kgr3BJLrpeHEekQhli/cdst61ExoWUUPHIRc9QR7
rETzH6+WemuH+LIvNG8bP+zYPYXXCJXHhQVJ7o5q7XcfVI+wE8r6cWbdDShbxsK+
v6MNoy9+Dtfff4Kmu/uEgrwO+wD2hj7+WrW1okVvntnD2IdmLhj6aJm8CnYDZLIr
+TeKno+3jFt52U1Qq+y0QZCKI/9lBGP9pFt2rjj2KwRmiGBBqAWfyAJtWs5FbrRh
CYO6NNTvqZM01U4Qx1mvxvnxeJC4EQY6k2gonCSo1dAfPkvFjCoLOEOX1uN3/ZmR
u4EFF6qvWd+WWPhtkNMjqvVyLcQi1OgfwwSFszM3YHKI0FxUU6gOP+5DTCZguDwW
sjW+xlYRXmE+SuOBw18VZXx+v8eb642i8HgDbYzK5M14ytiIkWH4Gy6uv2vwdNfx
iqIYFYAxEU51idrKOkpLeP1qNxp5EOwplyWSx1CxUfmtjW/9B26KVEB7RWvzjIz8
je9hcpddYz2YyuqWVL3jqHYdNaglu0l1R1zsBAPOiRda0M7qVhJFZPVt/JteNmeM
eiwARCOgPnb5o1yX3ptOtKtOo8j4OaFcttYwfEynzNkrc2DEpcdNgfvP2CzZd1ej
V8OEOA80ha10XrQy1PVEbxJwzTwwUXcyjRgdZVK54Os/HgUosFTnyzWsFS4Y+ajT
dXgt7gJ78lnLYlfbtJjXNLmnGWCpeQBRcyL7tzCPupdOkPZ8vg+W3y5fiKdC/LPx
PmrL8sEo+6ox6O2lSlKF+lTQPdq9HgprqMelublfGBtWpMiZnDj3vX75mc0MYa8t
768B6zvYWOafevJXKiWX1WNPu1xPTeRFYM5LxY7qVIDASUMX8J8s1C9BN54v5MgZ
HSeR0jbYbK2nneF+dju2L7T2xRbxcuPAeVKjVfKep/NYhpbVSprwHtWKucSXFl7l
yPYHN0KbIcOvAkFnq+jD91iTvEb8+4OVxaJISEnBZPM5eeTTfhLvqyy6DHqwBjrh
vqUwpA27w9+JB65yM89an6qRqD/AULE0szu4YFsF+7h3rHUGVicxyQO8D55FVrPi
Rrgc/AhibOV0D3o8xNRBgaDy6jnNBvDutVLamm/ZdSPfXE/huxCGInyxib4nCJqW
+Juz+JmTkTzvFI3dcHppEGCoQWzC2TSkHLEV9xh8WpzjaHvZQzvZTwYS7fInrB1L
UY4Rwc/eJU06hV6XfjqKaBwp8ys8kwbA1Gjb6z2qqlxwDdTv18Uz6dHmWFUN2P1m
c4TCrUt+0EoEe1u3MfozLnO6QGh+VRBCFKfIn3oVDbljELafuy5LG680kIgKfVPs
1ck4U1Vk344RHGKVvGLiXEGWud7+iJmwvcTR6TCrUUCRgaCx+Q7n7mXbwJHWCsZ9
fZ3Nr9C6yzBIGY2vd5X8WKx4KIIJM5fipU+uDPzASPwnfFg+CCjuDCzRJFbKjQGb
hUXnCAbLM4nuXIY3sw/nOTPAla0pe8a5kOTjnUmVcroIZHiUukHnRftnsOj9wyBA
vFymMWUyx49oNG99tIImuv9KgOs3pH0EC3y3W1zNK3lLwlxqAwggOm7CYfU8a/en
iXXmbtly7uSLb1Wev7tgW4v6PjD9QANk8aJ1VgYdrsyJ54uFvWv67J5zWINtk+nP
qwVjcsMoldvFwoTMfIJOnIkrmb2ZlSGU8ebyC2cQbphlLNJFx023wlfvqE9Nrygf
gFwbeOD/caH8zsuzywIKpZX/tW7tXRy+UEHWfYQY+yv9VCGPNJRGBRhxp97O5FA3
Gcduieakh5pvxRyBkFDhLUxo+BAXWyOrb8ad5b9zuCl3WWRItgVMIz7bhK08F+Vn
L0T/Nf/9mgYToQbu7sxYvWEMiVtgz1m7mooOtNEHM04kzcRV56kb16JpiXONF5mZ
dVjyt6KPW5HVTd/qjpDTFpTngyV8cNmXd6GnhXpmjSHknHg8sHugDIAWAbi/lVsF
X64gyzyZaK2iqpyYMRrbdeSvjaSK3TdToMEIETVH63gyTzDB704zsAygqb2Yj0pw
DU7IFan3Q3tOGUnSZRmC6bsdNBG0jnenUd0O4nhxSiBQpR2b678MCS5A7w1FxRzL
tlsWhedQVvkafwf09GrSSCdap4RDyEbPpGIxZ8lZ3hl+wZH54wvpHS2pShLIu25q
yDnRdmurhzMd6IWru/JLQWagtF7UZqF8h3vodz4kjwoLlnWo7uQX2mrIF6hVEilq
SuUSGStIvUvktRm5JIBvwHZbdS4fVNKlGzBmO3aZ+ftQu+TI99ojdXPuVlLXYu8b
+8Z541mRArp6Hqib+5l9A6ksrL4uEIrtDdno5PtwrkWMsquB/u3wfRJ3WOBgtFgf
8wip4rGI8aTxHeUKMwmZUmHSrC25q68zK8t0j3ak7hZ2uuxV+SWHOYFz7SmrHUL5
11OsVtiXPPAcYhLgRr5LKhtecmmkhKUOLp+VmXoac6AJKsyphQ1g8NMnCBLw8oyd
c6DwHLziMQvmcPc7QqKdExOnm8e8PzQAda3YsvPW2Gli64PFuesoTYjTmmw8+o2S
HL9v5daBkDmd0kA0Fkd7CQfE1o1Ct7vteW0DW8dixu67Qy7/eFVC4bm9jUiYULyQ
DO/mDMRsmrXfcljy8EJVSV1W5q5PbHf1083j4qKd8Stp05wP2E2H9pHJRdRRpPqA
5AzHzspTvh1ERrW43vgOJeHgCgpaXj19cmzbfBh6VTkDRBeIi3zCu4Gz5IzIas8L
GgI3O7UN3HZmJWSuiZcbQRLGndqLbaHBTnnIav8EkIZuMKjqaZisHjwdmpp1v34Q
Cl5Jc62Rlvkst3cOJ1UBGto25/tiVgP+bVqdQlT85swO7q9mKPTyixvyPbanPhKe
tfQ31Cc2UJtVf5NXrg/0xwiQWLtX4rr3DUenyug54crwpoGTe90DT5bO4nUgIVXH
WZixcmVtSh7tyJxVwDBNSmsptOHozFEGiBgJhABw7DxLPLdAXpg/gB/lWpn8XTAF
6iosrdnVjCLBJCY5S7Hq6tdmRLPusyePVmu24BNmZTWy6D3uX5KfUcxmBkVpC9nk
ckZFjPFqxZ2jSEVZYsYWf4r+srfKZi4aB4o/EcUvdpw/thgTXjuiiIBwV8P5BHKO
hygcqSigdpq9ATpx2qx5zzj8JGwNJwAxbcvjONovIFmrsqhvuCdZNg5pkjZ4R2Fu
mEh6Z+mScItJ6yadfkrgYdUZh8HIx+9B+RQp+FyH+I5MXQsJLJPV8IVnwzimUGff
9oSJl3ybH5VyhhM2fVjUuqTnmYQ9jJjxaPhfXzeN8lBfLs0GBHS989bH6DfWnI1T
CWT3b4tVYuFcIt5WM7VISdha/hfkASo/o+CzFx5VEF9jeLXiA1aNbF+y4svgzwLQ
pj/mQZUzQ+BC8JyqmvtXB+iLkGK0gM23/VMi4gGAhGHzYX4mLBLxqZDmv6r+s5RR
JgFV8fUpmF6dLw/zvFz41pXFVBIgPpesYaNo91Sv/NH+ePZExDuaAhaQs7qbunnS
xJB6ljrKRcgvIklx8hObM+t67tBrX6eiVToGjJ0thqw57mK/dtqcmbZMvTYMWYWr
7fXvGiXjIqgraa91ZHeIeT0lsve8cx3WGnnP7E0e+hOf9HFRZeG1AuLJOzF155wS
ex96idJqIpknfqH9ygeySFDpE9C3GlTqx/KKatl6lSrnP6XwBMyoULZYgfiPhtV4
`pragma protect end_protected
