// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:40 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PUiaZ/73ZNPGhri61b2swxWzQnZd6yNGjUJYA4L+nHIEb1Vv7kuIn+SBcIfULqg/
sHnC+zvyL3J7ZUJwAtLYosbCe44N7/D5MB7QIISUwByq0wnxbvc1O4MGXkm6/ufk
aOijmaChtZqg46u82IqP3lE/HMEiF9B+fk8Y9i4HrQk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2224)
yNNqJ35GkRfaeE1CyCfy9+MxIbkDeV5P23aXrU2vksxe5m5YFNiMS+BKkSnth7Zg
WURyzoZ7HSDlC3wo7J2/8lPFOCGgAf8uj8xvZR0+OgG7pLLHTu8rULDsx7Z9WlOX
Ux19oSQACKYep4pKPWWepkKFqbTd+OCi3KTMnMNV28VrvwJiEbeOtNlEAmF1y95t
2GNg2r9TDHfo2zyDqGu4UQ7xCqcClnMTu/uk34zolfh711r9WcfHeKPDdzmyjdcy
IriK88yvPWgWKRYdDESDqnUQoGdYvefvpbws7xb2TtsMmXqp5yeaP5xnqO1hjeZS
QnJ3BHhRtC+fN8JuBZF996fi+19pgbv8vL3NsezrzJ/K27dcoy3Ws3rkS0io5hS3
mzSU8H2zs1TgBjiA4RXPr6m65qSC/9pJePkJ6VKn704EVtW8mkBsTzzzlf+QixIo
Fgm1B1OLsvakcx8BErSlvlndPx5E6DB377rwSFpWE6xLfShH/P2/WaFVHo1c8bRw
l/i85nPAcTJLaUS/028iDJDYEVGEmY+kbd58V9uEOnr0OGognVOsMO1q7986Iluk
RH4AiNLSv0QPOWcMsx5/X4bp/nxtRmr1mPkvr4knyKM20GJh15bpV98uBMly23vi
qn9Y9FoAYXQ2HMXI3ZYWDUGz+dimB+ye/il/Uaawr0SRl+deOlWbrr86xKMIHX+I
rkAkGFVDWvqh6uvOm5ewa2Ccj5CXtBmupMHgcpBjEJYzM9B44DZN7mjdD+QnZOuR
PtjEY+LTJRqB5qRE//WkWkDGAnLLvw0ThbUq8LtWlwbMu+hbPbVu7oq2aMhIWamC
klWwUUEXtFSYO7bS0DK0JN0iHS9INITOvYUU1TNcD6CEkHfniTZEH0wBjDhp4Gng
5FlbBeHyi3PwLpqXR6GATIGXvnKYTgLo/ZwfmnN/0DgbzT4/gtIJxynqAEbdC8+p
aXFMb10xL1bcFHl83LWgd55kFcnWFsc3WET2+MQwd310rb4Q523hS/glnZuCr/Lp
LzkDVTmdRJ1K8Kw575QfqkrW8uOGtxrCsNjY8EniTPG6v+bpt9s8N4/lEuDwjYDF
sSjBqMJG6i9hs+DcVquKqThLwii9gbCUEOf3sTr4dmze30FyU2/8N/F7fdSXVd+l
KD7TNtLHYO5w/kRRGqTASWIqARHpWqOv6MrKA+1z2Kz8Xirk7raTFFkxb8te9sEk
IwpYKFA54m9Gg8JZ7hM1zcLubi+oOEdy0ssExXZXBGcHFZQf72Mz6VZ4MompI9Vq
an/f4gmP2kr1/xjRGVp68Ky2xj09S9IBfEc98Tf2GeluHkwnEWCNE/AM5SMs1bwC
S/uV/w/1bvCtCssltGSBn2CwG4Bd4jjmFsSCaN//3WTBa4M+XlXjU1b3+opqGmVI
od1BYIrEaPh83O4fl+mfMUdh43cYSZNrx9tNO44VGVG+eCrUquWlN+EGcgiqiENT
HKjiZAH9CNAQYYnFmzt4MBYIYN98jv9qPB5wavC4gREm2g+dcu0GuPgHheDCHCM+
7OmvdAHJJPgC/KV67Y+rXS1YN0MpRUg+p+Vi9GgvT7KMc+72puMtLfcFeQMD1nDq
X7FDTbHKwAQgGADDeATOnNN/JxvBKRUMJwap1OBpAEFI/gzlNrwEuemRr7MQjM4D
k6HWZUM3J/RhEWeetpcWMFPdNP2/IVD+jq0SHm9y/wYuCx8avvqtrlYl5oeN+H+k
ZtqJctdrr1nEZSv5SQOYc1msoxlwhB/yVs6p6UtFg0g6xUK+PVZi+lP6BbGW6ZKM
7aJU43PmJlmoPieuix4w/3p3q7jHX2iZeYe54q0SfON6rBbw9N/PXP8CzPeMhO9f
WiPUzvhMI+AJYSiAm15G2ik1lnisXPp7Y0oGRTTw/0mK+sVXc8LqB/6SzSCdGMiS
dusP4Zoz01GAKYj8xAwtf620lMnWay+hEL60JVcNWh6xCDG0VtXgvvAQ22CSU2B8
wA9QzOwZBZ2gKvg7bYGusLLWXv5X69KcheloOOe8mj/UtD9hw64d3Ulpt97k7WBD
fzh+70W0qCh6ZoxAkw/6IoW0S1hg+a39yHOKsWRG8cYkAi4yo1jvEXhxjnoiI/dy
8S8dmgmVDDYRqFUM1ggKUlihj7sZJxItA63kgd6ZppkzIuLzdzs1EclGzkpvdcZH
eVyuU67MMQchbajwL+eZMDYd2nJEcZ8K8a5pP5owuRmovf1MvVCQxAreUzh2gnBF
WpgIfFRgz+eX9cOTNSeKx9pPSTEsOVDpksMYfET/7RZExlWqeyySFglKz/Didpu0
KxCQpGrFnPoGMbr14scliklM8ex0hgIAfOzos5bVkKLCb5KsTvoB9+7OcZqkyiDT
JCGayW5uB7+UnE9FBTARgEQ15ThWKH7iPL73aehd+k3KLZU2X5G+4Pj/7Pw+BTx6
RWzJX5ELVJ4XwH1BLTqUGDQmAsK2rZb20z/qH25+crogrZeebFwRWs+jFJQtc45O
TiO5T3zlPVzQKZO8xjf2SoQD4KxuUCzcA5jzQ+D9knDX9iNu7EV2zeVD8o7BZMf7
KTa0PhAEnrWat3pITcYDQihHOhvzKr7gd4h0IaZj2Wzh0tU7SpcyWesbJ49lHkhB
K+x+CHikhKWzhlzfrKfgELrao5Vp1Z17a22d7r+8O7/kGjXr2y/BPj5DHXPsXxAy
1Cqsvd8YWfu89EJpAOiP+WPHiQ0hM2zQxSS4qzHhQ5AsgwnclHMjiYcwQO6W5ZTA
HWTqnkLTsVc6awvYrTG8uGUe21RZeeDMZBrETk6O8ls1YE07R7RW7SxeEsd4iGjw
ndb12JqoYV1DM3ZKw1kqI1nkbV4/c6/DC6rIIMmvyXvKM+6kajyFKXgaBbMcH2+P
rSQ+vMN5JKOa5aVItFaEX9u7nILTucCNWSG8NxfW++9B5njFaeHqDTTEMtPwUkLO
EdbhY4wyW/u2ZWN5xJtuAA==
`pragma protect end_protected
