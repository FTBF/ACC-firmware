// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:07:01 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ad1AG//JzqqKBcJmeDq+Rh+ikFknMLwdgQqdzxFlf5QQA1NiNFNXO28wn5RC4K2B
csK6fk22oR3zn3MUVgDeKMv8Tqnl7e0avTN8IRUt93op/HNv6EWAfDX+Pp381oBr
MVEzLabV7YxAllGIBuixIoV1FMueg73uRLFouI0Ys7c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32784)
rEIPHWmTIIMYYIK3dqacfrVqJfiaUmt1zTm+VmCSBj9GEmR1+m59yYpLgm4Iw71p
i8g+wUnoqzwBgzIr17eQhv7gSthqh6cqAe1TLzgVkLUhFkPYmm/IVcIqHIqLeuZ6
Wz8+RlILNpmOE5NE4dOkhWMROxilHOrDdZR0vsT6xdgSmRcVa++tbDcxeK6fFXvt
d1+J7voB2KUqcxyY9kY5NIwtGT2WIhv+jt0lxSgj2WgrW5IGQdv0+yTWNcliV2yA
3zNujPxkq+h5BDh1mGf7n0aKXeU/+1QmBeO/lwEqqfk09c9Am9o9Bqi5dRscEd9p
oEuY7svmNNjM509EVW4jCPZ2a3uZ8NW6NGMm8xYH/iAH6EvJV4d741KdSKjPzseE
1ThxxfkDOgW/1J37B/Y6khYPtLfFWjbJXD18D3m2yvY8K6t2XgMIfO/lIyyWYwil
k68ChoWOAyn0tdRbPV/1jzzgTtYHpzzJznFaI2J/oGD7vy5od6zwLrPG7D8EwE9i
CfAK6/kd+PKDXw6u1DJkILF8/auo8KbpDgrA+lA1yHDwWEialz8W2xY7ln3cZjLI
Ax6nGXnTfhxa2Q9XEEUO9b64WA7bJMAmpsORInKBa84z1APoXdfEL7lCRSEiLRJm
opexnwV2XBFgf0H3uZmMYAQ4weOZ8sfp9xlpFEC6E5KYIoI2MMas/Hejx+sZimXX
ykV7bfyHN4/ZSoSOU8pvsJanuSsKlCzZ6S3U3kp5TOTzqauvJZCSj5pHgplvfLiW
M8/azn9LHwe9nF5p1Csh4yqChwWIrOx5C7oZoa+/8KTiqx8W0+O8If4OPu51Nbim
ikBlHRPjcLGJhIIvZoUG7HFXr+vr9NKz9dQ/A/Y4zgeu37+0MMm82nSrcEV5eqEL
Ane8fMfSjvp6ehMEcvpj6mx5SlY3xevOFWJm2Yu32Awkh4kmrmFfxlkBAXsCZZmT
6UvEw0c4g4H2hyGqalbmQ4dk/fw+xGQeMdDaHp/BHrwgE+GQNKNayUnZ4vzGArYQ
D1gEqBnqDWNALK4ykH1H671dTXBjlo/wRk23zxrJ3/sKhO5SmA9D4GDQY0CAcnPJ
AopBRYy76YOU02vcn9ok7BuIuk4mkcVXJY1TAzEeQLpfEDaKCxTVIqeYVc9uGnwr
givO+BK9WBA0INhs3YpvCymaz4hUWMimy/5Fg1iEfIAZnn2KQRr3EzY3LU+EmIzP
xuoC2EqrsqsVyArWIu/Th2l9yJfZDd+iAsO+7k8tf9hjdnvVaY3vQ7KwJOZ9kP7Y
7uc+Ed+tbbV2XHkB6t4v7JQnTrQ8VvVIRycbjtrdwu7uwS3ocaxEuU0LZF30m/OD
7i7ucA6+hwd1AoKdSY5k8X6hkfHbydgq5Y4HnL3HMXHGf60tCEFcYwh38Ten0fHK
6nfV7u5NtYLvj2TGakTy6bSuCVc/zZ4wf7MrIDv/XuyDv24w/wWM1f1EPGQ9JMni
1msqSN63CgPJmriagW00PW+nNf7ljhUa2bEuQYPRAD5VX/KuWbLRt6hU5RUsmvUO
FGMIGrBi87WHbEaa73pXrIPEQkBPZqSkh/5+y9t/993ELVOwHBzFvtupdgdlT1Jy
sWFAd2IEqi2jVGxhR07aE0ueMfxrH5lHPuVI0JpOjB2iZvQWceYqL/apF1sKxSfZ
EhAqKzAkOv9vmW8rQAhsdS34C57pTKfAl29TlkrdYcUoOOBeD1JASyrYRjVVBU5k
FcJPmwCFIwUHvC9IxeeNuV5F6/Y0VYBE08Zjn4Y8sell+7qa8ZFXZ8IwmRVAlo4H
6OJkD/uJFy0XIwUxf+G+PWMmow6xx9Pb9JcAjHYg7ZxzBHwWuMcJHNPXmIhlJ4Z+
B2O0mvuGo6VmGH0iau0eLK2DWyrH0Aqy3GQ7XInrr/6sB7biXSg0XNJHdGqPsD87
ShmrplImyGi+31jXKpS9O/9dCLUyZVkqFuvoNycBIzVY5w5s9UNdwPmcRyTFHcYe
IqdcV6ACbWERBDBrXazz5Od1hAFxwsTQtfacuRq5nxL472iFny4yh/YOkCAYSBQh
2xGDgzFX1JgCWgFXGkO6qBzOE5EFWP7hp7iCrO0X0d0jqzqj3zELwqZL+i/Ksk/u
tdkak9asQOI7wBi8q5r+ixp240/cf0zcSrjHtNPeLpfC5RfPECLd0JYSi85sGDj0
CRynkI3tban1E8AxbnUkuU/5xOwih+IUBLBuKSPOg2R5v6q7CIi6UF3UUp1j4msv
0zR/vHgRJ1mFsgz0Sft6z+Oph3V0jl50Ux9vRryUclYUvskmomAgylp2hi3AWXre
ltPO/RO0X9zPQvgUXAVkQbNtjmVRw2nAtbHIemND/WGjOaPWWo1LxPw9ONpmQUsV
U6p4q+bFMY3WuxDsRRM78lLiTOcgtIhoZCtqPqP3cVdvq76981Uiyb3KZuc+fJHa
UdCo5/CVsvBDuAiasaLw8LfZCetMQjemhYcfo3cEl08lVqrqkhGAYA+yHtHkclln
FOmxSvykrLPLtXVDoEcJMyy9xasekQF7qjRmpSWwKYPwczQIdSXY/uIzL672CrrR
GggP2dtEhELU9OSTbVW+KPAm8GYYVwjib/AUXAtGq2UvnM8UB1KzGiz7tGhK85mg
i0tSIolZL9bINXsn425BIF2ttd2GaUhypr7KiuHeI9nGNn4f2QQ5rB4HCz5FdMXv
V4HorsuS4n1mJJVB2UtzK1QLb/+q3QBDDU3tKsSW6fVqLlf7dwzkYFkjnMVHoCvT
WYN3HPDn7wWI8LU5573i/kv9BpLPGPYCmnmttBTv3p06jMDKPdqx6FbrJaMZxqxl
2rRRPdaUTGzLhCiU0kRVqCZHDpspni1FMYH4tRggGNupGOyGikusZblUtQgotjXF
7MvqOvZRw9plqR5jY/NSS2EymAWEDD2ZcWK2mPbCiwF08H7MBixh0/KP318ghfEl
K2yu6Q2VLxnL9r7uZXJ2iJbPt7DcAk4noiSwyvc+4+J4oLaQoUbmbMJxDZb7s+GI
Z72iOf64qsIL13FeGcc3g1o5SpmoJLHJ+gMwZV6qXwBf2yUc1f2hgcLaiGYLavPQ
kZ2KQ4wrByoGIyoPXZqW5iG3pIuQcMKstdjSP1rg6mHFGexba8zNXzaE9EapVNKr
rCLWfCMzU/9EcQ9JDB4VWDonahZeZovCnsZujFF8QpOa067UjbXIwdNGggY53nyH
eBM9LOSnz3aXG2vNH9Zazk3NGSXvxnhGAvYjCqCt8yeGYgZL4XoflMVh/qssplVB
nRC1lkn+PNYJouyymTUHA+fbrUZI1d2LgQmmj8agWSjn3SuQcHkt1qT/w7Or3S5C
dWUKBquTekf77qCnHWRNi3jPS23Atk+5KL+BSyBIUegDhzIGH1nl0uOzGNak4A9P
KXGr+yvQh+CtQmnG+NnqiAyrou2de9FwJZ0A5m4A/Hmx4yBmB6VR5U3MQv+a0d0K
t3NLJR+ReCN+yZEHxUmd/ApeD2f/tngoJzLGtcMAmNE3pUSnuXozyTos7cf7pL4o
5LUiO/Wxf2pUsMrPGdrFF+tC4CmUiQ0kBH8SHSVPutHRSExmJtDkK/e0lfFl0/Us
BXuK3r60W+SV9DnNBQL8hGxy6iK6/llaAfd0fwfOoblDqBIXjXIHRoOECz6AOeVH
yydb6FWYxfNlu2UIyv01H36iYUSG2z8FaHbNNIJVIxJZxt53YxuljcNMUPQcVvTL
UNoEJOT53zuapA1XuA8iat1l6s+J734NhejsZiWOg8HpG0AoF/PsR6MgpiE0Q78M
8aggK0APL3QYzK2mwkeGK7OVqg8vQOsZD+VlmVLAc+47gcWQNpl/rhTF2V9J9gm5
kSpZVUR3GvhoEDrC3h2AHJMV5Uou/UsZfknfXGDR9X0GRX5sDdKlBN1m/yHm6sb0
tQtK1PYcYU9q6xXkQASgJubPr6qKI0IfT10bZOiA5DpwR5dUjy9IKnZ3MLXuYwvO
z4G9sTCm761zHHhWunzmAXjNVw8XFXOP5sy/7A5o7zE7Lw0Cci7G8IOSvL7F8QpD
X6cHa32yTSZZyZUcYDhBQeDzomEVbZn1+BHXvNxBq27Ugtt9Ov1vpSBH4FZ/C7v6
9bM6y3s7ZR0byW/KwGmbSqGPzwzmaUCiWSLNhiYSjx+TNaeWmMuIeMb1Yocl1tv6
madZEJxPTzJ3DJaneZoR5egdoPhZzQhgbXlmXxvj/UckBCWb5QT+HdA0U2MNeGnt
Kc6AAdSY6Cjkr7XHPeAAUNfNdG2g88UNeK573vAkQQ9pHJgqui2pZIWEKbpi141s
lWOKnzOVRkjTfgDHiHVle2ib1aUqW1Ex3X9CuA6noC7kTnADXkqP7zTs1baqZitS
iZaY7qW/PkpP1F6SSR/HaywA9JoJCtUSRB/PbH/4A8FFZy6D4E1uYfz9CQDtsHBT
vC1P2acIJxROhby8dLvqLkaQ6NuDqxMBJeDPeAFkkI3qc/s9Nf8SKZwMsLW3HeTr
FWXMw+sO53ImUJHeW2N8hLxsTxaBquqJRAbXnYvy6Bdz3l/IKy7cfk+fNBiqhs7H
dbQnRuPJqUEBLxDyG0LmMrDVgaooWbyBJ/Runy80NaqQ/ouvNgGsdclsXbKYPcF2
0lhT2vfpry9TmqKsKmZ+k+SC19pbLAZAv5buvjCgBJ0aoAbUS3pUQOSKvdtZbWgl
2y0yYuPZbHEXRG5CENif7cddRpj5rw9SVmw5mus/ZlkPF51xH5xaVYDoiKbikehg
DHD6sObwkus2sygygRBB4fNEc+o/3wHAWJT6WNDsDc9VjHQVgg2c7IDhaHNAzc9P
K+xNnnOjkKn0dryibBZaHBzOdykNLS3tCgtLW3HL4bD6m3m5EkTBdwfLYYbo4ijC
BoDK5FqjARuRJFNf7aEklWBNxf9/l9k+iRrfLlWWaejNZ+/mkF8O+XpxST4qVtMf
j2p/Vg6i31lZqSrWONG2/PXQokcbW+1YUhFpKWpFbwJXJcIY1NCm2taagiaWqC0d
bHHDWo6A+ty73U0hxYKJI9KmQgQkXbOrZFytbykwjnImtoFl0OXBk13WooV2jYrp
ZiJ31roCGN4C/9mnaHMhleBzFw0F1JLFV7Obvl+wxoLcJKwjkL4rLL+BLLMlEkYh
oxUbTHf9v8KCtxyx88y1hgN5l9e66stflN3oX5aSVi4Ex5bYxfSlOrj9VFd9tmhZ
EAiVEW8DFS6B80W0aMDFYIXxcWlfrRN2Up1n5iRUBO0wIg4jqXhLDWuYC1bAiiVw
IDJ+Bjw+7BOdRBVT0FT7KufEGklW//VZX+1U/q+kvlKf0CGVjJpW9waTFEyMaRUZ
GEzlbMZjEkvaegH1zzNEJZ6FRHjYP7O2JEhASS0qvdPkJthFSfU9eYdhLGV52X2Q
cFmuDUKFHihATtAPKbj8MZFdTR0LiBq8Xb3EaX9cuMZ+jyh26bgXnSHcpTKLEe77
3PqIZ8HvMcM3o2XdwhfbbrCpiKQaUYYRsLxK+rIo7zvLxcCjrYcD0eYxKlUs/tXK
c6c2hJR3F1bPitMYv37em7BanUdOiF/IuZ1LpK8AuyReU4kW3IV3rbGssKTUPcsD
s8aXgq4I7BiVt2vSA27Y+4ZgzgJF9Vq8xDLUEr8ENnSk31AANR+9ic0OgN5OqKJ1
c1YBo8cd4+OloWYFZI2M8sod8+/SXdx604pwbz/mwpeROZ1CqaRzfPXC37NMAzUc
63NuzJKvaGPMe5srffueZOWySV1HwFZWleiSTc4kCd6soilOBK2RUnUUIOO1G1sE
4c87TM+3jcjMuqTd7LgdR+Epz21lT5D+OwiENu0cx/An26Lj2kHbBQfqxgMmqp6J
Md+xvlIzQNJ9qCttd043g7y0SfSpNg7CiBAlkZ4mXbUv8yLeDepLFNYoEfFVYaay
ezFHenyr+E8nE3qCtUslOSWNNNVGr5OXfCZEJml7Df6evOkY2G39Z80UbuPUXdst
msJo0+yJcxA9+6bwnDYFjk7+lFjdp5UfIdIyOaLKYi4d8SFV8k48YAYK/8L3ITjJ
t0EN4oQdlPpc9gfeHgtGS/TQoSo/eckRE+pSxRG6B3ZfjIwFVGCXMFTzGky8U0FY
/F4CTcrWROXb5ckZJo3lObglm/WQZUS0Z8ZlpnJX8QyJSP+LCATRNt9saWMGpjrG
Bdt60jIQCiU5b26uuzlAycoGtXgvexSz1hhkQyWkGJbaf4eIYcA5BtxZPwesti4c
+hOkcyLvOya++ZoxMUCj1SZgaiKIxcvWz5sei2cxgbsXK19mz+jwoOIpgxijxP5+
Co8fmb6zXmQo9ij3YTHdZE8oZLNRFZPn69TqOpJczpZXXexKScqlJ0vXSC+As2By
FuMxWGA0uFS61TP+Yk/Xamzd/CATVoCJp4W7DUssREXrc19dVdhaA0vekyp90krj
cXM8ViroPYukZTtImVGr+yrCt5/WzxOcaFPaHSB7tuK1YOHzWxG8uhahfqAiYWNM
9xepr5JGIBjL480Cz4noi1V1JzHykoBjzQJGXS3WEM7lxAaQ7IPfYMwStQsGWjjX
bdbB7v/TkiWkMDZOAR8dZe81Wks445dB/N/RKW7l4HRgUjb0wlih+wDHdmL73PRa
Gg2ARJlilIYHt9SQF5jv83X6b5RTIz1dw/bC8Z+g4vLWQo+0UgJ23t3322Vf1dNz
8RafooND/xDZCMNACY+Ykkp1LXxEOlzjANLYmNbkoepWkAyWaq1AjGHD84JYwpgz
qeKp5eCdvQ6l6lV1gog4jhwcGjZJ2OsfrojcC+pFkpkQFu6VQrQS26y4C/C3XO53
A8aFAA+UqDONUEG7FyM4zBeWfvKwc5En3UeCuyYs3ywBTfPo4mQASc6q66JppbRW
csAhXJylp6EIy7nO8qjx5sI6a+Aw4y0+/noFZ5b+Zgb/zzhYU3NKdvtioWPMxEg5
+Qg6fAvaq7rmDQ7TfeHtsySwvIRIAqxP/cgqYuFw9/bsFfrUiSaZyo5NBXDRNQrp
/wbTroaBa0zzAs+hX5fuLvfM6MNYbPk8I+IXA/wFB0MUGLwXjk6qii39440jvpqH
/ZTHD9pP6/IIKtPYjy7D4LmIilke7WiRLBmCvDEkUe5uhQZJ7S/U4i1vRhMQmkYz
w5653qLiEU2BgxOYlA9gM/oIirZ9JivdpZBwfZZxbw+BMUsegnsnff8DqAw71ZQ7
IfDaQCcc2gvyxU5PRmCr17anpRo+WRiuYlHbJxHAoq0vMV5zcZYT28ukglPXO3Ma
9kLNF9oZaukwbQzE3xmJskWy528WuAie9WDKP9m15RWnce6Us9Gd8Ra9G4pJQnM9
FaDrwgkj8v0NHlyOZBypmZsVaUTVhQQRjuSANHdVVNVOIkYfkzHn+llhhOFIJHGl
2LnTw7p4MR+7Ft8QtZk8ouYv4lioBpIWMPUvHo7HTMEQHERWRBZqBPu0kG4vaZJ7
de1yJGvCCg36qZ5ISNP0vVkb26srNKxf43ODWb1UnFMgNMV+t8zS9mjnCCuKG/yW
yayFT1vhJEkV72YTIlOWpzCbQcql1cKl6sd3YjWVbJOSzWDncZMBjifBcPgflq6z
6zSXO3kI53IHWzlrNSsuS+BMznGkw8W+Uz0DQgi+D3WMQpLQ7HqvVqYTgag3e35G
Daq4RVYV+fm/jWha3BK7GsvXcgWXDItJ/pYyLyTdc9fUoPqZQ9ED6n8PXnYdeNJt
+ZWM4h7O0Au5EhlkIRi7Gg2a/I0eMbMM/v5MF6bCVnrQ/aOYKFXIq87JU8QBTkr5
8hJU2gMYpZFcWLwOwhWdXiTPDn35Awg90kOZfl1MQP8UwQ44LH4qVSZXLNDsr12e
oa99zyBlLea5aSB2l6cpr0v5Tr/+CBGDyOlsqPEpuFXiZaaD1WFACRB8CRcz+1Gz
Pr7vxbbq1AsTeRUYfZV13gcnYFEmVL7n3PPNeYArl0+HxbfzQWA3/WPkLnRQCz2Q
gRFJR95QBhmqFrCNq1hGZiBsLCLfFkSgvSgNybqhuyNGQoCGPJ593nusmEid+gAx
emWBjQ/kRrRrxwbA7B9wz0n7HmneqV5MeLQ3mP0RbqtNIbLdTApw2zaHhdIEiU++
G+6KpC/Xb/KPzy1ctPfcmfxIYiDrseDPdJWXRftZ3LVmkY7h9r485TGI81Wv67oI
gwvmKSupXEJqT1R5aFzoTNM1REQf2VJJZ4jy3UJCKhZmmDjGH/rVQYwDVe9EWQGS
1qDTFHJp+thsbuP6qHVOFI9rbWEF8mDwXaF6EglkVg77O2smWgrezgFMoTauQKEa
Eba2EiBXTVZh6H0RWEK3miTExOUH135un3q/1QI5qfMnDkoj2OtmEiqflUps3tCb
XPOgM4N4CkO2WeyWXEPfa0EM0UhNEyOvEf55LK75IsRqlQyFk59WEF2w5NFxishA
Unim2S/9NZsp2IYzaRy+L4ujxyedwCaTkpbkuY/+aGKCW6CGNv9zWMH3Quy3XxvR
vDJTtCjHpHEr2xkxybP3OoVNSZAeAsI3Ux/jPN/O+2x5QxjnlS3JHZhH7kRcyRSl
C4EMi8kZscl6ruiyDuj42g1jzLc9z3cQIlJ9Co2n+D/QFXbxbSQUIOWcZ0eW64PN
+tm3nwtuNl3knAJENzeOcD5t1+BlUGWP1yzGobSeYr2+NPbb4mezyX3n0CMVRDuF
ut2ZevmFvuhN9GW6BOIZ+QzMByRDnMk9KRxorqpdz4iEn0LK2OO5NAdFql5pA1TR
RUfBHSe9ypl46abWIKuL69xMC7mcd8jmh1R2Bgt+d1ZgdObkBuky8neMqT5Aws5B
rS8UNIzoPWfHWqO1C5pLHF2cX2adj+resq0sOyLhxKAhMmpFnFd09ARDDEWZbsEG
1vgLWDzVvFCwftKIApsdlHA5AX7SSmxaTdvUIhpEFTGdTpyIluvYdvRY/UJW5Dkr
qz1Jn/9JmtYl6RNoHoAiHS3FU91TdiKjlAMMqfKVTad9yfRGJOT0rBZ9ShMR5ZYR
piNIQH6VNawxJxy+/SbEDQhTDMZPwHMPihnluAfFanWb9bzrfeQ9FcIXKo5ptrzU
J+ldF1MkPoQzB7PtUvCXQXTzw6dun/vDXc6s/JXTPzwuoy/YSE9EOB8Hmlsn1HF1
2A/9wddshlKynx05xf/9K9qvnLNC3xRj/iqQMStbCXGMoFxBILgSVL/QwENzWIE8
wsuKXsKpdHYcfV/uX/XmBJcvEBgXaetDwdLaYvjHuN6IqBBvyAgtmBm9MSgui4pn
/IMe8wMe9Q3JQsVNr0rJjjfltOl1v8MJdIBP0qDG7mVHbnCBU+WC0UTEHjSfNgHv
Sm4ZB3d3yUlFvD+V1z8jK4KhPrnCXmKTvYfyM91lhG7PNk1nRzHn72M10FcnIVEx
tSXHuwiUGVYkuSNnKoEz7VAvkT+BN1ivsMU5KntGGMujlTVAL3ZWTdMbrb+KaKO+
+zz5MysFUVQHN1CA05qbrJ+8WNjIQQl2wfIiC/ATjvsklpbdYqrlbL5Nc2zy7Ohq
7khDlaJBd2ctqxiw3gt4jhANiWq4/xi42jIOhwxEHmsWyS8VzWKkbNtAuYnbjQvr
k0NoUihsgrqxxqqsSXPYtVjcaeWEACMWvhozMrPfVVI9h6SVF93qOz6V4hVF0P5d
7n8AIvzPL9rwzuJvOj4ALR7QEVhK887aJsGGpfTVUQExPp9P5ZFVKmL60RDJslZN
m/Pf6RUmOC4e3odPTagY+sq1JBNltghBvyqWaezDPRPxa9QzfE5El2AtXu8nWmSI
8Z6LOPcGu0CDowD5QlMvggetVj40ysg9PSgSPw3CQoo5S3A8iUuMiGjr07hAL5X/
6lcxkJ/TdbVucSx2SWNmsOoXBgR4wy2Qu+PSdCGHSwxVxXXStyQZJEXHxTcgmtOS
TFaSLEae+DJhZsMVoqCKBXgNgE4iOIQUSPky7l8kygOH9bQZK66mCMx8RMV+BGna
97z6Et/+ThpXWbPpnh07++m3sf3RY9UJYtZR+xkZI/A7EOF8xTJGxale3pxcZ/OV
OUos+CvxtPz4745LUQQgFa4naSB7RE8xFRyGM6JUcXCV0oZ3wpdxhft8dt1IRzTk
NREA14vxrimbq0aYBZdA7JdYoI5rU3zKEmfIHWDCZV6Ft8nLxL24Qj41n3W4biKc
YR1whh8zPBYA5FloWQCfrfRoYYeFJc0dB3O5nbFbIAN7L8bHowPOfkTXU1QmTfmz
LycV3cx6pehEMT77FQsQIyh+prwr9AdWMZAa2VxhuK47pnEqe6IZ7HRWDWlObkXt
3n3ZN0/cKWdzfQKNLKYZOEaQr9K1rG5jfX1OdUckXoKa/KZ+1Ap3XOmF7zxieM4F
7WAcISpHAcOM/fAfh2Y05XpymCz0QWPP89VIbC+nP9a1ZiGzWOzuctNKrPEqAmUD
rh8K3UO+43Xw0RrNiwzYfkr0d0j34IkGUrEWMetL1LIUi+Y4d6OrIiAWhDHMxpuq
wW81fDFOZoYIxVGGN7ld7cQqiu38NgkWSMWFNMKnnLdSWUggZPdNWT08/27nHM8d
8UpbxUXf6DLcxWl4fNGUzkKtSJ3FOh8zRzzIyAU2qUM+A9VLJCOgWJnkMFEPg9mK
egNybdZ+j3jrOGAZGkhUYm4rs2jsddej0lqZCI13iLh7KgsnLKf0vlVc7NgKVkD3
Qzw7/uUkBomc+W1Y4+MNcs8Cl1xbhdJEb2qRzMT6lQ6ikHTflDYjoREl+Ei4RD5g
8z52T6NnPbA9JoDohOfK6w31nt4rzBpfldIrYtNem4PauyTkaeRCJgbxeFhARArQ
oESD5m9PALZufmHqwpQG69wmOuovQfYvmnxNFnBI/yv1YEP7NrjbSjvdFVWf35jb
Zbaetg1cEHIaIKhz0WSsIkfL6O2Y+BR8XE1Ut+AvDpzvkoAzfIcX0ETAzX8S4Nts
qjDQHhYC6WPRcEyggf9XCup2wahngP7baFYLpb2JPnY9T4MNHRJJL3rSMK0B5ZXd
viF3nrEAaNZ8pRQJrcJxGpMJFU95ZxucHxVlhb4jtwNSsBuxA8ccoZVFHtdgxoHC
tkoPBujfjOxVHih07VwaeHVGVyUBXEeJDy9adw3zFx29Fmpd5B/9Fp/NReIQ+amn
ayjvjL/c09gZx1yDx2y4t3B0rBDO3HIRMA48frVm+9q8lyJoPI+AGogkvSFoOkkL
vrxLrC0oeq5rqQYLO4rLyh7hy3NPEtGyGkXEnBhCWIaF/L8kngFUXKswawU+oWLY
neVApCOyduKjB8/hoeGjRx1JVPpdUCBEf1gm4dCa1uQ5ORyZXG17QWNLIECyt23c
jRBxqjCrUDf8sZosAW1CqRObvvHAJy9vatrtpNrHNagpozuI4RS0xS2EW/Avp9+b
R2942ofPuuPaB3NfFgNPe/96memxYPeMfBuzMLml6hJuTy6j369KeHJ/JlyDWA4W
OIhZ4dpKSoOUKRsL7Axix5nEr59cUDzGNIegD8EbBT55dSc35TKz14S9ReyOzXL0
UEPqfV9PVGIR+jme3hNPNiXTwgqytwcpKANRjASz8cAGFyD7JPjbYfbuIOFbLw9h
haEkDsUGfSJl9bDOjGGhE2/B7v52bwSj0JmYb8BAMKs8q6imBKsCA67tZtG3W/Gi
13NK+WB8PjEy40yqEUOaIO9YoBKJpRXAtGfqwXpDOwgimQVgUct9LhNsQQSJeNLz
CsHb0bjunw/vXrdkN1M3S2dnCNo5awx0Fnp8qONjXJ8SuFO9KdDu/v+I8gW2W9XQ
phUxAscLIJnzPpy3kk+xCArwkziZ1/6r/L8t+7r92/02vGJqbsL44/0BSMtKeQpo
CY9FzznqCLbMjkDSwLo6Yy5eClYoRt1r+S6MR4EtLPb6/FaDEIX8/RpfDMBnfA7A
QdN1bzMfgLtYKfU8jj9uC/aPeczDdKheQrI8w8M7HXpgc3Cx82JQFFtKmip2OH5T
CbvOVnB3ecUJw8GJwub1b1GD1HBqDA8NAnM7GF2uMcPgBHWUssM1jWMg9e1irz7B
r5eUNnGmXELfNZQveRNq36/G5CDyKDrerP3NdmxzGUeCjzgvDO1OASel5iGSi8Jt
eT5OoNoOa8CVppCYag65rLFz/npcmHEUpiSn3G4lmYt3mNYpwfGrWhqSyOvvqcBL
v+MhaSixhBlJuTVvvtlkpMMfH0DQS/cNcB3p0oLQDQi5VYMwmQOcYgFw4EmlgO2V
G5jdnu+N6IfbeEwxg3AEeIGVxjKAwSONuJ51xOfPHFXGaYHShCZH6e+AwdvbUhdD
R784NWDd1eiVxH2YxZYWltzAZyL8KDowMel9sytjygyW0Lx8Wn7Wf7i3YDf7qwFC
rwTh8RCcAoVBG2Zyt7XtqrKkAQIvO44f/oUkxZyIGjUwxvNshbF5zlzvLeqJHmDX
hiVlUhuz2zlO+CLFxTp04mlLQN8YuxX279f2dzQHn7QKLR3Ox6gOMBoFDp9CA6MC
1LYcm0nI+2oE0Ts9wWLEHKDBh0N/AGnFwmcWBuGZciu9unD3tLE7icziLAGx9CiX
siCwGfcx98wyOIsrclGsLcMUs6c7/WnP+Vy26V5T0bxobjvyDZ8wrFFh1jpSdn7F
O+1rjfOI6xrFKdooxB1qdG6qVjXKuz3q8EIJ5ckWuStbCyP6GLPt2u8DnQdY3Ve2
aEUhzCmkho6wqzA4kmSxAlPb74v4wTpDPXJaQxJnfiwZ8bTapFqCBurntNZid2MU
FHbAnFH4Vr2W1hlzaN5+mkqiCPZraR0TQXHkym5NgdpjFQ8O8+AXUzhnB7kgAZLC
7ca2cg56vVREBrVmXOcwLUucNwGzJE3pUw0H9GLmEkJbtSE2qLo/KaRmhp3wn1IV
kj3zZgszqk8nlAu+ZFkgOTjc9uBTkZTL19jAzixvmgM5nfFdAGM9HicxPV2t18Qf
laKmC1lm69lr+maOGjtoNWGLJ6IuafA605DGjDWPo1MhyPYoIWtyGvPuJ/nwOs+c
gASoXz9Vn/nYkg+v12zURYB4U9+9iapXfeif9j1S3Eu5g1ZAmIL6bipEdkXeDfb2
eGOAFyhatbG0HL2aSp1DYxQhZovM4w8UMUl2MQ1LJmcgja1+JiOUQIt8XkjKrGBe
BYKZXiZbZtoFV3ZpEbTqBFpW0SIyzXdUF8woCy9OugvnppMdQjVb8XgMlEr7EigD
HnnpJg0UnVhwc7XUfU2+0gs/buAOagujsInmrMFOgsTEP9Q8PmhSLI2KyplLqHqp
jpSG932DRzkVRUiqJeZZa8GE3gKNvfsSgQK0PNnfnytJ93hERKK8qvc1zcDxJEyc
UJOGixYMU+lfOI7Uu97nkxi5ZF6ijfW5fWtceAfjCbpP8KvLpp2OsYFyPeYmXsc6
dgJc8n0+IzEknu3w/UzJOPvtaTm/YHJo9HddsfqH4pSoJUfJU7pnTIZqF5si8Jm1
qSHSYjmcGRYS9uyq0Aznu5z7lBeyBGHVbJ5xHhAyrDusrCBRiKLNagH/q5Ax5y6b
I45FM947hful/IZka/VXyqG56CIYlzh+LqDZzCjeh2VmMGRYRssY7P+1nn4BKVZi
xTXQUj9GWwEhWP8M83ox5Fa3ipRo1WeHT5Ts2di8Wn9yyjd515PcHlN60VCT8L48
6/deQ13xjjEKpkHd1hMjIbg9efNVCyCLj0OWZ1sE3BfU673hQ6009zmE18fYISvE
V77Lon3S/OoerEQBIJRME7wpAviEhRfAqKQD4PZhPtPSnptMf6x6SpqFnAudat3E
KSkMnvUofPUq7M4cKMeIY99NdLJJMerM5cad8pyzCRzA8JOsqrUoOhaueVzWdzd8
umrupNPLekfGbhadPU4EPyrV8Kz5nMX+dZS/+QMY6L0451OiOOxBXzKp0BStcZxF
ppR4lMfUH0lR5hQBF85i0ny6KbIPj1MvEOd13Gjb80bkH8+0aSjP8DBJcr8+beju
EAbdNiqb+X78TbHCETzsB4FXsLtYyPJV0x+aZr2+zd25F2Y+7GeaE/sYW5KeClE4
vDlHRj3nFlQzxEfqwaiJ5wdH3fNfgABHgFpc/oBEmcTeBTyv0al75Hqv1ka6RbA8
do7/2OMCKXV89QsS5Vl4n1X2wQTpGcm3U9c0XgH6E9RtqecazA4AAgEsHLIChwlD
EJdR1t8uXI1hzIGJemqgLt1TOmfgiTQ/5hIMWps1H6OeA+U4RDRPlcnV+yw/dUuX
nSdai+7Kq9YFmDrOmJCOAPo1jXTiHc7HZ9UTPN2QSilbcI6BrlkVGQvMY0JWWZDb
wI3OD3g77FCE0f+W90VUWS1dVKRb23kX9YZGTcPH8NOLW5rpy8W/N/wUb3udWamg
QDmDPdc9EIKk09FUI1Aye8i9p8RMln7+EpCA04DV3+7TbUR6ccV/o8vMKA5liS9c
L3wocnvQMTmXymZNfTgZzeXUR/k+yWl+dXDE+0qCKLe8bW4dLUaxM/jBtSipzpHw
GK122kQ9+9x7qfK48kCicd+GbX8ka4IxgjOg0/pwzYMutbb1tX8JNeuqbOV51PhT
uXronorxS3cBChZhPjq3oQY0ops/X5Vs/Pp/bg43GPVl8AaMiu8y5bGIdThU0cX6
sxnE1SCcIgv3aUSDk8VrjhUR9K5jNkSviI85HwNY3kAwoW4LZyzluhsIjDfJiy7s
S//IBUOmByzv4Y/jmznmdbrlNzfiq8fbBul4mTXU8lNyj8MGlqdPEc8Xm3vNB5sC
XuVziKkqK6iFUekIxL+XRkna4CtUuKJCV00LAgLs9fxVcSOALtoCee8U/03R1lZ1
k6/uzo6KlZwC4IrcUjdA97zFuFckeP1SjRPFMXXGuzXZ2IfoLbGwry5TGvhGSJi9
nw4FanaOZwKSaQrWnMXIvPx6iwppLPVIkWp6LSoLbmuc8hxo900/XE+6wXBoR9Of
YQMXH9UI+naqfatnB41tW1ZunDtpkVyqnWhm8uh1m9P033lNeYyngFlkUJbIFcpY
mVby29sAihKoV9Yz477oEzc9PhVkULOWizwl85L5b/bM7KB8zdmqGiXZP8jRNw8B
oB9L885oVK0EIP8z9OWySDUI9AsRY8m35uXd5jAeRmS9N2plAM8+uvgOuMaEmH3Q
8ZJRolXZDwwkf6wta96Do9V9FOvkZvhQ307QOA8UPTE3MoJ2JgTyTWsM8hCDur9D
KLByVlCP7JHeq5f57gqvT/AWrOCCZtLRMmHvFZm4iFaUgxhWw4duqzkt33FMZWCL
SbRxVl1CMwmJFDqYduaacmok3seDVCzma6cDd5HQQ3vfkulM5BnF5dhX2lzzo4sM
Es7dHXvUl4G4lLQiFFvNy/6/6AlEkGBQHnTeYtvSuQcjy+8NHhuEQT8fmeAgt80t
4MF1uMG2lOr3ONd64VuMTc+vIMc8GAMiREUYGK95s/1um4+AgyaUcDHBrbO8dzeC
xWUt6BtJS4b+GK4liZfCZIM2BirbBaeJ7/GwVu2jgysGKjzr8+v702RSc56IFXUE
f3SmNvzjUKSwNiOhOI2r6pciq7eKyZpEqdBvQiNfd96R8BA61uLE2U0LQk2hNuby
SO2xD1WwITF61s6uwXNEmcKOkpeQd1Dr8gBoe/ouHFlZjHUzvuyEfD/4hHCv8wvq
Vkxu3QR+izGrSmWnMVZ+sZN00izP30zrhnmmLRjoouo85dYEPR2KbdhlLA3TBWKT
naO1eRY7kCtzO1jq2yLpgws2GE3UDq1pK1sTYjbRqjPENx2GfktFk7PIhAK5mYHo
HPixEINyZu39CIM4FfYdUXU3f2xZi2Ki0Bd8qn7i9DMCWqQQCtPo3p6To5P2EDkN
pQgbfUlIr2994k+Ay+SEb538GXsQRrX/C7nHCRd++G5iCClpF49mQLL0VwCGi//4
bxUcb8gro2xIFHHEuPh/1It3z1v/TIyzw/bsFaFQpaZNc3eul1nMIjGT14G9vMSL
IhTSCmh5qQpS6nJbNS5RT/90YdesRKhl1X6yiDKAkf4fxMxChYwLESf9t4aFC/8G
SCTBoOzuDnqylhWY9ka9tchn25BIPEpxTljWYLqBlGfgl0nGWdrLEMpwQsxehinn
CJCfBP45lcHCL6jQRVOt4nobhzx/9is1dVkAxUzKUEymhclzyixCwabCIj5hzNss
hr7UGrIzo9B7m/cd6bl9pvubOJTFhHlqZGan5TilIdX+xOhm0ZUfWzUOzydS1V4g
ZogUkwIiHJI5gKxEY1I5TboJJoZZgbmVYgPOBI2vA24Ia8sUWL4Z0VpHGiHYckVy
DGMmrL3DXObTDknxblzt4ArzTvJt1jdJl1a1Z9977+Fjqc3DFP1DRxt0xA/uaySB
mopL4+X39QZj7ur9d6uTf9Uxb3mcPM+hQ0zEf27sYWpVgK61vJbKX5weUeBczuDQ
Ew7t+pNNbpeekZn96Yq44zKPQ9vXDSc/NMW6AVMKQSWWQllGP/3O4aYtyst+9/i0
7s/6WISb1eT8srBeJ+K05K030M+GMA0PxBZKevEsaxMHCIV8+jmbF11j0Z24gZu1
EQnY/s0j0ZVHKIS/94I2t40oJJhfDqXzRyHruDEx345Dxc8Opc+2PSRR2c3wb+bX
I1ARRYQUH14JkWVFhozG16JK7aaEylgQ2D/U+VshXFuBDwQps/L217M92XFgqLBL
dv9JPJj+YmoOwfq0VVfEVWbzihCmiSlorJm0Y7Su8acWj4hetj0X4p9/NV6fVP7B
af0fhvWdwYcEBfmyyjXHwhgvtGGCRzFNqWZWaVEJihvxZ/V5AU4+CG/5gZJkHt/W
EbLfqwUE0qG5lyC2Rf5fi9UMNccPGxzbHBId6DLtacxznrZB583mhnAq1JumjMsL
Z7A8nDEnnGdZsmAi74B+3ePtiQuuY9T5Iu91+Y99OkM2TBeKOUORpBq8tLJ1e6Kn
gSAO0dhWKQ2ot8xJ5W7YGDJRqEqZpciMPTfEHadpLOyGwwtd0MPmUElzUfx7JvHw
SoK7sKJBxKCwk0V8dciJOa6FUtqnpYDtMiKqDT8r8q19mPgIqS/HCXQO/Isf3j2G
JHY44/cOwiLm/EYqizzz6NJdmam+h06QT/qUt9r2zVsGxcBj/Kk5YI8zKGL0bcMq
jamRckrObhd0DcijcIPhUHURSekBHLFcSTiY0rcxismQiR3Vvhpeq2M03cdPoDbo
Huu2LnkW8igh0ZBcmK/wZ8fxV3ePrNCO9WFibOiD96ZELSj4/bYDg+HzM4hGFENw
bi1gXZYP92R1CWR4QikyzWNeAF4ptOLEhqgbrEQieL8Uh493Qgz7htA+wbrocaNN
uROZ1aNH2Gb4bV9rEgTKuHo0buZRKtRJwBch/bNOanPso9G6ZW/6AAlCf01Xv+Wa
9LAP74GkRWUquFIxmPiTzakqS76GjHPN5sjW7Kh8/gPP5/Emw1lMJzztoyh4ayE/
JPI70NOY3rtv8TUkfIRChEOpat46Sd3ctBW7TusFRCZ1UAxZecS/bwMSHyI0bev1
CSl4EJEHskh57gkEQzAVU9ds5JpmwcugNB0nVI0At2CsAFVjMuL8vwT+0R1DiaKX
aT7bJf0pC7GnLJWNCYZSZQ+LeXHvCVCLvBIZegzeWIXMchMaZpjzbsC4uvXCncdZ
v/mfYiHDuCmRIFk38pniHUmPYB7YZ3v5CzUvyJktHrRzk100HwFTtIMLYatIItEE
7T4mEcoiQCyNfe+nR7bz0vu5WcouUkhJCxLJlSe36QNx3p0R/NQw+N8+0cIbvKPQ
rCjEfE/fc7mB0Dj0pRai8hYw+v9Sf4gm+3VOaEy5zYDavwvQd4n+PcK8vzIbZHjR
tvAN1jlwvN87VL1Covaw7wFWcHyVowrl48eX8Vax/2wzAN8vybEuBEDFyPq8RDZJ
3LgvhPQnZWVzfMDxhzmBNqHVyQ60Ewicj5mjeRAElHd/Kwy9W2xojlhvw7C67RoB
HlIG/9rKkNm1QuSfEMtEiSTfUiy6wDxkbiLhOGOn0rQDiD9sZcD8ZoOQBW/Un6aI
wbyzr3WDiS5kCB13scEEu5YsN6REo2gQ2Q9dAd3GBH536O51N8eHbx1rYK/rT04M
O+qFkQVhjUdhpMe1/qQOQ2Jb1cqo//UCMANqy5rPEhzL/hwVTF9A6Zm85Ly6aqOA
oG2+AdedCqHg6mHUI7c3kHh8skiTZIVOQ4ZogrkzihSz8XDvhdN5gkhs+QB1TL4L
aZyaVktt6QeL30+GU8+Y5naUBxA1vxQwUp3pZdcrKwwGvfkeheCUq+ax/ALMaFPz
jpw0X9jBsctmCMHnUhNZMPCz0p5niQSD+KkdZTw01ycs8uOr4Qy3UloCWH8j+0RI
rHBetwllmswWzcXWfRnzV6zvqGvxbhoi64tl8uU5h0IHeF6YNe2FbfrcZ6WIK8WV
0LBl4lxxWfzYXby/Atxe1hmDTD4tGAXZ4n3hTvAhFyKvZxsbedHlGxAAvGZlw557
XPD10WGd6Dkq5wfhBS1gcvk2gHNTr8jdClHOSxymBij2GT57Pl8kDlkdoc2CQbJ/
doSIg5gCOkZcPY0xyjntzU9QUkbhfJDU3J2ZLt4ldtQZbOrAbJXSUqHM7oyWMadM
cG5fhLtEUcnacUOsyR5ubQUlJUgHov1XUN+KOmtJwXK/aFwUPN7zdwmAXxw1ceBE
L939QAeT2vDZihnxnUDOkX+6kFkjZhXbB91j5x1DpzwvADDb+uhpqlyuwgTUC4Yj
25lm1ZNfcB3exgwuvsEMrjbgf4T6DeTzejgGY++mHZ7Pj3gJOPqO9yG4aiqbi55a
3pl7uvd8ZLSG3OSY4TI+K7hgRQSazC+D3ajPFmgk9X1DrxDUvTjpCIUy4hFf1UXx
wacG8okysXb9o56aYINlccC0je1/p1LCWvZOkpDYk0vqr+lgRQX2lX+vBdZ62DGa
P7PX/7T4ypQq98kzqAk7uVcfEGL5PhmLL0fCWlwn1zJfZEMk0cKxpvsae2Lo6Emj
nJ6NGyOc+dn5CV0/5lLfTayqS6uW0SjW51toRWm5uuPCgUHWeb2T5343vZhMM5RE
aFfzMwUd80mrSHj7hjxVwVFSppT6+yfi6kVf9lTA8SlEq4GW6IzwP7T3nIw+58W2
wH9PFp19wfo5z/TowDGu9cn5hJPztb2CU1a58qxJUVLx6PbnH3/tBvqcbz3pxUS1
TY58U+eaDXIWRLx3VOGBs0m5IqiJ3VUJ+n0MbwnUzrpYlxuFE8OFFU5uxIzdy2Rm
TgKMI5vD8bkLDcdFpE/1SjUWxwbHYqkpAyoF8g6Eum01zCcAZYmoMHRm3G1E4qZu
HSXLdg6WlL0ZvblBJ26GIL+dcYxTykdLNEwxsc8MG9mWA5EP5v0pLINSmgP/7APJ
XGJANxrzYH9Uvi/UOuj+yLvdWpB2c6mAd4ek8voNVgK7ZS4YSxuAnGppVNajYCEC
m1C5IJup1D/zAaF9XcT61Z+J9Iig606RW8v+/7X0mN3Zs5KjhHEIW3uVPdP07vS+
lssS7oHl7HgSuFtfUlIvzKaX6CS6Pl6aj6aEidWLcg05k8rvVcD5dI6QqRBWVCC+
M1XAltadHwa5im8okN4DQjJ9N/3WzTIJApT5DPCzUwViaTsH6uKcQUhHZI4YhWPl
ijqvX2tsOHOyMd+3Gp8QAKJDgXTeSpU+vJPjKc2NxLWpVRrFqmOTYlGDqwIOfoX2
iGtdkRNuTsZGtD02uagAZdRoboZkbtYqU1E5QNhoTxZkyqErikyZ8hQpqbL4+W5s
mpsJIiALIq4HPL371c94IpLP5IuycYKH79GNbAZqGWtKkkS2g4PGYJ4JdZk/mYVZ
qEjK4Dj3pLE0bfTLvzNk1myrs6OKg0jFTq/OeowEBoq5EshgOxMf3T409LbKB4Vb
1zG/+zevZntvjqKJo1kXvgHjPnF+9KmA3YoW0g7zsWHYehNP72oBpGgE1xgFtuFR
uM4OATZFV47Kqq12LJ1GBsb73ZmrAa3kB8c079hQEy2j88jeiZ7UkQXtcWJrEQbt
Ggg266uBVtT2f659s5imZVh3zUjSVum0V9pVgHS3oig3v0IKIhn57swvm6J3z1L0
QaQwiXENv/gQVY6zn3rLguKKRr+emZD1hEIlHgDPtHTSv0lLcKzidetMvlPa3GJf
hDCw+dM1vpVp7JxyeTbWEJxy4zte6T1bW4gSGO8BOWF8C25Rv1TGADWKMrgO9div
8kH5Uq7a5eSIHAwxnhmx22jXWpTlu2noflwx5620AMeF+q+FAUnwA0cMspPDZdNr
HhEnNR8tDktLt5Icgr8phomPc6LNZ/1y55TEVSQKNDuPyzcTum4FUjdsEjyPUpUB
IeD8qxb/ESb/LCbdN7Sn3wdzYq6zMqzPLTNRa8M6SHwhcDWQ5hVSikwzj3zEMZ4/
1krw7KO1XmJ+G3pcMBJh65NfoOZI4PdFB2o0qFeN/izED9JseagRS6ILWm2WRsQD
9eFRAqims1kvIOAdOfclt+L3Tu7ieOts4/RSa4F85LKGeH9mGZ5zksFNaUPrIySI
0G0JhM273jf5wuXeqMULVy6ovktsd+Q7P6KW04kNEZ0Do36ZwUAgXcmg1EoPQf1I
bw6PyNPhgor2akgZoU1amuitmITCsXhpqAuARNIlx4uhXyO8MA7/NI3O1ABNGuGh
samOjrBkuQ9SkJw+XjXzWnGC81CkcLwqqteZGK+Xngaqzk1may6OQkI7SD9axTsB
2d8rEwWBR/znp19CB6/dJCOiIQQC/XKL4vQleX7iIYCeOL2yrUqa/4RA6sfcYp51
9cbvUGpHwhBDnadBkU6icNsRoVLfGjbHVRNLD2Mx3fRzhVB9VwUkGnYpzWoUmeAG
6tEwYdhiysK6AadItASbIphCD1KJ6hvMsUoJcOkRpZSYmpEGvsNCg+D68lQ3pxHj
4t10ZHLQ9LUioblwuiej7l3enewTIVg0EP1pufRfku7+X+NgGuyob2/vHsb5YlMS
AMKlahRWvWesF4r6dt6e/UZuANbOpABVIUFD0DT2CUTi/1tB2z6kn6WVZBIunLu4
lWh3kZrjTsZ6MCtnZ0t0+6lPIUPZ4V0DXatABrvekfjlBRavaqSh+TV09fSB3pmB
JXiTspvZQcvzge/DWE1eUtiQZcvIuAOVs5ZbC+bP9y8YJE97m9CWnzZWKiOAc9i6
2vRtiMhQSAK2kXFrXYziztgBX8HzJUGi17SF0QJw/4WJPpDYwpJejpu/3VBUA4/t
R+ktBvSer5mgYKAKSr6IBlmOF/dCPawzIwfdSebXXmRBnksEQEJQx92Xcp2jIUnU
YuSMotctw41WVIuU/JETCClEMK383Rc2bFPI043tk51Aq01732H2l23uO1eRx7dn
tLj/MaFz9Z/xzTx9cmG+S4/AdWp2ozVqCDsrscX8m+Y7GiHWq5A2JA3vQ4V4S7pB
5QHHeNe7QhJCrPEFFdX2EfX+U0lc6KeWTEv6+VBdGUlwfg5+o+8y730dhJBQoZGe
Oxpd3wbIdA3ZWTvngNLwrEUDa4Lwgd9iR6JmMqtlV48XQ0RI3loagnpDqTm9ENTw
k1o59+SEsYG5O2prE9n6RPY3iU7d/ObCC7l0TJ+HDpGC+4r51ZNjQWQpTiUmOlv6
/7D1qmKRbOBbSA8zgJ+Gbrsq8QgNxo0/B8aymOSH1DwPqh7LHVIHfzzjfKvPUQka
JuXJWR52cN6DgXgx+YqLhMGHNQJPQolq8+bRdMX1x2zOeOsE3OMTtAFqNicpqeQ2
PuiED6MkkDRXEotQIa1F33mzg2nx26Tqi3cw4iN5/EFCCflXaKmUlAuv0xeIHSIH
bDXPeUEwAkXWJjnkQ81zK4NeS8rLZWWhfy+njfKhDW3ybqhkAJnNstQw1sOjooA2
Lt0oUyjyO2UplbnVclWuCDpP/ZkAn6HeEB3UdUQVo6AFhC/gS9/5hwlJVuHRA0ry
dsG4PmNzhNZ9M/gp0e8UQldI8/BpYU0iUOEfE/pG70mqjF71Shh5iJtIsu3MzcDb
lkLbJX4gvfVv2DqOKFM7V5p1AhxS6WT50cJoasSS8+/si+Dyp4H+IdFIa0FNCFj0
Wpx6AElApThA9vafECN8WFQWeoyccjzhWtf6aEDYL8rWhwrVwlLf3oeAl14SdqgZ
SGevIkpAyNN8UDL4vYfl6LxXfIodVtUylvf5McBpnb/HfGpNMiLeUv858icF1dkM
+wB7KyGxsebRN7+YqqUQ4U36mpvLsnX5QPQLdIv3FK6lIoTRmA/Kt8dWgKyxwnkD
8GwYCIGRRf+8xYR/wzhT1ZHCFeFmy8wZLau/hAnRec/e1X713AQwP3shJNJ/69/x
H6BPBbA3Mi1Tk3AyfvgndKHtz++Y1JxrOD9gF/seMfcKoLexZTbiMWuUCEe6F79X
ePHZtC0TL+ecGdokdTfUhFLnAHWHbAxzQ56WXj8/MYVxGAM5zRBZ2xX9qTIqUWFP
bsSwygidlX1aZYm1Th05Lad656er1135Z4WZ1yVia0YVIxxhMdn1MFBlZzWB5wc9
AySXOzgr/U05Jma/i/FqDK33zdh/npIKMQ56ySM2QOn+qTNWbCXjTqRtQkPhgQVc
OCz+6SB5KOml1twQp5LjbkkvzJu6TvwG2tfYOU3GZpUVYFwlX2YW4cR/1pyNZwJy
8SVAIbJS8BM4LIUv1V1S92otD09I8zaH+/af9NXQzElAjCk1kwRz/oB5TMnusWeq
bfNlkCmQZ1DcPecsBUX7faWC/4x+J7o9Bvm95pVsgQRsr6f83aMjY3ibfno9BNca
Q2ssqwgRlUQe272V6k1sb6PmHPMw5qJOQseNybGJEEe/75tAxWxh2mVgVZ7VoQtp
aTXtOA9fUCkqSlJWflEQfDBzAK/r7QaYU1dIDkTQt5YPeePoFF0YXY+9WfKOTqnj
+IKrhb4gfLpDcRzqVM1oIeRyJ7PGPWbb5FK0CrSq1twT4E97ggK4f5PQ31Sn+wdg
w1xoLNegLpBQ7BJCGecXvNvlHOUtY18g8N465ayXx881+OJQTMo6ZnpZxkI+zKrr
JbURZDcvSZNDA8Cyevr23XPZeCH2g+cPj83qavMFanmjZLCHiF6GGVSXKlJip05O
luz5W9hfixiOC8Gg8vggifqvPGVf0/tzhVXNLPn6HJ/M+xuGhZwi2QhWFCCrBSbc
4GBud3nKADWK3suDzwPsnnHC5mvfzBvcOZiu+o5/zyrNWtyvgPfnta7ExFizVnNZ
QuSMJPWndtUAvf39URK/wnZfkggsj+Vy0DlCPErThD3Hkyp56e6M1VD76ZymSr+d
QvNW7li8G64YSIEUq8GiGliza3fza6278XvRaRaEpJaCZ0WbM7fzxgWNBW5l9nIY
+MNexZ+rYLul/hd7RK1XDFvclNg4WQiD4+9fQI0vAdWU1lIKDfRcm0nQGnMOq2vV
kZWtKbnZqwRgE/+fInwuTBISEbbGHCPRLGPK2l9FfafA8TB612OGx2XdFBJLX+Ce
KAlVp+uBtB9wCBavM8DkhqECG+untjcre6QYgyE0bsPWZ1sXUK2I1vNZrKyvJGg4
KMPMBnto0wIZonjIL2cBD47EyJS4mI0Yq370oWDLalmmc+MjivUu6mTmj3v9Je+j
BC79s15Xa6qfai5DlUusfTF9kudShelu7G/HEFLP3Po5H1Dts3xb8lLEoq+lmJHt
lYzdJUfDba9ctYHU3+/OZQfFn1FkwXxkBZFN6rLWYfGuyToXO/vsv/ZUiEJ/C7ZO
GQyHVkVByV+EO1uFhUi3yB5oCh0a/WO5m69qRN0nqMYEWIUJG8h+Io5cDXbPF3tQ
xINra5RPboJsNJO12hFhJyF+Sse+t3NQDAmKNWbXNWfptbuCFMeVYxyiUPtDOMV0
19VDTu3lMR7jL/TDXAlKK2jH/nEfAyVSrGe1GXUuffIPzO2WJAJcHbXgh9x/qLNL
iD+1mkU4u8XsoUNqLdMKBqDaGIF8Cnn5A+PCCUIZiouWejNz47/z1sl/kcHzDbeV
7Z3W4Vs86AZkYjCgqnkPLtIiTkcZlCNP0cPXUhR/jFJeEFAi9vX29R0KygSt/Psc
oYHCG83n7kc3GWuCU06y9WLMEjb0oVJ5MQguILLLu137qkPTSkhYm2al7YePPjH0
f22NDShjyQnNv47CIQpZA2UGauQd9PVfy8YQYHQSheKKbv6HUHSr0D2k4sFSt85r
WjgX+qfcfn7LQUXQzwoU2UD2yW3si+tKMaF4WXEFnF9SHTaFQkdTTqQTbqdQmEn+
AzCzOiIpLdE2zAG2RSZNTKGRvAkbkOwiqO2KMAS6fiDTVKT3AliQR5XE4ELEhYtn
SyiUHrvDa9+KFt6S0Zf4VvGQPSodazTfhlppFE7qykg3yvNbrfMkD3t1rP8tRedh
mSLi3atmm20hsjK2PizAlzlNBq/u676ixaqoTiZSehhnaLvlPCqyIN44aWGh1wHb
buWc9kBVamGitlry15wJlyPHM0HSbQwTiuXmbnWMIPKgVI0S96KXwQVSu96gMZok
3B8IaFd254CD28puxKC0Qvaca4h+uI0T9rpoPU6dL+vZThfGO7Q/Nr0ZXQtGw2GY
m9lo8+cRtEKfKeqWWvJWoeVr8FzMAdSgt9wYrycvsf3SMg95qqH6mACzOX/kusQI
aEsrPT/TD3x9MKD/C9t3dhAgJ4so1TBu655D1gYQLZKVOX+NTXnIA0F0MezG5R2S
p2Ih7RWTwWgIilUBjX7Z4DXoKz25jrBdmuXvIpwU6y/esfgc0anm3XTYDauj9URo
AsjEivwySN1Nttv78p/q68gUw2U+b0Uy4xcUYPvGEXUgJO3idFAGriemjubOqnvX
y7H0wUo3LYP7iOL4uT4ldR5nGgFw08rNQ6ghPa06AGdHPxK8fn4ImAU8V2/17MBY
hzUW8mgrmByf43un1SgU79SaSAkYTzsxcdrFw3GXQgwCll3hqNW5J2Dvl+f13/7B
z46yh+rYjp7Pg3Syap9Lm9/rqEjqPsuwKAnugIgbfH/cjlS2/7rdyofoIv+JTM3F
I+6N60UvrQeRS1dpHzB9WwCTqi2TLQJF3To/NACy60uB4BZIrnu1yWJ7tQraz5Sc
24xsnHe/wNIVdawetUkbgfdlpJQxp+BmENtruPQE3nyhyw1R3zf/wnWbpbttq+Fm
UoZ1ZFGokDwigdrN5HYHX7cpXke0UWGFiKC4NQAUjVcQAFV0dOmUDQWrWz4+RU4F
Gz/OPiuQPMi4kMed/5psomCE3PpzhYm2+RvAbuDfGf4yTDs2JruSTC3j8quO6dtz
acJP+lciQ7HOx+aZ4appsFWMtkV4btAj0A2zivlTDhYduof6mZYZTs/qxl6nFgzY
pobuZJW7siqvoT07N3S1Xe03d4ChTAqoLWHKaha1ToU6v3fXvYco934QpDGqTurj
GJoU446Bmg1q/PRl7LsQnIDbgyA5AJ5H5hf47/8CU/baO5AQA17gDeIEYxLm+xn9
xj5Za3XxlgvWNSHHIdX0jPjS9MXCraGa3n+dCOMrwDaJhFOmoN6JvUuIUmRGPawv
wZp0W100//PdYd7gv6BLl8g4J41JDwKKtFSKxPbgQz2o+qSRkGNohG/yJERQnI0T
Fc5WemZH2vGkRGl57W18qfxL3AZCHcrP+8Gum9pLzz4e5kiV0y5KnlAn+IQwSqm6
gBTzYI8IEtODc+3/lqxPVBnO3kpUIdYLgY6mAV2CuC7Y2wg/xKXa4j8HmkWDV1i1
jxKPcxCMxTCL6o9IoDYOQD+3SsfFAzMbxpqn/1EhE2aaXYuYmRAaYVxmHbhr0QhB
1cLfKqkF4OsUhUqrly7tBm2QCpuIh3JC/qutS1hftgx/1AliawHZTVNnhzdcpYgd
08+rgtbTnyEF8A81hFH34EAHhlpC1e6GNWUyaWNbMSxvz7uI2UwWGe8MEaBjFogn
GI4idwM4OEfDPhi+P3VzhCPL+f/pzMVI+LvHDbpeNGOZKJKqyO2X1JL0lU39uObP
SwW4vP/SLNQ5rteq88vxXkGEn3eHKvKxqQ83O6FQINSpnx9wrjmjoy1THJfWhVmt
+S06qhUGQILzJzvOqBNC+AZoxxOwY1Ia6e9x4Ubrd4XJ3kpecqzS/nrQSFzavCv+
HceDlShi8pyh5DhCIRqEgaVNJqcxhYW4m0IOhVP0OEmce8VNvepIXn6PQah0TI+z
mQscRh9hgIP+UGR8FTZkkGBC3soro4+wi6JrYCN/tFtNbFRm/WoVZ1YTxLV0ZGIk
4VphiVydNdUzhU+SomDWdUtgyFdPRMr3PBHP2fPv4YFfx5/OlWwIlPipYvOjNGba
wy8SWZ/VsRy0Dd/YbBBTvTRqJgs/rZhiqzSLL0ueqZxOi/Z13FR5q85YI6jSN5Og
aF0xPvbPl/3v+YX5eJj4p6up8TdXuyKyr2VdnpT+yT8w8yc3fHQwvtCbb6mkEZpS
d03TATf2ssi/2AeJ12S40wwnq0IspLH/IwWOywFpaXsjtduOdvbBpaBP+epXBWzR
9+Sa0Hb9xAmQ3NuaWYbM760u79KUciM95CNfmroodfwovqHx6xdcDOOQ45gZoKNc
EfUaLnIPFVib6sH6I23ob1u8kJyiumi7TwILXJ7NjhBllyRv5LFlEdSsEygSFbfn
tXSTmcal8joGEpTxvKKQjgChudmcq4BcLVOZbL2Rj3TX8lCliw6vFeTx5wW9GUJ+
G44Qp1poveeNUOjEx9ME/MjDyE0+IZ8W/CFQ9EkFRxFhTmvogqiZDn95yuhwrt9+
Mq0QU1SgA2NGv2MjSvkVofqAsfGeG6NECSN5XrrhtIoshOqrCruH5yPM1OAK3f1L
cG+StEbC1jnjcGAbcqAKqdMEsZ+o677hPndhgikvTVRjrsxATbbQENY2Oa2ftHoh
C13ZdW4znh1YruguQfH/tawQwfiiFiGa6r/IL6jY1I17KRpjc0wzcl2EXHogFOKr
ymRR7lwaqO04KAIzJcGNL4U7azNX5SqLH3U1fqgqflsi8Fur4+egl10iStuWLG4y
WUEbCOPmLLotzbV75fNkydEGK7Elgu0GyY1rgR2AkI0HJr7AEpqde1ejMyZOFp3V
7qrMubPhs2rEJE86dLUeV2esxre9nr7wIQepxuot7nwpBffAI3t/gYa/xX9Mn+EE
PDvc0elBt4T4Z66O7Z9OUuCyrVmquKyVryQJxHCO67t0iboETTZjXpNPjyf5+m4K
l0/RsAvE5I8+se4W0ELD1V1dcxpZIVIyHAIxjA6TbVy41J1cXv64DLChbARh+XwA
KTTUzL3MYqB52DVt6XocJxw8uXGx/fV5klYhbjDnslEKcKBCXrLOCqYcvr2oOBMB
XwjzQHPW8EgI8tPpQ6Hx8Dj2YclS2W9lqPIhauxHb6gYXbiFOnqLu9RJd0Zauq8X
Rl9le5o9mg+MQ61ZOHSAg/Gn4bS29yCMfI2a3TosfeJ1YZ5Koc3aTXaxPdu/ax57
ZYDRvNXo+xvWCmr5Y19+l83+h8gm+16gMaw/OUU3lAeWonGiYGpTfR7WmqJIeVmD
H1ceCjjD2R0X31qriByvqeuff7J2A0grf1CePq1EAJy13U7QOL6O41oh0IMD4ObI
ynG50Olz8VFxA9WSHNOy91l6XaCnpgLjyfI3VwoahEZJZUwnP7KOTGbiwqBaR5A+
5C22c2WvmIFJW3YkqBCZA7bnpY8cBXX1kI/DOgRieLz8KO9V/ciSJluxIThhKnSz
0YMGiAOZPjxawXEjoqpumzljb+Wh4WCmecA/csrRIS6RypmMoJw8W4ikqydDomnZ
XeVTWqpiCydAWkrJRA5NlddjIrgovw0Gq+Nxr3g7DbcMVvxdPM0/LGAdGJB+VT7X
ErqYyLhYOt8zxsUOgK9/2nsVoFVk1KgJVmKFWlb/0IMoMyKbmWSNn6rs8Cwpr7jj
JI9+Loox51ymvQMYqUf9nYcwPKgP3uQOwb8ZZkfJXb4uGiLDrcyehJU9eeYrspps
SPFAHoVdFkvnNWtg5VCPKzRpaUJ1aue+a8Xr/+SIZfRxyhIYoIJT5P9wvOdnPTFe
VHS1KcUj6CPeNeQj2cOvJFbqMipngrMvOsZ3SXEg8hHDRug09rXGTIyGGIe1L1S1
3ZqgsmXGu45iGGMs1aH9M47dwq7KMy8vMQ9nlBH097ifxbtRupOKo7byF4LbMhOU
x/TpD+e/eY4B5DsRtVGKM5xat1mtrcFNthNkjdEc7kkoUgnT4+GHFzDktKnOMzDy
XUSZq65nPDDEVGoVEuQs2GrnfyK8FNDAptj6qrKckg+ceewDhC2sPz1OZ9no0aTG
al2u1tYyViGUlFX2D0wfkXgj+IkzrDOzrHFfHs+RJDIXgldbekg/TYiArTXqxpd/
VQe1grko0fvaFL/ZWECg5tA38lWYmodGdAtQlI0BcWQ6vfTR+7QymKDOnybKzOej
47O2JITKpWTuitgcydVJMQCFPjzMNQqAYbr0l+kJJQySr5XPVL89YI3axvBUtdwp
wmEA+fWOY8ibMxX2WAbhnrPLuQ9gIa4g8at9qQP8UpC90god+Q6ixm0/uwBlxU1/
K1z0lJBI6mDdzHNqV13T3drFk6AHXo3XeNLoJW0oNYp7jWhJzGKF4pfHPLYcPZJ6
2WAB1yn94lmwR6IaydHr3BNXqq17rWZTP2wSe6v1pNzdnUV3C2AuoAqvm/7Juu7U
qBEGkzOKR2lf9MruVX8NjhNF3vmikPQA6AipS0KvOagGhWTMiHCKioCLP/Kc/CRq
OWcxzMZJiy5/2ITvkS6Y9zekbF8qp2UmCN6Er+aPg3nZwq7jDyZQ4htSt6z41Klu
RufyxUjOoWEfp22eNdn1WL/EUQnG16hgj1FMta98oXQ5tfziIAuvfJ/SULwHGeOY
0ypxoypAK00Unw0I6bGYn06n3eIAFm4Vmomd0Rq0SBlpycYHBn53b1IkV2cpfb9w
8kV/sQ3++O1pHmyEeLWeEQXdDPd0qONXh/9Y0hB463ZmZetHxa7TleXLqEEeOCYT
3bVYwXVy2X1Tqrv4M5EKvyuWwHXJgnvmxqtnGaJFrpeNyaZpFRHEGyx0XH/OQym8
xpcwnj7UaNQqobb3iJgfYGsiyB5y5XbCbBUJ1gJePzKWJMvoknhc5KGBKNV505E3
ravmZe+UzGQv3oasXk+JXiBuuiVi2nmnnuZxTpLiPbtNuEeDU72x/le93iOCzZYx
CVDO/rFLBdrYyXAI1XfmgZ7MpqzX1GoF0Yu+Yu9ANtGeSQBv5iJY5mxE9KXMPsuU
jAwfQJM9UI98Dkp3jCApfRi0GR6wb12BH1BqVi5lNPkspt6rLQTFThDuxEs2Fk4W
C8YB+mYMOmuu/Fh11nltkDcMMYPgQUzuFlv3lXP+RC3xV2U+3uaKEjOlHc4ZbIk3
3Wk8AW8jkFwnkKlzWMNwwjxQnJbqq1OsTJiUtR/eQTXVVNYFcF0uI/4kNSZ7pwtX
BV8y93RUIE+wayHU/Rg93EkSLJ4ly4GmO4W92sqFMjafFVQWogZodMDSWzANAPGO
C4JGpIvNswBVmmvWJz0QgZjgKrzYcAyHhdiOxlXLNiIQoetUswvZk6vVB/EZgPX7
BKAcWmdSowg0QE0DEUV8awIuoFkD4YuopqdDLGoSZxiWvsdTpc04JemK+ymR2WF4
Y56lRhPV2f8FPj6+S5jPpKuJU1f+QUgop8HG+YYthPBlvWEldHnugBx1MomtkXwo
zMnprvs1vv1ojdbn+50tRDj92YNOTgsFmKNTSTa6/svv1PAeWNBqZKW8IJEc5e7t
fUVR2qDzmZL18S9ZvcEKZecyy4Xe9UbiceyIUu9PxHrdYnd1i2QQxoTdmpEH0kjp
17y/2i7eUzu/Z0VWt7RCPvV7Y2PuOPbnFMZ592vDAcsomBcbHBo3qIqqRiOcMxRq
loCW5LTxptYzwPH1cisrcUv4yeme6zGr9yFxDog+60oRDX7dUVkmrD5/C05X922G
SDyoxNnR3xMz+Ga2HGXP6aKgj8bZ9060cWfLW37DfH3grytpOe5HQqYSQbhrI1p/
RmIYFBSv6RQB2ka25DyLaochNjVvRJ+u2Iy5scTgBqPbo8GsfGvF6GSdA1Jj0UZe
LkuFyj9HK09JYhvp5MXaIayt4OHfylAqGzQd5dt/zqEBq/4/oftPXyEMoe5OYo5y
mija2VZzXzIPbRlH70THKA+Gd7hcIjhn5scxek1Tn6CoB0Q4KKWMQ0qTPp31ylHZ
Bvupmum8ZYDr7Oo8cTVHplElgiakwFYi5F5zCXyzFNIb6/rmn5ODYQoVlY1dNi5b
gmbM+vcir8PP9WhrGBgUZOKJqOEZ6AzRRKXQrvTAMdaEfRPnI4ppOb+fuaUj6mjB
Ub7/t06D6YCklquKTgRomyz/09LZMZkg8RA80/hAIqkSP17u8ImUpo6b5JUmdxGh
xbv8dYDZNgxw+IaJhZP1m2cFGlEPj5NEy8BXCkn9QernopETnzdcg5yRQH6bbFP3
Gkeb1aJnnBWIO3/HjxqgeNmDgUy3tcx7BG8HoPbo0IKLIYj2G3hS1YQrYRGYhKbE
yVxDM1O7JNEo/AY3DE6wTqLSVDUIxdb3zclCTu1GXnXfIWBjNHhznqq8zm7FgTI1
bWJwSzRGlzhvIUSASVSN6jGe2/sv6P/Qll2J5/DlnX3mcfAz9rWfZeKm9inS+sKA
d54b6ulBAGaWTCGM3LK4CwTQfDCpolYt4tn344uyZWJ0yoSrtZM0K4sRrpcovlE8
xMW7H3TXv1hS/ekodyN9fD9z3/mTnKDzj6wOXU2o5lfuy8jyysR+0dD10nNLweeG
NtYWAoVzEwe2+HiEGLJfcJ561zj4RcNea1A9JYjTlSQQmrHoHCRshnD+adManFPr
T/PMR0/tG/l9ykwLIMcmPi/MvJ7zc66QEvZPL8W4lKt5TFbC6b7EwyvBZyJIA4Lj
Aka8nuGtwzZw39difglhRhi0BI5FuJ8nPBk7gCRPJ9V2TcVC/5QaQUaT/Jqw0bf9
2JK8dcp0jgYMaDmI17roS7W5Upr6qPFl2Lmyzhw/mfOo/mTil0E8/IRkOhqGrDWO
+uwX8j5dm9w2dxmAZB6gHgw2rdWdKx9EK8WyjbiAkmVk+u2dbCnnf9tspZVeFqPJ
z+Rkr3SGAxf0LJ172fYb+s82QxTV7WCjN0m3focQ7PlxOw/tz85x/qI8MqkBI1s4
22f5dPF2WiDsC6ydm9DGjRs+sIjzVEfFodsJ9BmmqpN6cdC3mP5LH3QLDQoHFOoE
IupNtBDq1kSoDc6BECPYrn68lpIabu9GI69T/Ex4faKMPl1qOyXp5sQ7lxSDMdCx
izljq5DYIm0Knr2M8aBIr8V4X6eRcOU11YgXWh17pJW97XwmwFdekZd2IEdvgiOo
EiDUIRJhzrbTU6rMRCxdFR+bevKoYAFvv6Sumlj0o7YmBZIefX2/5JJ2MiRtrUER
eE1znzn7yuP7heilefjogyCxXTE9uOjMCmTORH1srOLHpnFc9cq14nFJZswh6Gxc
PQKu0/jqntMACaGuLNZqX5DxMvtbp3msfmbiC/kPX00iSSFhAhI0Mt2FpUNLLl8b
OM80omzy9mkoFcdrdFC+VRQ8927eOEIGEB+abcpb6y1G6b/v9/9GNiaZxX9U8Wey
3IXsJRve+OXARL6q9CHCUGzvkJAex/oONcWq1nnrd9CQekiHhCbRtBAbVWASM5tN
RNZS0nQHttEG1xR6alkjwlcBz7X8+TMn2jA7/Y9ux4vx2kESDgBWEAvKR5Lg3RBX
jlNhC2Lmj/icCzlP7aZsC1ywZ5zeswDAeormzO5q0P5VaC6QkN90P5rFewA9G4tU
kx/7dOm9ZRrHS1Z/Vs8mLsFPfKipv0wqwdARwP4/BqFDN1Jty9XXLSpw+PoUGNoP
Qq2REotx+UAi5WLyE7eS8wMNfvp7PbN6UzZsteKrz7jZBBH+0C7/t+7KRd+OiUr9
XqNTCFJmoNMxSyPnn3vL/G1knMrG1g+tWzUQaaP6gaem4+B+sNnKSuG8kiGF7KA4
TtPp3qonBZuC2aO+JTpLCcdRdRIMBdsAoEXJhtECGVdxp2Xt6m/hht/tEheVE/ES
KcfSedmXFw69a88eGSIYpJpAvrT4boBK9c6RfCj3keLrENP4JOScs6fMEwc9dVwX
fNMiI/O/hfttrzJ9tugWor/OrQ9jAaK6i2CbialShhHzzUjkJszzOrOtHE/pDe5S
XwPmz0TpByLcrfhS8dmey/TstIdkErCug5/lI+JntwcXyTZcn55UHiZtz9sSdOKR
zfPlW74VxUjc+fjxZKgrTrUgx2p/j1Br8XxRHPlyj/cpB2nUEalm4v0Sk959o613
AVbyAGFiSArMs01Ql9nviAMmoeugK0w+8awnAHC61QnZ1/B52XOlWaWr5/kIaEns
/e4HsvzsoIIK2eQdD6oqRC71DdFj24hUol0FP/whp7ac8r8F5vgHlqvaFxTpjiCm
Io+t16VXpQaiUecfUkcnXdgySEd1bi25Ziaon9Zhkcr/i7CwYf2DmD4smWYTi8qY
zwjSyZ8vGdc4ITAsJO9nvEEAJc72MbkEzMzg9hD27wsTX867hm4cGDXrBVped8Dk
RPTKGnZAZb56UXlxMUtMB5x11NjSmjZ9HZpyArWOdeNHQhtehnUqhCdv3pybFcDf
JekbuSUO7Tb2PGr/9sg8pcbTWqkikJNNmvvDXTusiiF7FvcFTNTCu8lfR+FLmq3Z
MW4pyxP+T8U0l7+xETrsLj2etj/G8hwdiW2U5FD1einZduEGaD3iXs505QVEjSlX
n6glX5Rt6xSATyOaaYSGPNXIGaQliJ1UOyt6s7Q/80/UbdLW0/axq0AzAkU4cMHw
P3kEoMBQqesFgGuQ5OnoRWfOaiLKNM0bEeT7RLwVK1a6DRUqx1bPqQfosXCyHRwr
PajU1E30Nq1+wisk4zjl3QTwiLIHRy/pLXsx6TXW4bDoBK/v+XOYbBL1NqxOqzmQ
fJwR7GfDoGIDZgHr7xEWchbcW/2Qs1rbYoHjKAHvQpiB5HtSWMbpAU3xQxNCibz0
RRKgtht1CiYQcL3VuvehOnQr/4S9SydEGvRwz/xpgIPq6sPOcR+dWHB+Nn3SBw11
rSqRz5/bRjhLOz69ocjpVowINpfMpny77qV+IC12ndgoPczXLDrS+xnzg2OBZKCS
/4NidsUBycGjarcmudlWdXVJ1+aeVOEQPQPs1oCOphzsHk5+Ss99mvnyKajT9tEs
y1iLHO4VVFFpcF9u16wzNmJwBmFzLXT2d8EvR+9VRVmkmhCUKNwl27vSn08hHFO5
4tbYQXYwacNGAU30kgff+0jZV53I8zkBB/53ibMPdGjN3pY3StSV7WA/eFIhJHqd
EA+y7h8tYArYEoChLtD9aCugtmqSQr+9QYQGFJcwA9hNCWL8Ab6O3aPsaKJQSoO7
b/lh5JAwhjDhG1XV9s8RxHMVjw6yVqBVTumHfElfqdLPPFZk+ZwK2F2LWtW+UrIz
MCMOB0Uq4xrEHq3b7qW9mFTo6QME84QUnLLLZcS8bVijkxfTC0bC8rQ+Mh0Kul+Z
ka83pM3q2lUypvb/Q5yF54qm++JITjIp26245PSXhojOf5IqGWvNgkpZiQyHjjsx
LkqJBllzgnLE1bfch4zKqU04X85dkjXKmFOSQhW9opJsJzwWfSsK/PTmhbXR44Jk
jq9craFdkWMx4xiOA22ZkrCWlTlwsv1FMpUHEpBAfCAo1nLJp4QJNhWBnf1sz3if
mvT7SKtliXbZZF6fB6fU6+Tv9Y3GSBHnH8oUzCo1NVZdQ4Io8UujQI+oQYs2ed8W
hPYzMPYCBnXlCUaKHpMPYPXh+W+Pw1uiDXKuBvUUHE4G7Ndkw511r6kwaMVEfz7k
gJouY08gs4AFqegzMA1r+DZj1J+K2CBJCNdythUJR7gGdwcXfTgDInvh94RU4pCV
k1qL9GHntQxviANPbe7DCxw4PzbaYkPOYLy3Lm1lN9V9sxgTZTLSQcN7x6Pp+BCV
o8Q/suxpHCBLPVYhK/CNAneg93zlYsCY+5/nbC4jvoJi7blTlcjgx0KAKz8ErTA3
k66s1Pquwi1YoMWmSjTRRGuUkOSs4XYmLp1nP4jDv/eOy78EuoeD46vLZNyLB11s
Mbo1daEIX/9rzgvh3EaxjoDDilJ77XZspJqj/e777zvfd+qxkEResLWRQau+bvWx
UkZbqKp+kqEns32uJ6nXIxXkSN34HbodeBa/q44KRH118YsW+DNhy8BbIpnB5YbJ
0tv+wqTVsPHRCjyP7DneXXJOutz+GpejRWR345d/xhDCwOMyM8Rn5Sm1MmjCS+QT
tN43L7ft5C0Ld3G3Qtka6pNKOowAp8T5+iRUtotQXCQO/A2oPTtodmiqV3IOsdq0
RhpIWZs7PxgEQpJ/I5+RwtmPDiSxQtbH30kq+YhHOGORyNTxSIN9OTQunC8vEKzp
qsOFYzpwj8X8lq4VswZ7QyhRr/kUZC9kiexrX1uM9Zb4s7pCNteCw3NrkqL6ncfr
Pck8Dd+DF0djSteuw6nZeDrcGFfw+xylq+0u1yQgIVKuUXkPR3c3E7IjEJjC3h21
AK4YMrc/4I9HFk5+ythaV8ZJx3tSoNdd1TL8boYhYwZE9MF6WJEmk0lzyGRgfXx7
0Dhe46H7guSK0xtlfdUgjnqsxvMhU74rkv284Ef1o8plSsKZF3qyGZmI+a3fsn0k
W1vFYhcKYli3o5r4XKa7Cyyu8lEnIOuOXlfnC5OxjTtJwm6oltlmhOnkecfRkfNE
jdx6SWj7yFvAZHw3MXdH2ZFF4t3AonZgvlgz0TXMWbOPDmo1IW/tFq2hDnx0Xp7l
cL+U/v927mhiNejjij6g6MFyF6K7SJO7cxtqLG5PQuJgAv74k0fA/jvMbxvwpI6m
ovXn+9L9kt2pJz9yRdFj1hznArEH68AWe3ZS5YLvdXvwHq9A/m+eSXYWit40CTgE
U27GooyxUWrJCC5OdcTxqMZ5vKtilNqNaxDHQ2S7qsFFTgTXwoCcb4IFVaKDy87+
TTXJd1q38ZsfVdC2HNiqz+U0vM+q+SN7u3hqRPKhMVY9y6fxj+tABE/IRQBp8QPm
qju9m93ylMGBaKP6rElQdN+0FkGxno+To4l6Clp2ydGd4WatzZO9hSqHpZ7psriF
gA7k8MV1hLsYawNZgdC28BigacRbhNtpOnEyMrEK7fwxRio3eMM1rPnLAxeE1/gG
Gy+ikfTU55eWD9oHgy7T+Be8Ki7xV8cOz9GW95PFFu5s+jIrYfR9Qjed/4p34fuB
1QPW/joQwJNC2l+9LHtAzqHas8uojAUa5T3V1fp7m4A3+xfon6Vq2TPMJ3CUPVLu
wTM3rP45T9dyP7ZYA4yRrPVisNhuZ/qByFvPrCZCIDwvvwwVtdyY7dqEUuJrJ7an
JynwKASqk/uKakmATcJnRe3ytLLRyTd6uCFwZeEVybV8nmOeSvhs+wXOdv9+v/P3
K5S3PfLNO+whBgEv609rk95Up7HnyMEjN65EXQMysZx4atjJH82YHJnqLMfXCwmk
/vcQIwXOSjZorVxMi728SHlyhYtN5iMoDeFhQYfzDT/eUOyxeZf0ppKYMlQfXWp6
cakwYM2HPjiu8XnHujpUr28yzk1j9iubBoEW6rO8se76UphNUG8cPZddcxhgoP2T
3nGJFMwcTPJCfzsCj57GwsmlXGjRIn5NFZBMOZ9X2ZRtlQ0YTw28g1hQY0x15cTh
zvQr8UKahI5pxBPNOCqYYdaYpIJAHIa0gmCRljLIUQ5aPLSpzRrik4/3k9S/Jzta
3IY19blDOtBRzM8tbdEsQ+8fV4oZTj6gMi8WeMjOGzO1MW2JPwzMd9/Q5lzD2bDo
7AO/7cCotgTrO1jXMu1JnJXyEnM+xkXZxIzg8/0iqddAu8MpokBkNlGF5JhrsyQO
Us+LvdcvFTvPpnWyabS2JcXYDuI9UKHoioaavzHzykNWsEdcLIF35eUPCN8RiBSM
7nJW1/bmQ4G0xiuye0T3TIONpDyCsXVgdR3gPcDmr9F4z6VAO5oGY3VbC2pMjMhp
AMnrs2IYpmSxV09+5v895L7QU6SLJrdlvHiYIaPfPHeoOsT7ImEB9VQkttux5NHJ
NxSWyIyp/bcy0f26y1B563t5vmu3ZW0iMC1iKfF7SkzTgKhJ45kXRivYgOu97ZoG
USSQPmnpKY/rq/ElrgFvVLGZpGVxb/Cz27zFj+UMas60jh2b9by9UEQ7ZO/pD2gP
OstLKm/G/qsCoN5QcUkjb1Plr+na5D5+VmqN6sXs9CPbp6fYZ+Kk1HgfERRLKGqH
AjpKeEmwjIyo1ksstohJNU35yachLxPcOcP7BiPG05Hp0wClkOlkygEu2C7QAq+6
fOBpQVn+Fo5daUpY6OttJDawU8hOCAId1wgk9tK/SYh9o145XQCQQEL4HCc1bOwS
sneagPQeQp1Aht0ugiaYrOS43+3zxVAEJH8AK6cEZUbAhnGWC7RPzTcm0s3ZgkX6
WbYS5DwqUV3cppGJhpi961fhcLZpuvTRRbE/8KQXbskycycIkfT2S87nmNo3M3UD
6y0y0ojZUtBbsJ6kKYSudk3ULgQpH834//DCUIrlYvLYc0vmT2dAMd2DGdtrcwcm
3qOC+HD9Dl58CU6EXh1L+srK11Ru3lsZtqI6TLz568JjWrM61azX5LtoroKmCWTf
BpzNEcBNDYOum1gfUAEi7I85s9rQtX1RNoK18INd+o/WvLs1LEiVfxGWjNDuSLbe
DN08YDGLTkVVHmQSy+s80eOpMPaydf52tHbUTguZ3ajJ3d/GhyAFvgC552TcLs96
7ENPdJ08KALdC9RLeuyxhKjtw74dC+IRwUOEbcqQwq+C3Q3Kiz4anRfUcq1KqrW/
P+wKO3BGdLd/wI3XeHA/xXXiJ2YtRM5p9vFGCbON3nWAwpG8n3UWFEitBpVGgSLt
K3GdCa5QUtl9T+Skf6v7JZYVtOPvUo/JmjUCsxF6DzD1+51+GTScIQE0BNnlYnzr
Sz08zWZgK/gScsXJuThTIgu0sbatbh1qgyJIdUB9GtY35y9qbDguD7wvtfdFs1wu
v9Y7qekRcWWdkwmy4lCEMPiZhvUEQ/mhlAcLzbEqT3STQcVnOKkSjTtWJ6bkxN1b
wgxBmpCz4RqU/Rhm8BalRtzMyaSuDVM64Ars7hdtxSiMk8HPEBatskelJLKnNwNT
mO6nF7IrMos4mv7QO9zgR9nBDsSETF8KYSfzgmsekD4+yBewZf5ulH/HVe++T4Zc
LCoGrAl2lzXplthE60gohz2IYLllGiYU53F4YtHq00OZx8YSz6TZyc4tC1pfQ/7Q
RKUi4r0INl5tWvcm6qjrrHJ759oMf4Jbyr70I3mTWWENglmD49Tg51mb3AardoSZ
Ytdfh8gjZaVvtPeSEZEl818Sqw/ex11Q0opGJ/tZEqtL7DiXkLS5+4WIBra+FNrU
vB/17CaYOFv0vwXqhf+57l113hikyLFeAfij+P5zoBHP9PKAB8LUQZZwOHqGPubi
/jbQNxi8aMa8l1Zq/p9f6h7x0szOTLCg3bnsGB7WkdXhsyOwtNQMnTZKOrMocKVe
FF/mha9kS7o3wciIV8olr1CioQZM/rZUpAkLZAfl3Wiz/jpED66xR01le02oYEkc
46Sj32h+uzaQPhJgPf5kIoX1atMlpkEKbp5maAxZEf1pH23eNOHcjRPKoUOe3EfS
ylB2LA7/WePeBvUY4XQexkM+lIdFkcjn8FAy0v4mp1WMoL7NI+Kx3i0xUgOwIAb+
rQUY1GfDkOidZ3rvOvbVX/Fn+/c6+fUDoqb3j2l9naLFtc/OTIETmEj8ATIROm3j
8v0jjEMl0jEuIR2Wn4k8XbtmhVdc6kr0D+MGVjJmMJl/iLMf6YVcjvdEZSqzugOf
3yQAyMLaUWcxgqw+imKjC98Xvd9vnaxow/HOrXKq56XbF+0I2wnH+sJfdteBo7Nz
JhBgCxr2B6rQGfisljk8GgA6hCqyFVtHebrtY7wESjgrqbrNaSH/2SI830I8MtUM
00pdi4nBpa3L/d0BXtf2+OTpfw+TXkwyXa0IlFeCLOnyaKuj4+3ckkv50wxnRXj2
oQOXiUbbskwkm9OJ/nZk9j7iHSGYzZfoLUO3ovUqRDJ7boo+zRIAmqKAQYeCEvZW
gTUyTKmy5V98d2glwFrpr/z0BRWZjo368lIpH3/D5hJSOY5qC9DSjkAOBwoW35AC
AuvDdTxmoNvqS4FZianRgj7u01bPGX+cSfUA7vYVkC/D3nGchRS9mL0bFBqvFcTe
iBeLRv+BSbzAlJ7K6LN2AlTUNKFvCc0lyisaM4UfY6ofnk+xAjMVWgeJ4kTQ4wNn
S/U0qGtg0KjXzs50BJ24r8OmPF34p7XUiMly0QQciptipsGUC6wm8lVUu6aEiqpK
Upbm2lfXTVWHTPyWMBmBZ17TqPisJb0SwdXkJpsvalnEXThfuU0SsH1LhrqzHhRT
27/vUazNFpBa8OIop6kwSZmVZqZ7+8DhxtnRcWUSiiY23qr67T0nYW4N5NIgnFMd
DeaDhiKBj+3vMkUx7y0kz/QvqO2uzJK63UUv0WNUbUAw/y3/slNdlGUP7Vi9Q1/U
bLMlzLqkfKW0foTWG7P0MAr/IGfsSaLrs4fmYa3hiAJlp762yibv/wg6/BOWOWeV
M3IlQlN/C5el0q5VOskWbuMhCnk5vs1C83ElbVI9hfIK240GO57NEFPSI+B4181G
+44lVIt11xvPZryqiVmnZQoVxYA7O8vB7R4cFjVLs4puCaq6lqqyufZC0+RKynmU
eUZBw3WVMMGazNmkRukBTLMKCyEbLgyaOwp9YDSATK2CwAbFMA6N92O4PiykpKae
Z3h77SaOtKAh24zWWccgbUQMkJg9Gx3GSguyCWShzOc4L0OXIbm83sBHOGvnrEgV
HW8vsl5OyPrbWQzdKPoGK8hJ87Q7+dL7kP9ebbJcN3JVd7S7QYeFHdzIR2+Br4Dz
67DF1melY/FVFqUEb4zAntP/oz2h+krvFgi0FyatSOHzeon/XaJUmtMXHh4OQEqI
VP36Mnetd4ES7VLhh1nWzMZ530oSxjv/zWjbZs37tkL0HNU6E7kWAywXe+cmQYeP
3Kj2o6swwDkcJCdZrdo/I92sXn1M3VmfVH3rfWySqWP5KKFDm0bF3dWeIRzy1RQZ
wnxVTuEf5gpFW6WQD76K2nfDQBOyFnwmtL+FmYj90DI6l64hjgeMEz97DWuA2nOd
V6x0ot55XCFs8zGfL3cAiGXG9SVx5/E7TIqLxjH96ImXc47QMbocwWyQzLDuNi2o
JQxDl90WUO5TSKQamthEu05+6J+1+T01VipAJKZTb+atzVBp0xlTQsNNuYq87uht
qWu83rkHURURdlRBaowS7uL3uAccTLxld29lohkZ58nlpDyd8TmTU42eWDqsXccj
PBtmNCnmUFHLMY5iToplqR5MRc/RBz7o08bdgQjIJZcumo57h1dPBCaswv7a+XUX
wbRC31P2dGoxmObbn6mmigoVj+CS4og6PsKubwSesKLpmwlHa7TIuwcf06VRvB5B
Ro9YmLV3GJxUEHWg1l2rdQqMPEdMBYRVjpJPTMiwAXKN/BjPJQyPd5bekNy+2yFz
e4CILdqZQL8fAR+KFGYkEAkR/Jxnh78Frp+yGKHTahtNaDIEWOnF0FtbJIFq87xQ
dbxVfrtDOk3puHOQwpw/pxiuQljhbTUcqRNgA6QrjPVzDqI9IflPVvaf36jnkUz7
g/qHbhvF4jp7cukKyRtNSVZz+UTaOAGlmCnfFBtg++dRqs37C2jaKh1Gz5w2vtq3
J0nligCXRZzq7CsjqfDJaCjyNNU2kj6bRJhtIJMNvZchFwSwEqguZ804M4rifDSI
zW3L5cQnsBobGGvdhYsEUFuXuNTR4OFFdoNQ1vFEOuBZDu5PNuNY9kfAB88LlW+w
Lo6JDotxv6bnrwIs8G26BlufjPR41vebeUMtQdQ6fttR5P/eaKnLl2rzutEFaW3n
t1He/EMMgGc8Ss4kFacFUpFHxX1hBIVA19Z/Y9VIww0eqNvaZvn3naPGCiqqqUsn
A9Zdx7LhcviqXqPxAP3H9K1u000Isytlo8TUL7mkAw6bCovAOqq5vbm8wHmPghvP
crzprdJ7AFilhhkX+HrELen4kFBQpKzg8QsCNmEpoeAbAuofU5PnoNMLyZrT4a0z
md+ZOlne04mrd93g5REhM7uVxxM7v0UAr3rZDG3kNEl9wnG8hSXj1vPbBPD8DXYS
GNa5OmkOI3M/GuEnN1DvqFo8inmvHyvgP4Rvw+wA4ltXESHomw4w0Wg0m+zp38sa
Q8jCa+Gf+WW4TqcRIQieEj9v+cpfdvyP17g1fTkUph+ULGHljtgY4H08+AmA0Gkq
ql/VV7LgVnz8rIGWcpbHX1xcol+fSK3uogm+USwiDOT7Blry+g9uMxo4VPK0X5Je
wx/70XFcAGkPPTmdNTbuYV8L2OGohiYKmteLgA+m1c7YAzawyg+C/77LB60c6jvg
HQEXuUyu6ZNgvMfrg2sOitjqGECp+zp3yI+D+EYvsRmnQD7B+BjtV0lcOWQBpA4b
0GgmGv6sXuoaCmKW8lUIOs/LYij0AR18WPjk2J30iuKMef0lo85EVe8p1xqIOcX4
rohKp2GfA9C8qOZHLWswZkCFx5iui2oCoE7PpnKZFKzEH8nD2Pc5BDiOV/p0TbWQ
HxEyViDxMysTZMvjQoPK1WUWNJrKi4iF2qaC4/pEpN9cFSaeEpIrgKR+RHTo9zAa
IDkQfRJlfPbAGiN0v/lOGmJ/9iiKRbCPsnZJaWPzucQjY1ptE5zlKH9VktTRy0sv
WvkXg0rqRLMTREkpBWUKAtE2g9kzRWT/DWT/7BJFa52ygVCgfjBdO1wvbTzF8O8x
ofiiIaYH3gdk2B4tgpijrpJxLUGNUYTF6qmepMsrqUNDCHpTaemRdNwtX1hs8Pcm
y7pjOH7xd2zKBt0TEEFoxHy328DWRn+JyXCp9DPrMbv7rFSUDz8bjG2VHEHwFn4X
an+5Ruq16MqQXMvoj1QP4ruXiaDkbLqqZJhEbj68dlVbYNpbh2rj8XgZPaLevFlr
5ggJfnM+iztBJDHDFsjHvB6LoJnLMJTZq8Qr14dU8TtS3m6et8UZgAwz2+FVeL5w
Ra60JeH0Brd2i9rwW+5QsE9eVxplRzTMa8zPVbV4GwjpraM86gi8UofVXQNCW4vK
J2LJkFqWjvLKAv1rUHKz/KHHqiLV5Mze+prDfESZVCQF9jbyjaEPV4OJ07DavdWZ
4/lR04u3pwfYhy30aj7go14QfuYg++OIEmJJWDKpcM4g+WykPb+kbdKh+piWlf/S
L1Twl3nI1QojruEX8yYWXNa3byM5NTFlsUa7oeQmGRI8l744ILUumL4GyVOvIQuO
ABNpIp9wZAzwm3UoTySiXrBOWd7LdMgf7xyXmOMejqSmgCOPbDoUwf9XR2mKdDAs
+vx4xL/wSOrNHJq4Yrlzfm9nvxKBK1xvCZphPhoQxAXoM3LPDPvHqc/NWQ9diwcq
I+E+QiQFAfPGETX5FPF0d4i720NNAkfHsnxK0ynP/aH0qJZvmwToDKiTXM9tKnOv
W8IM3MLGtneCaoknAWhRG4HeyIF5BFjkFA27JxgRjxPf8WjmGgo1D86OHWP2qB5U
RNBVnLu/LIWrghy35WPbb+w1wixtX85Q41WRJIeKNNQ5or6DyIec1Bl4jrZB/n5n
T+3X2lZv9NB/pkISTZdLX39ikTZ/YYBZcu/yBdd5MSx+ivBfka1d2inpPuuMbql6
UyKJhwqsdzA1evwSoNm97z1nOLkRfwmOchkdoRF5QbKLPK8jt0h8t0OzozGHHvKr
SiQpVFtm160UvBy7txfdsmea1R2Op0xCqXx0l7ZYWaEQLahiODMoiqHYIeb4k5H5
a1wn9+aqb5CFTIHfLZMBI83wKxd7CYV9Zxj1r/2zRGHvvX88q3zA0Rdv6hmh++kW
u330fu2jT3QkkNAuhCC9j8UM53v6GzrwGdRxjjzpiiLfVcoEA/6WhjtmVI+KYVNR
54HopWf16WJ5mXMinI2gkz8Ie+tXp/Lf6bdMP61AVnD55aXJJKRt0z5n/mdxQzRa
f5gwdDjF54mQWeucdDxn8+4XvIeN5X1bzcq6aqkaopvDAGKrD7SThccZ1MIGVf3V
8euDJcyv5enMwdw9jk/cMyP8qMNVjp3RV0HCrCH8agTIlRSx4jjx/PI0wG5OdDf6
vUQvNo+PxSyHFbW4PLu47tLtYlh4bTrn6chW8bvo3cnl1Zhx9OhDqZzQS2VfLF9M
Jk1gHUaosn9c7SBggB4rTPHJ3wXpeFipRyH/h1i6AaKCK8uelByrFIguTF2Edoz7
ky8uC/20dWHIKL2wQ4q4N1vqPZQNJajKruT+64J7461TKpNhsgoJKDhd2XXaqWfJ
8Ks8NyhxiLfUYkLAuw31kU/AKqBLQb0Kj2UwMeFwTn2mMvyh4BC8kq1xpNRExitz
C4PADkYEIfhnPycxo5O6Wu5ehrr/GE5BY3I2t/n5kr+mdETO8SWpO4XXmXzc0iaO
MUgtDS3X6KwdamHQLBCR7EJyXHNZjdNsIZ9HOxuZcFlKJ3hR1p7/K0qumeJ0u4l8
uss+mSlp3kiMuPnLtt41ghpl1oZlA/3aV98Y01CA8k5SGDRSb4LPcKyV76BsrrUP
x3K1YGq5Dwr6er8CwKOj/WyFGF3lmmmFpg/lF9XPxQ4oOWhTw6y4PNUIJqdHbQAe
9NzYQ6Q5mLptAsvpUwU2D7VozR+uYA3jcAjFqa00iYgOhTvhuY2EcZSQ7TP1b+pF
Y2+1NxvFDFAJSMQRt0M3H3Q0rMHp8Uz8ssDk9lWev5sgu2HWm7ousBAy6BkgmZHh
3j74vDXeHZbuAZsOyjjaSUcXvW8vaNa/TOIM2GIwlA+vJjdOAj4NLUGGWFxbaB+z
QzZLwhUQcu3n77WiI1aJx759Zgy79va9Ys3c3DWsFDX//fA1yqc+MKaSeRxZPLxP
2dtPs1uu1XoWQrCl2sqGUxowwXUcNa5qm0d8a7sSW9umcIs/wWMvEswgaSzYxvBf
r46HNB2R51lMWd889g4ZoPB4px7C4ShEqBSNsUho1g5eRx6i4RuOn3vmZLLGRyIh
k69wVm6Kcf2VgczvW1PsWWbqUSGMtGGJPQ8gfMsvTvmOSjX1YL6YwBNAEqJqfmsZ
iOdQHGUpfD+aGr3hgjKCW8T/tmoLkrLU4MA9CSHec+K7A6CMuf7AcZmPxksx9lze
XcXrBRiTFfnlWT5TOg1gnevHdDJ2Acke66SgJY4emImJQKfIwas5pKuJ4I1sOWhh
m/OSItUx829M6eonuuvmjh3DtwaAuuBeTxwB2EbYvDyLBmYYsfHtgMSJCzOl+eAK
i1LR0+Un6Xha/vOLVaecPa7v1lqDkbozU5YGhirvgbFpO8JrBNHkJijqM75E4AX/
DQxEf+HF671fSZBP1vyTqs4kDIGTQw72Tfuq/v+nIvelCE0gvi6MTguxzI6B7VKZ
o/VMll53t45CQ3XMSl1czVDzlGfB5V7bYy6GR0+exGPn2BwVDjYCyMfGZj+whFF7
mhEFlqvQHgLT66+THeWUWBv6QXy5MjbX14VxKcxA1pOBGkd4l+4Mu0zAfUcUDQmg
gapgk7AvrvHpsEleF3r5IIO/y5zMs6pbUixiED6qy39eJCAW/FxR9mStqXhnRVqy
irHM/TQN03wjJ//hWIr4aMwOY0/5TBUNTWqjBebzttmMQACznCa+exw3ksIycewk
8HYCw5tTypjEUC6W6sIrB8qmnWmIP+2q2JLwc87xqnzGhNW/zSkuHGdABggOUV3o
`pragma protect end_protected
