// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:58 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
iIt5qymNb01tTMJrvUR1S0O0/8b0DkhD2QZwUgujzx4JO7cTcbs3A+aHrFFY07TK
Ldtl4TMb3eC5TLcxgkmQHtX7g3b56bsDbwXzbUiwSsRYQwq0vwXwy+fkyyyO3ibc
mTEeTMqLrPCyYFw801uWcusTj/17/gffPJNolp/Wphs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11472)
YKwUsAg2AxCrQ0IkIGd6oYrhV/tcuN6eo04vCy7lDyKXyqkx5guzsoVsbzvbUzRu
uuMjtkQnDq5qBfcEaVPCRWSDud6/cox9MS8OVKQOlRE3/rEPgZl/UdBkYdStc9en
trTAYKJoXBsE/gn/cn5R2DjItSPiakBZafG3ygoAS9DRNxR480BT9D+lRxggdnir
bA3fFb1bBfToDa1RV0Sqv//iv40hcC/hgJ0lP7odoWcwulE/0qwQ1w7CZGalaAwh
88ixJC41m1+lYBQA+eTU0iUV0AvT2XTY7x0rW5QRV3zU9s+y+6zi3e5/lxNn+xVV
79869pSRExXAnQxvnwwJlgbiAu1NY4Ye3r1JEmEfX0RmicMqA4Gsxdk5+GM/TXzN
gYcIEbqewXmO5/lrggGpWV7lvZPu6Oa2628p8kAwjIX25O0l8++mctgOBCBg518Y
p0vPb6+luPXffxadoyTfq8PFcecftAI+qd25R72gj9y4L441e033INLQ9s5Mmfgo
S6nQ5EeBhgHc5lOrwfrBq4FbBhMMUi1Ml727abQMALH0H7GMSkE41wK309/x5Oi5
JCXH1c14qfU57Me4h0OxdhGJLpvnAFHNsAMvvBCLt+Jz0CCHI4yrdxDQrVXUrYjP
ZQoK7g2MuTwhWuCLXy7tXo+brL1EO3PVF4SaLwtDW5bxyfN+kP/8lmuAY2pqs1cC
yQjx0S4tjQc+rVxXkVD94trptZLwJOgL8Rw8b0b05vogzpj3ukjBxUBsvfcEQF2N
9tOZwnYqJtz/ev9pL0bIOrEyDNT/gWY2WqKMK7c3lf4oE+Q8wh5/maAVo0i/2I+B
aCga/vwmqSYYVqJau8gGxFEpCA80telcKRLv843M+eRc1wZ8R60GErY1fxAKbJ4v
lZl6ZbJMWKJHgoW7P+ryF2t+vP+UoPnccbQdLj/5wMTSyv9v2vDl5lZpZLnY5IDA
YiJhKXMHsjvUQWbPEMa3wxoINx9V/UoA/UAB70FKgqJ5YHyYLds3XD4GNQjSjPMg
biCPHO+/Subwapq1dxCSoPQ1hLj27iuCYCWwDLow0B7Jfe59UVtK/+1NLxDMX3t+
8FGzcFb2qe6VCUrMGyuAWQsR21QguPyRAkD3VcZwoqYlLfyuhWgbNRhbjAcaF+li
u4VI0chku6NUd2eQU30fUmNTHGJ2/RcJyuPzn1f1k3xzZRuy3lC+zLaGyjwDwEce
7N87dN4jFKQo8QQgp6IgyAAIkLQ2sAJnvDT4mCp7cZCq4RoTau1PKjzXgGDOM4zr
CKWW3AAGJbOsoBt+MebwLoKIdB/2xEJCqyV94vyBu/ONysd7GZ8gyK8EtElW1Log
MzAQPDb48bZWt8X+aYNFhY8DSLXnpDlKjHMkBZoKUxJFTTbe7Utu2tmPla5bPXxB
JcA8aWT26u16QYHdE2zReC9o1n2IO0wRtCAGhCG+kvZBohpemY3xdw9ADhihG1ZS
i+NAvrXaFPiSlvE3r4Bldb/WqDBhru4zZgPDOWFdIY2STg/zh4f7B1nxHvX9zNBf
sPkpcokUwbUxRwjLyBTJeZZeRp6TNVwPQZPIw5HiOQSkud/4lCS/phq3/xWnmpMC
eQDwDmlC5ecAcsg27sRYNlyPrGTTbk7KZ+zBzqGwDugx0wuFiAJ2KyfrzqR0xkLK
nyrgikyGbqoLI6jY3cbFwEom5rf5Co/LVQ8Q/YGvnhaol4CYx3EwZ3aEWzxKwySw
hWHIlF7SL4W/CVSwo1Gw2Xf62aZNssjimvNBwRnF4UfutyoQZiKyBpIGGkaakNGV
31J1fXaeyIcCwxk6hZgfNRWEokJrhIO3DwCq7cNxAk7QnyM/ojfxh0DMShN+tgr/
JbVVE7v9hl+c8pM+yf/k0anOtgmrLNmZp0Yihs+EKnfb9fCwKsShXx2owgdLb7oy
z1iIwtT+TtBQTGGv7oB8cuCEm6V0o1GbyOEQ6ElF8U6pzxozcMQNFWimXK8TK6Gf
V97fXxKonCCHrBXSwnvJNWEW6ogKl/GkRTaidCnRGEJMjIuqF1cfLWSm861zjw1B
u1RHWgopVaDeAjdpGywBSM3iUo706P3rQ7VO2hfCRERm4xduLrQaMsMLPhX92x9m
6mwef8sEslCIRMMKorcgPsmTY5p4DM1V3gUpTjAkLmpeaiG/kAWL7LcDFX0+wwZJ
bVkQIL5idU9j8PRyxNjWjujTs0M3znmzQ/b6mxcW135tusxQlDdilNsg+KgiP8/J
dYhEZVCDYdut+K5BQQt8rU0xSTK3DB4X8q66yu4dKrrNNq3wg4+8eorNcgV8/UIi
VbkmuQz6wK3fKt0s5t6e+Jzx7klExh3k+qfnxythrwenqpfA/1D5kWFQDv79OzEL
BLiNDYrUc/SKPnFsNhwhLzVMI43kfXWNTij0HipWOqn0vD7z67sMgIGVmzdyJp2I
aZWUgI2HWct6E0RcPvzSW41RNTBomviAI9PzFUNFuF8YrJEMSweA5NpGM6xYq1cG
LlpF0qm/TPxWrR2jH4Jsm8ji03i9pldDV9eCFsY8hEbvjOW5mjhlNyF5F++Xh+GK
tSnhBNG9M4P922kZpiAwIhkDU5CWrnWX18Zl+uEgFo2AfhXiHBN2xzxn6ZZqEOU1
B3M+Jhy3cCNMQekakXX6Vojd8gkFnsCIWO1/erJPV0/8a6zQf3ivMe2Z0vsUQ3fI
AuHUsE/z2pwAyPrknjaAjOMnpbPYahCRKYWcDHE/yVQruGwPKh/+zlBLKCfeLeFT
/7ORPo+OCBB1aFZN+y5MTojZkZF0cYKTTTupxD82goGM9DKOjbNeRcyq9kijeEQC
GWXSGHlMmQhrDDVCp6+LFrwt0B3fIqShw698wLUaTDRWp7Zrli7c8+EI/j+8UmQ1
carrDt8OivmwT0K5X9rJR6vs/RZNZgXna9vzdylRe7IaIibuKcAB5Boaf/suFfVT
iCeJjea735g42BpwY/N65dH3P+6IirKUdZlDwpssKRUOQEnPNIJjlvkn+h2rlM15
T00/EO2IbNqy+tJl39a+KXEze3OHxzaz1fqkS48re5H8gkuGRHh5im1m2hN6iePL
rGm5yR49mbI01wbZq2Dk8OXeC+f/ewGLp+4hgH3vIB1OF2wNUJx7vBDgvwa7pVbz
M+YlfH9lyf7eykSyWOs6hDjlFDGlnbrIRg9n29rknNedyULrhfDZSGERI8uEQjQF
x37kMaS2iDuq1QzZdzfFFK5KRrlc9w7kwkwsOlr6Qbod24gT+U21PRSM3E8V8o8a
uo+thbpz5G1F2PGHvxxLELhqSZKUv6WxVX5MUTGIoIGoI0fNPU9qe+X+5xq+RB7i
4WxdwCdcM1qN50fDkGHxVsnMWKVG4GOIGJRImB6Se9NhnWofY5jSOJQ8tCf2LFYJ
cHRaGICP/9bL30uEDxwtbqrF8Uu8FpHZPL0iPzMj8cZ17h9vmZZI/RtTrMaNqOoc
xMEb0F8DSZvAYWVB7eJhNDnsKMxCmCwdBEBScSigNud52g5+skSTFbvlD0lphzfA
lMBGPin8zF/Y6J9EiPOQWio5/l218bgoMb9hgug3qC0PJx6vmTbpm4Z3zh42BTVy
ZNf2ZWcwCMzogzJaD5KX3DbxPvRw+HQErpsdSKA3gZucaQUsNXNx/Liu+269cvNI
b9XESINoFONfqa5X8bB/zCUNkRRxEsR9lB3jUbrdHiELYl2S9FzN6WKbijLo+iC8
I+rfrgXm8DzRhMCDw56Otu6xkUXqKFtbaJnn9/2ZIDGSfkzW70usGOqD4LPO2F/o
pQcvqqV9QdIK8B+hpYUgIbbntYWakCCEMDLZvH5CbRlS0NRhdQ62mLQopDgwXWwf
pMkA2shTQk1/m1DCpfU5PwHZOLnvl9bwacU3o2fgTXmZyvziTcb7tBS4pCZ1MqZS
DjZwUQuJUHmRWTfRivTJGsZMv5Iq6LjQjIde5siGgD4xzfSHLtSJhqZDqwcpxp13
+GjASD7mpUCL2AoNV2yy2+Pz4bRLZfNVX9w9lMwhYDY3wwXpeG2OaXWj+4dr1K1F
eWeJNidlfaZt6C5Mm+rbMPd/eMKmFVVg4ZhrkCyfyRc4OW65lE9OBDUbxFGpl67G
bbyidR2pO3DFlvOyuNKwyy7d6b+WZjDAuB4GQqwjrYQ6R1uL4nAi8K+iVy53e0wc
q7+tVmyAQViGMVFWG6nlXUQR5ulnuosxEZJTmA9vZaLNZkSjlyh5RoEjPYV8g1hs
gD3T9fpSmm4xFFnM9lyaz9YAARbj2apbGbtBDxSg7vDYnE+RZ/9toIWFOmsP8hRh
yT0CF4MuZCueHu6KFXIPQspVU7eE/y1OF86IULRFzTwoJAi50NwRsXVRqvm3s2yX
uVDjNL0AvYx++r6a9FQ52OYGymLsMXnvx4ME1LYw/oWcZNJ3QNOIWAxWlQr97bBV
/XYaEi6d7cFxJBNhTBRGqbpkHl1pwixaXcW3SNSvMtmCt4PVzlXlqfouPDHgDvvs
kuqMOLP3JsIx64+mSgh/sW8yO/5ZuMzmpOnDqUrUaDx6X1dJjZ/yAx9C5QqQQ2eG
PvVt8RG4enMjB+9Xkp9Sq9COrE02sFN/VD/8K+hpBJB2xS+9LOcTumr15ncWKAhe
jDJdGHegjWr1xLibMNugY6gY/4OhcpQfdWR3zrZPMXCJlmG63yGzKnmBDcAlmZgK
rkiqYyDhdTZkWaPBl3zVy4jz2jh172ZraVplNpMhNGfYC3ipEbL8X9djB0K9jdh2
fd2SNFfS3WLGlpl1YfzzRyVnYvviGQKxvcUdTMkBEd8lGeLk20gCsp2h6KVbogeD
V+2XYdCNxQMx6lVQhupp0h8a5lwUn7KTQrBtHoc4t8SgWNvoUncW6t5SRqv/kOmk
I+VbAxB4Ve4wH6hghNVwGDH1wvM6h0avj22st+92QiRBbrnJ8G6uToML6w92/ETP
8L5cT7E7CPQ/HCTyNZbYRK7atzYPqbQA+oLzSb19G2u1gNbHLFUkkTSOs5DvWUcL
1HOMj/L0pO/s/EKX7SHtAlUwIoWn6Vk6HwdZqg5T4oVnDPfe0585ereWGrfJz0vX
pc5wEG5VaEyhwf0UBHZVWd7JDVS86q1HOhTYN98etq5yHhdVGoSMR9JCkTeBuV2K
UnUE+hiCq/EmLZ7p6WG68tXSQnMqvuXxK1ah7S/eGMXbiYn8TVchRAsmYe1b/38i
L2jlzn9Yyo0lYjFb/rTs+irtJsTv3PG51mzjXLN+qGgVGU9x5MXqE4KI86Jnn2vi
fhRcE9OrCduYQD/M2h76EjfNyN+a7aRVjYGqFnpwiL/WRYsLUzG4Ukg9GSJXtRzD
+EPHaxTev1ZLJdmcH9HQEVsA5WZAS+nvl2oc+Y5vGmkTRl9RqQzsFtUKVm6Tx7St
k1Xgu6kVliGnk2tHM5wvPgAoMKMiF2ggn1jm4J8GFOFpDPqKhXHlZQ83ereb+Ud7
reL9y3tM99+qmC7ZvgWxf5pJaZez64d+6BQ8XtR/ipVz5F4iWPFbSwOx26uXPCZh
Aa4324D3Ed0rcRZ+ab655Y2YnshZ4xsbEsjx9eKOVUhoxm7IH8H7bohT7t8ldSr4
63M8/YCW6oa5WJ/q7w4m7xUnSsO2M++CLNlQSPsPPOSmnUYN79iysJ6AedihcNy4
ivnIEIAK1XmKu7hfeUK3HZ68Iv8JZlwDtYffpJ9xwiKzipdUjpgNNfTGeYuIKWAN
7pl8hTjoMbSw7qIFFLWii5zdSc+JcTSML6Pt71gRoCHDect85Ip35X5feERzH/+o
oCeW1CLB/fQKMDCPFIVEJQKFSfB17gYiLN2iytkElxe1F0NeL+mh8PW7zuwt3JPf
9WzGseQk4PvMcDopr9Ax7t+AsbipygbGzTjrhn7Wr1j6kjrAADKfbMIWxAcumhac
Ecv3OX4p9WqDnFd/8Lf7QYGVc7o3VbF2YIVjM+/CtkhRqcoltp05IJcK5Gsr4bBJ
OzihMk5sXgGEmjClBSQjAMRFO2KxVQikbcPbvJwOhFGB0z525yKgZc4aJ0qjQz6q
CCi401XCne80Hb/4heDY8zPEBDH2o+mqUYolr9/HwOo6pTUPCpZLZKYgYQx828cd
ACLAd0YZPi8DUhmIzAy9HmzAJP7EipM30dOSLfrQkzCx4uRgn6p34cF+7xRbYwq0
0D+qrbZL4vVUDp1OCgx4DQ64vpcsN0SQgktY5BzFrcnjBbgh73JHZa7PCTzIKRHR
ZMZHcw8gcJvGrxgCuyFxnpghLQKaQRrmkfd1o+eCxpL2nkMIZgLberGhEouR9/Ce
aT3nezggpgGkyhAybAp+QQimxG6FsJODd5RIf/dYa/KAk+XU0ZaQar14zdp+2Tqn
cJ36IQ+8hvFl3O/cz8DIjTcdrH8tblm1wPR2PhbdYamO4HmiZz5+vDoUGK+0r6k0
HWogbuqU3H2oI0G/3q4xOlGwot8vmG4nrlgESZ5yUrm9luZsC77kVtlR/PxkKWWo
4szLSObGx6/BhH4TOpoMD/YN8JiJ5kFER+6sZjzPulNstwAJ3WD12DWiA5He5Jcc
hFoDr6vGQicpfC8pwmIf2lnAPV1YXZaSVKCylb0YtbVc5PkCV6l3jr5oIPZ1Njm3
hHKVy3jwTpxT3RY+XOk47dkntT2+jEYbxh0zjd4BRni60tHj7rMN/Faa9CRvoQwP
YYwqte8mYuPEiS/FPq2DBeZRCuPFd3U/IR/jQKj5Jch++QB2bUaySlA3MvrZdhhb
MvhOPwOxy9+FRHLfi8TasQSFRI0PxtQqjaUsrLW/ACYQOFoNGIZgJsw1gKU9bQyK
pzVyPG/vH1BQE9+jrc/liLjUMrQAw3kpgFqGVNgogOzGLICFczVw+adpuRtwak7j
eWmKNr8RgFqxTkeNf0sqGAx1oUopfYyjba/krHLdScK8SfrZiBTb6hw/So60ZqTG
egZD8NkMccNMzrN9F/v3zgWayJZ0qMME13JmJO2An4KLldwK/Nm/KfUFo3YXCEXM
Odw6dini+EvvPnBmLlYz5OsSiEW0hXl036gdD7Nhysu3zcBchzMMWeKvUUAZKJNH
nYcifDkb858qz92WAfdResKlOB4Hh9s1Z8AyrIGRilspEi1lSyiFcXlWC0yE6Wk2
roAnLSwql3L5QmAbuRbSJOkoCvNtsrqh8XFWr/+CESuPdvymv1TZBuAgKQ+LeZ9T
2UyNS6aRjW5PUhLrHjaYfSotqsvzwwIng/j4cV7jou7aR3yo/HVMyj6OWt/w2LtV
/8sIyoS2uwsUk0fCfPEKAIjQIa/HQMdSjNhGfjM+BgXJSgrnjkXmRba5Ul1bXgmm
T1Uh5qQ7+M2Fav7ad+s+xidCJti3S+kNeI0wgigKqbIqJZ+FQJs6FpXo6795lWy5
IspcahY+bRaf5vnRn4FVWWzvlwLd2FqWChVdCLkLejERQoVzTX8d1gcG5Z1M9xpL
Mbm8HY9Lq6sF0SSknhl3e32IbvmEz24EqQPq3v7lDBfe+35caVHhjkOvTB6oN/Cq
ZNa4Qz3dc5LOyVKnwJVo6Ypn/O5noN/wENiJ4WddxTOfIdXqRyIWT6Hu3PUqzxDU
c5RlnNey9dzUwhgtB7bd8UjqKqi84sDyLLry4SfrSfn40skNO7cI+wxyZTlRkcoM
bRsJaQsp2NNOhSzqRYkiCIOwkxVCf97PV2dy25fVxsLp+XakohIpviVUm9F02K47
j0nNH/G9XYNUPJoTbbZFl/bs7R5tA73TqXkIx2Ih4B1xi+QbBAUOcH//KTyr+Yym
uZBzSMdHnzx2dC9QnWLtem9iUEAz+TcDe67pwzbjLyi65JH/zfV5QaB1Jj+K0w1A
DsWNzVIw585r1/WbhXXu9I0EcPn/xpzcXjLmSdCQ/OHIpdlFqTjQVDt7IScElnJS
+nP0MA+Xd8b/9uUQdDhJWyWr84ODgX7/f+NXSg27dsS1oSl64yZT5wvv93++ZJfw
uIyd7QZxrFtCmuzGL5RwQYCo2PoY3u+AEJa9RA3qYkup1rRx+66UG1rScyeY9d1f
0uVVWnUJkJfpaDIxLMRPg/8AxAv+Qivvh0IUb1DowZK+9HJgoPXiAo5XcwPdi4ev
Op70tRD1lkJ7tOuqbZdtslkbYrZ7V3AFQZReVLGnwGZmf0jK2rO/K5TisevZ4/2l
PrW2IIlSSwuC6975DMO1OAL02TUgx55AzSyJIOmf4wcnXMekJ2X4fQKfoEg8qT54
kyhy5t7VXmYqRDUjAvryILbraDxmna1ZkzPCRo8vckAFgshxRhAZUf8mgFfxMuct
4rn6J3GjSF/Xsk/iIChAwj5MGruJ5AiCY2UbX3pJkC/LoIurTqfze4sby2Yn/5jI
g1/g0hAiYXgWaIUCpnUV6luIbq8AXT8wa0D+rVkX1W8Ui0EpjDg2RHDN9SYHFDvO
mAywx3wcz/58AIGWHNcHn7+v7khFBWmDs8CWzoJW6+uJHQ9XaMg9U49+1uZKIefz
EigAPoondKfDzpFW2RZbz//M8QL9uVAho6uWHmshJSx94OM2REnsEGLfJPc0juD3
5mkBGuZA6LAmhb76kJdqYzPKkz/dUQ96A2ZKvnAp52SjtOGWdmyC4uqHY9CdnTeh
jg+fvyfpOwX1jSIzzZ1qoZrXRjdgEm5DfpuXVyoRaMf97+jA7SiQGuXqCVKbpw97
R9rGr87YidF01w1NwfsbhxlhghYjYwjCawOpXEzNlq5r1Hu2dAuwUxZOCoOSgz1A
NVlWxZG0lqYOf+dEfbUXLQqK2bfdjlf6Rxfl0zLGx/d20r2PJaO0kWx4IDFobGXH
tg1d4MIwlLBeFONdgXWTplRanLaA/IHmL/tDgspT7FCy2JM4X1HKhvOqpsG4IPta
YfYQBcOeM2qzXtIHYLljXABLkaA0D6qqDvdEIu0ZUk5PcpikpNNErFTxTrQ67tqp
4bJ/jqtvObgJ74VdbIwe4hFs4sZwUmbKSiu/bU1P2FoBfqtnj1aroSuHyBYP1Sy7
lr7G67VqOfkNnaHVfBq49BQuPuyNkqjRCH2BexWvrs4LLMuvp0zYADTB05u4qUHI
lt24KwhyvIBJHqVHLXa1mZQyYwXU92EG5eZsDoU1wJC70xAhTOgSPWkU9JfWQOXu
ru8KMiTMTjsx/679gOhr8F2lB8KSkS/HLukbHKlGlxTHbJeEgi1+yb+tlwG7Q4EP
2DTSuztdLgpdEsAhtis3scavZ7ikgQUS/SRN1kV143f+F0UhqVRZBV7yeN8vFEzu
tFtWzpacBKx2HVdylwxgkrFc6txViFHLsJrefnSdupXkWcfJIXSB8kY4vw1hSq6h
/MFNqhQMNr0H5sMmww8JQVjVhY8yJxaMpjY9vHGVN/nxt7mtilEsaW4ySvx1h7Kg
XrBELDK85WCo75sG9n3Mp29XVNKKGXVDNB2aKA4m7gheZtNsoNZBDTbYonIkoPKq
7FDx7s8t6jg83u201DcqqJN9nLou03BH9EOR3DGdvBeLdmjsABAkEefzWVSSl4ay
quA2pEnGXKjZIpKBuEbtgEG3BtZeQekyXhHLME2zP8p8HgTf+prWqz0u0VKaO8Ph
7HPagwfnVM5eaSHRxTceTdW+5FRe2QodO0cRI2Ngzp5kv0A1TKY7xDrStcmMcOkJ
RYZ4BcBhMRgFzKg34aerplfXGooYwtYgH/kHv0U6iCxFK9YugUb9y9TFIYkdJn7a
p2M6zO4XjGeA3Pq5ccIuFRKBoyx2AtcNI1Xil5d+45uA7Q4FYGNRi/gvLYbPwJ/V
tkZfIemt0NpAD2kN1ioSLZEZ/hsJ6vfSdmPiScnpkIg9t2B2Y8MQeiVg2vAxjSQR
MVSnioNqwycaQOJhnpOIWg5j9374va0ifJQtHB9sOYEFaD3CHBR5YlpfWIJ79Yqm
mlRNo9M29fpeTqhM50mpAYu1ObANhvgbjor71NCN7vQrAkyHoe3PdqUb+RBSBO+r
D1IBjEpBue1FFAcDRSSgT45VKpX/HHKZyclNMaqySY794uLeinPo10fC+H7zH85x
HLP2YpUZ46UCwv5/pOa1Mdh85uwEXISgnzRl2h3Y2OPv5uNXekFoN664ZXSzatgs
X6wfUMN+bjA3KSUHh5VY4j8KToPnozvn/qlToviMXt+Ax2oUpv77EpKUZZUREBIv
Gn3ZogvinIMaGlm9//K+VnUtjCVjk3bmLjN/IhltqmCfry8DrveGJGVv/Icf7BoT
9o9mxQcg/VWoQD7IECx4S5v6vcshMVX7v82LmbJObZmnszxXCVrvv4GhGSrakMu9
Z4KIhU6tchYKFtInX2zM3+lWooHNsn2Yi/Ufk/DTYoz7OZAkUMAGWTXWszDl/ypS
h5vnIo5c41WC0/riIYPjVgPrv6n+n3OZQXduukhuwLAF3GL11npZNFpqZBmLFBxX
pxWP+bnFjWqr5M9AeY+rhjEKFzRFk+bl3+z09GBxFOH6RGKSHY3QXWdDTCntN1Yd
NJ3FfOG8oqSRg0lL+N7+u7PB9p1U+gGUn1XQQulasIkCUzCXU88FaHr+Vb8sGwNY
8L09IJDvfbLslGz8Jx5RegnXjd3mCI1PMIqBRrMVOqlwc7ZmH/vb89TFKUNMdssz
YY1dP25DMIKdmfVtlr7C11F6RD5EDgpmuNtbhHGXUAXOC6cuQV1L4JU3158LuN+z
TGswyrAi2ILbLEHgM+nA9Fnh2fLZSP11JHcQ/ejPfQoY9OPRg1vLCp7SGLugQP6U
DYCisSPctgYrTWq+vyWTjNf5CyFQu94pAZJNFxgvYNbrbPcPlFtRVmmtjHv+2T7N
XKXjCa9ThBYMUwepcdn2kJBmr0GZxBIDWp8SjXJyjA2bqdrIP96RiKpNUeguEh1+
wYYMGWKZSMPQXtbaV3af2VD1y7XlUSNvSFo5RgE4+k0SLUcZFxTcQVqbJxBc08zs
qthRTcjpvSDF7RBgdtyK54wI52smreMFEtFmcm1TD9UWrX2aOvCrGc4cug0dBDGW
+qp7o+qvTzAp5CLkPaW8S5FcK1eAiDZmxL9BCyGkq4LQ4FRuxbEhHZST7qWfs7JG
p7DM5Zas+IZAmVz90WxAKwEpkIuOHswupHpvHADEJ3r4xTDgIkyjZGzdoX52+KJL
QmpH8qWCtiSv1wUDKbMHQy13m6P0+3IpC8A7R5BEShiqwlvGRtiKUkASKRbpNRZl
dY6/auYkgP6LGprhqc7kw8SDaYYG4dnMJXDZSBfuYmpHwW8NNQ/IIQiKLR+MXGQ9
u5nbz2Ymzhd4mer3KCS6KXoi9x7DAqAurq9JcO6xstdlYRvtrMdbfwnL9M13mNgC
c3puCl9bzM8ccdv5fy4qbZ6NwXRS0mK8Cva9y3nc0RD0mVJFKoboYwu4ELOgWdaA
ZOI0TfEj4cCO9Y7vYZ9Irz1hytq7e33KjpCvJ5UP81DdmW8F2eEz60b8P0Lb2QT6
N4RIybe5STCEfKpAl6y1PBmI6B+8YLGJXkA95sY52q/g0vAky5fQkgcp18zmo9Bo
G5gy6f8FV2qFKS4g1/P3CEkW69ch+DHPjdfm6/Pceh/UVY7qDeoaXsMOEFo1O9ue
U/VASsstYN77jFScrP9u0ADRYRTK1og8luLeayw+ZloSRp42crEa/HS9UYLy9ezb
UPqRkAILenDEFPy/FocP/aaFWjNxuVj7HJsjO6WAd9X0gUriMajZtxj6HFK9ffJF
n3IaipI4OOjYaaeR0FMlLoN3sMnu2fTf6Z0z7Y87wvHmo0VsNBQ71WLMEbe8poAJ
6rueksTu0PIk4aLYGSJBA2nF3zM0er/lBvbsMTxWy8hSVRyzFpChaM1y9e+rknCA
F2MEVwDT9RkE5bWGFjaP+0LUNY3pZt9vndXEw9HXa3poAxLJswmYfeVczoNqURLp
VqIhSYmVL8clTbWG/SFOPUbIice+TRhJPoY8p5desYQpWfqPsnp/ApBBTYLlLBGK
innj/CAigy/1thMl0ZANw3grFh4a5XWm8kZwqqubohyYjUyj6bf8t1KuAbeWBS6o
O3JwflB4DAWuFz85nfqOtZKOiFWEU7YshzpwnoP7wjlN3Ic2e7B5WNd5c6R8Phss
1FyxM+YOV6jsPrz2EOW9y/Olttbxtky6pmte6OpNYU+a5XU/zXs3ZEHWhnXHzpK1
W7h9Ze0fHSwrNBHjQfkKjgLwQDhsXQpKcZVeu5QzL8ur9xPFt/oSnMYFCULXJPIE
eWGQxUAbGHZ89fV9Oa+PsE6bC31zbZY2fxbxp6rKic7ItitE3mBFvQEydBdl+6g+
l6IvnYNmeoc3ZS8mmK76oPgaXWGip8goC5PkYIx75kDoC6kIyDz7uoyN5x5dwNl/
byhKB4rFmN2ccIUZUlpcBuq3ByyDhj69Q+yyff4D/ZFDhuh3hRvXAsMRaW/mWK2/
GANyPIDn3xa4fokihbvw4SJUOotpDzDQDRYZoWF39RZAqXizu3L9zm5UD4RwHb2R
YcZrFZEIUygx1mIOCEV+BVFnbmZEBLUygxedkk0hmr3UwgWXYjvOXBb7vXasZ3CK
6xAKFs+vzV+t8Lt8aRa1q0fVTTOH+Mt2dTMMgnju6qHzol8MRw9+onZn7AjPWaF8
ecKTFZua2km4JbTIDgAQSSolKTxPZBqr/DTdmbiad8pb7KcpPY6of1BsflvqkYgJ
EVWmrZNRDcGAJq+oG3FBt0snxrMQaF3LKJlPSg2FXpVyIuP7Y84gGLceKJND6FQV
MZZhZxiErcX7gsWQqlZVMOcSx5g6JyHf4f/wILL0KZsub67F3EEvdWccWw4xB4Nf
1kFqQxX0RZ2G5bdpVMCQum0XkV/7dJ8Bc4Mhj5dxyc3Ahmds7ATJXgxBHO5JZ7ko
vCxuvYi1S5xJnIWU5y+mu0d0KSEYp4fG48Aq/eHaGROAC3mzOj0F3QLiOQPgW4Zh
POyGKzfIUTzHQ2FM6RQ32dj66AkKS99O2f04lSAG1vDaw5r3nfyCY/WbrDp0lKK6
9Kk2cTLGebAb6ABtQ4ZMfExCacjFjlywFNlEvHXDURoeRarDkDoSrld0Z/T9SVxh
3iRfkx2BtCRuPnqo8F9qqDqmjn+RR137wbbpbvOs9hgypqROzeZh6MqyV1TDlRPY
30awa/mzrqRm/VK2SnFMIZCPeV3mzT984rnGsRh0P4ZQH9lJpfSg2S/v908xA5JU
SIqyHZZlCr8MQW9YAzN+BmbrEHPDGcA8ttQXnDGTS+Q/bHGjt1YKxJ7EzuqLVXeo
QnEEVz2xM0uyx9FlWx5qO0oZYV4ONIye1MFX3bGtwoVUQOolYByFP4quoXn8F/mh
R9v5dv6HYmBkXjULMLEocWXTWEChDtZ/zzolzLEnMSKYA7itEoMRxrWxRLRaAeZ3
WyEBqqNKf+RmofWtiqmmQ8LyDz5VYAcbXc2j7ag7GE0dtOiPqn03+3CfQVjV0Avw
dZ8SEwF/iugqr0j3ab7KFbPW6D+DGCkc081v3yCfwjdnCJzoa+dkL8anBiq676tN
QMpVafqKKk1v3sCqYdWySuarN5KBgipvLf9kGn7kzeiN8is6VMc9EMLD50cuuK+g
BDlZI5MbA4zCd5Wv/0G1zwRYxicTzIqwXK6uMGRq++2eCv3kVuwiJK+0Sghe3ZD9
goslZaSpoh4wZV9QJriEDTqLsMaL1H3AKf9OQizsDd6Jo+HdxHQMP6/tbrKF8SDG
lq3CeZibhB3IzfgzdMkvQszrPAcJAiyBOa+dJugX6vn/TEjYjwuZfLazosGdvat4
6moTkn3rsAhSLyAKfRDl0zaUTP3QjYFV06GrZ0UOW3YGRsMLX46n+PWP3i9K4PiB
QBkSmy28x9iM0GTLuyqvD1l/aLn4DiV88ARWtD7vlsVDorWOdbNgjPXBUPllJ5Xc
njXN6j1cS5Pdjm6wpuUz3y4pfMpvtwCQLrH+OQFrUBJejk3oFqP9L5o51Sios477
h4xotLRsJKgsqc90H5Ib32zEMdeLl7xmxpqsBw5WHSnK+hp8Czy66hJax+9GAWjy
0GEPEnbnEklXLHb7Yz786b8UK2TPqJlFEOl1EJcJdVujMCBt7GSnE+2kwu0gxM2h
jyE8dQ47KJenN3gG/Z8e0D9BoGeQJZieRYLCT6DILKyRC9m6nQ2g2yAM023tfb2z
xopqSenfIe47LBTqvoIVZRrLnzvboqL2HiiPyV9E1L/091K8uVTvyBWsrb9BqqKV
o0a0MIe1D3ASaMMfT8AGRyGgN7mXAA6O8DP8KixPQguVo48vsrEF7ZPbzQa6ldYk
FiFCUHSXuGXc0BXC2V1EMjsXxRcmzAleZj631k4PNK1XdeH2Aree7E/eMxCDJNI/
ju714fE1P4judFXdsSTVNBqEV0cAazcwmMt1iUDI87Ei0n5+WsBJWbiTbRzuS3FP
IvmNBQVpM00dKH7SPSU9SydzyX6PQQ39dTKosO8rx2IvRjJm2YyiwZ2ikuBhRkwL
xWIhTsO0hOnAkxXctlfPu7kFzroXcPu5NrT4fTFasbUKOH7X+HWAAiODFYhqhir7
wteMlJeETCUdTIMhRQ4APtHEtExq7mIfoESVPlzO2ZD1x1Ip9rez95ANsUZx6ml9
ilRzPVmedYXVx0b5fvVvX5HnWdqrYOho7SynAdssuuB5VCzUhtza01Ot9hiYNr8T
9biy44jx6IbsmGXKsvLeVkRnXUhyZbH46YFwyJKYSEkpxMwQf2/YsJ/ekSeaaZvP
SiUm8HGAI4uMK8AZ0O7qHyoXBjn0ULjK5UMCrXB277xf6z+9o1v4ngIYRZERAY+0
EcvmhdITvgs0tYKfARv63Vvv0P5+N7mXXZ4Gy7pvqh+QbttDQgfQFrvGRdR1btkJ
llKJ6WLSpjthHFpOpr4ODH7heVwj8qgeDr2lytErdLvbQ1HcsqvUG5dDaMrp/a5d
rizxd+qs8F+T6J9e2EXVLEBZtcnGWTi0K+pu/UXRXngp24fWh/hbxpkmoaFL4hwZ
Vm1bsbXfCraakLq2a4JfjcyJwjF9yrIID3DP3zmFSlKrsONn14KU6zm0BzYUJr/5
SQoLzKcFlve5KZmWaSnwr5LnY8+lzYS37+paGI2kCrARZfWEB5pb3SA0CjMP7qbn
12Qh3B8OmtJEIEM+CoUhEJ62SAfzkCz/Rmh6dypw4T0XE0txDQE2OKXM9oOxv/oS
tXFS8OBLs0SIR+WOlJ5yG7E9qU57r4ug/3QlpwZ4NzLGiuu0pzICBMM6nsHynsJ1
6HwvESvm30UvD7n0M299cdQ9f7ibJH1l8NUFbynXGV6GpDCK5P1i4V7HeVvNdj85
Av9Dy3GyfaS1cXsMMjWxpdXBOOajU1OuBeUkerxJBu25t+0jSjStOqAtC7jRIo8t
`pragma protect end_protected
