// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 03:56:41 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TLOECHvZf/8PT+HurNJXH7w8lJjaNyH8+7juqQdpiMkOcvA8H27u2hqgiHc8XqRh
A/t7aj/ITfIp7n0gAheiLoFxgFyXEQst8CLDutiFeFXImsZywsL8SyrhPkPU7xCn
ERAN0+LQHCHUlUk6bYezvR1Wm/JN5CSU+WLmaaWSUp8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28016)
mmvk5Gwkkxwl/ApSx1VE/CTV6RR5PuogJJiGSNaSeuj9dRtEmk3JdhT3w21LwivN
zNgMUq6BRhf7kaoHRGREylAj0ai4KTGDsUjAJChilZLRH1E4eKbVifzCWnEgKT8v
QaUCnAYP1iveGktlW1U1nptEGZdcHyENhsvhtpu4Qn08H9SgwB5gvRiGELYil7rd
d/IVoU/zeP1QYdBi3tSM1n/k2R0gNg6281HpAnajtwbK9yPkbAF+qpI3yYZUjQ89
+bjd7F/sLRV5rMDiC2sNS3+BsfxeU5FOV5+z7GPAqsPYBfR/nrMDhPms9JlzDJ31
iGRDfAFtZde0PZxHpgX61qWONc/qNmr2S5Zavo2mz8rNTqf/nuyzuu+znyOL6Sxs
pveYh1+P/Fh4uFRaLx3LD+rd7n+i9843SIe3uDc9Lm23L4G7LBHBAiuN72ZeIbfV
vSdQaeQgLI9k2p0l/Z0GdGsJ1ckhSmNFt3S+FYexzKWIWNNEDzlWX4JNTWND9xAO
0B2V3+rHFF3tvG1XX5a5+ppH+qNqFFxVdKlKcjq9xzYIH6buDW56u8xlcMxfvkxd
kBOZXfJ1AwfABYgikVEUYM1L3EDiyD4H4odXf054Q4qSXA8l68sTe8uN2Qa6U4vH
cUmxIdGHcOMKAJ1uXNYJPJSDIBNI8zob3ZeSJHi0jmcGoa06x189WmrZrOpB3105
0AbDc3ac3K6pPWOThdX8aaPgn/sMkNqWM9QirMlwJpNzvkLjAzNVOSaKH/iLAOaP
ykTVqgkDQb20A0deXbb0RdIBsQKxHnN1X8N0j6RytXgB87op9R7I13xrRgjWJGmV
sczAc6MCz3jJp6gdcnrI5nJdWwMpjEL5psXeo58B2/BGDQR+S/4A8+wYe1ZWVA5y
7QhzB6POaPkW8UEOwxPGtkezMSC5Z87oXfu6eprJnXhqcuS38/V5mufkQZFh8ki6
6loUUPhQSwNyeHnruzwmzSuVnUIBIJapsMWxO0R5ayS1/o7vaUl21qhIwfXwjCG9
0+GIaNxHVaFyrY2OP7wkfH1uC67PXsHuHIArqt+6etTZwamhlI7bjNp8i221p0aq
q+i9nfHPxRMdEpSZcCVUrC4LrUPazvcj3LQqyIR4fB5deK+Rd/P8BcKJKW5kutNc
3DNRM+TmKi7gl5GCtciIBZBzHVYmOk4F8QWaVxC+u6Si+rimtbwgDTgk/qkacc6b
622rcWC9ZpKEffd+q/mwymkzWzESjzEUrtrMNN1sQ2WpePRhEPDg4Ghwttv/OBDa
L6YuD9H20fod77SH6jqBw9olUx0opyt4H+S7ZYYa1JtfIOvScFLS0KfZLNl+abZb
+P0IXlIkTjt3eHT5m8/5dDPmj1SNth9z0PRR1K6lu+hLBV0ImsaM5uU18RvWN+dT
oLSBB3s6qsBST5s+9weae/T6LNLq0r3D/srWWGTuBuBRmi6rKZ/ffOUO0OeTeHfS
oE0HBFHeq0788cTaJ7Y585rhwEA5eeO0hiZiJtt8kPoQ7NBuUFDhQjzob6wcElNm
wYNkuAokPygNOwia9mSuiQYZv7Id7RIticUTvRcXZIUViNNsuzzFPYfIqHDt1hM2
YUYNTG/CQSjsCna2gkq6XP+HMcWJIDT99ftXhQ8c7abc5vsF13G6ilQT+Q+64A/l
MwIdINz5UpIigDqfr6a8/OeT49hBBbCCCg4nbdUk0Dbg1/14oHyc0pcxf+M5kuEj
oWqjxq9e/TiVX0O6wjG8lkXXUmJcOglVfcVZv0ExhgaGMxqTyiwsvdM3KEUaHIvB
Mrgb2TpiLVOT+Jb+wWByPcWkjXnHsA1+FQF3yz+2ElYSFCXAJzWjFRYaSNefliA5
kspRaELFTG8mWG7FydOXslrqMruvmTC6Wh+a9MyBLuDSvXh7xScLp7raiYwL925v
HONhZNTKjYfTgvtw23E5RMLiEsMcbhkmcWixBHvwUNajFFPq0/r0uhmZKzb7DTHF
7xQKWx2pa/+0JBoS8Q3ZOGDPWKVl5SxRHknt8g3J/v+AVgj04q3TZeCJehf5hbCx
bbUpKn0yiRjnvM3LxZttf8wjVxRDWYxHWwaDgxLql32KL67PlXj2w+9p1je+mgrz
4Ce+nTkAzi9Njdto36CkTpF/jqCoBMLTw+GfLuOmEVHpktNDJHSwaXyTgVBJ9/bh
EKMfW+EImq8QAzATlOtKMgP+1YDzYTuW2X5saKKFPr1aD/hYOgEs+wq2XHUw4Nkz
6Gnkxe4Af8Y1dCrGMZparGHeQy6u3/QbpNPRaTEf//7UKGNfJj39fyxFP19BvFRL
1vELgu+hwYiaM/8VjHP8xvY07+8FEr8+oNmAJju+8zWSuFyGzA5BhjTKNEa3lVEI
2ldu1Bi5h1+/j7EsMToTN1UTm8QUtGhvt8qqvjfzNjMYrClWSmuazlzKgpz6skCz
WA4cMYxIRm8WsWkr6eoEZy/eZWvzoIxBCpBQMBetjtNDPI1soOOPPce3sAMOhWqs
bqan/iuRljcNkf8hYNPHoJ9cxAdSVPiwzdeeFGhyZ/N+w+Ltv4NfSNvzZ5nClLry
GMQSmgVqqw3maG3Ic9r2uFCx1SujGIkuTZrzJxxRot8j2RiPnxaZX+WGzlUYADoS
GrNJXAGkoliJSuL0ueVGbXnXlTlEnv49r8BifjwWFnqYQf2UOcPWK6mtlKpyHhAK
pVlEX47eomTDWaa0RWLCphpE1BKuh0g4mXFLbhGaEzDttfnMS9ugx5BwRBMiDwBp
lkYdbfSFzrFz3IWlvXjGiw2W4IrkxLj0aag7jg/njTQC0IR6RZ6Vmg5sgYCVwBWj
98IjBmmvWBQq4qkNCWHaadyTvTXn4Y9f1wclQpWooQ6zUv9VW2RJDfveL04d8XZC
yyy6Bv7IKiudLfsfL1l0CF21RKBqpXbCqnNyDFgsjCH+8LTKpP8DwY/XPN9+yrVz
/hbCPzz4xD0SI3k2n/pmierPnuyDA9+/YqN2Jf4J382XO1USPo/DR3dIXjBGAKkj
ryXZJbSB7gjAi8aLQN3jFpbA8v40xO5jtWlRgk8oYl5A8BRxCcK8xyffbnLP0kqU
VJ7gu+l2U9CBSUmy63+mqONEBZQqNQ//dvsrhBGVpbKPaluczutiwk5K0aQg8ObO
Tx4ioIacwOmrrB9gxn/XmQyjsJq+x/e9UIA9GDLKmtr51BRYExtw9enBSt3/WRhm
FLbOjcF3tGep7htIzFav23mYeyB2V5pIPt021l90xZGjscUlx22YNahPVL6ctQMc
+X2h+/XeLRvJ0fLwLSZ/mBqDs+ohq7pxqVRbEFsQmKLiSBT7TyFOsnKo6Kfjk78x
jzFHtOUFBd4zj00iYoiXusGfiftKCk2y+4QMEuyRBrtojzrtM3AlHDR7lJyiik31
c0mbeKEKcF+2G1Fv/aKxL+s5f3C71BeyuDYtPFh0n6X5ETEuNi1dzjTAd/JTFbD0
rcUACd3lBQ+GK5h2KhexxjUiOF3hptWZ7L98pDkRb8XZPi7EVp9g3rSEQ0q1SVam
U/5DC79q+rWTMUy41I6KHHNLTL6INxfTcs6JQkq2XSfNDGJ2/+GPmQ6Dyh6Ibkol
wYVcHKkz71Yaht3fwUON+Vmw+XziBoBwMUO+o6loeqMKTpPyBOOObIGbR44WVMKr
GLNZgJ8mGgsR5ldd6KmVuJ0YUcdl6hdJuzmJrPgBGFdJyYwIIs1KnfQxkEmVY6gh
p2ZoDRvEtMj1BkzAZxzAl1VUcBFr6yEy/a199kYQBHn/z8ABPHH2PNPhlzJbHHXq
i+mkT4BzyNC0rgGMM14836Roz4VOw4fLkIzJ5YdUA0Fd3JtTeQXPSwruoN8ihisB
NlIOeXO0Ho8JAcGBZxRHMsPy6RFlicf8HMQUU80TWLH09Mkl2Fq6TSklBYscXp9L
RQuf74Jv0dFW9YeNrCAPmR6P97kxXOZJU5+kJvIS0taM5iDiEI+n1nSItk950tjr
yDKmPS1Qz2O2ttIANkuxRirVOm0jcUeBL5b6vS8zahvbYvf2ONYWj5lKOrWJyp1U
EHwjpSiiEZqw+ZmJd/lEIRYr3pPcs+Wc+P+NfsJNPkKnXJ6FzYpTnGX/Tu2Qf7MM
L1gVaxHU7xBcX1U3ZI/WWJUvfDqWdStODRynDHLCOFta4wSihIQ+grxo53piN9LB
mfg79aDmznz7aXRT+S+RxsMy3Y/tffganLJK/77IUP7ICMGN90nNA7Ol9i8WoliE
J9Go5zXIDnmdZE2nYUGiseIjwL5C4TrOf8X/vhhYgeZLdTaIpSS56fV+K0XCh67Y
XJPjWo2uH5o01iCOs00iS2Q1Tmf3jb9CjX5/m/7KKr4CG05kPZxp0QFwTZYFZej8
jHl/xD12O4wS4nsfXxgbojT7nAABnOK+10TRzijGyHmC0SWLaqfMEAmH98+/4N+H
bl6cD1CaBcRkuMl0ElRhCzUugPWYQbmehT1xF2qyrLmXCODz1r8m6D1euTFoD7P0
XkbN+cz2TQKfaT319vM0b/ysrJBaUrPEnuVsRVLas+qUw5I/MR0Dyrf8/bLegjja
LAR/sckIDsbhaMYOuR9B0WV8CuNk4anCqctWjhlgL0I0BuJX/vAs9P0RALszBYix
JGmKq7SToDlpmUXWuh1X9OEKAb0fsFq5avAxcNLMnm328P3P75VoqHRc7DVocP8v
ZXQGfE3kQF1q/+WPWTzbP3cH/zh401+51UWo7T28SkNTlOmZEXvHhBWv6dbPny2D
pPN9hBqocFZ5pBmT5aGScjz+NjN7kzvsAYZrAq1LQ2O5RACeA74pMvgVOVIm4ssE
iCrHItve2yLnhkaGagow/NFC54yvJfFbkzqLnWzElWGuEDLfydt1DeiF4oSVUETv
RJH0QPEJEO+OZLz8+QM43ahWRXYXTnRH7ctD2XMdu75NYYxeFNRGRftLEdZLRGyp
1gO2/FeVAeF9cdPa7aQCo5u44qHzEJXD+eDXIrc7E2CQl4Ic5PiPSHecp2RtAMS7
vV4JcYNU9eUfAt0p8iS3HdwL6aPoM/MYUj+wYtV3oeV4KlOwPblAbHKRhcj4ckRH
2OR7GaX5MeeEQ1laiFoFyWGE0cQUzULEE1yOiVN6lle2y0wKH5gMvlUJYSH5hH/5
jLGVbsdd2CDc/t48A3n0Ep9QG9BfxWHRvlfMWz8jw/uArsYnjBNDiMfZdXx/res8
RGf/kLCge9Tnd6Lu150xXFNFt6g7gNtLuyITx7ya5UcxTJkHcGOGtDk3YRM6dML5
qalMxh4iJr3cffySPGttGHF1fwXTX6ztUHyKhuBsyF74L9pFZADzYy55HxfLpezq
xqrOtDSOnuBfQU1jx4bbP5kbuivqdU1wviGGNd2yKhQksYj105em88kidPj5zp1E
JVhYQ8MUTHCg1XEEx5MUBwbph/S7QUYF8mZ7NMwcVCCVtzWyJIdf20VrDYSp8TQD
R7aqEKPiImbkPJwM7zxpdGYpjHGsohKOr79ocfQZI6A/KX9P479me8FuBFuOpk3B
H7ISEfuk9/YiofUXS7vvvZuHIofHtSgNGC/7S/jiSTv3Yw+/7dF0HQ5gSpJk/9Ml
O3ytswq95nCn4nZkFSUBZ/zgLNnTdX8eD0O+6BSwQnmFxQ7WBPlW9WyhFtehyvS7
DPSMC0QG3uRzYU7eQx+ZscdiBYEXriNhl0LoUfRPswyB77CWd4jn4jvgSvafHeS+
zlWArhE/cfPlnr0jx3anX9+pFJTtYo1gUcKkOMALOOwDqlEoTjOsh9f0NplvsCjf
EuBtTvCAfpztJUnQuiLbi7ydIrL31TUNDFWadlm4ChslBIFNGX/NUmbMShr/pkPn
9Wliro2BgjAGLQsXgl6191SijqwbxAfrm9BEPN7vsAkP2wZL+OU4dEdWc5BWauJE
iRxNqNVOlvnddWLJ1EEE2Hj1SngBjMvNFBZTcRA85fEpKJap8zh6KTTO9NuBNKfX
lNosUjrlON/hwxv2+fQUoPC+TaW7DzIFw+Ne1iwgUl3zGyZOUHcGpL7PAlilg904
gi4H3mffk9GtX7cJXgAwvPwbQvBiKpc9TlNf3b2KAfRWfr0fXQ2IgKnvJU/fToKp
JUmYECso3dyGePFaMxcT3r9MDSmZ/MLaqq1+NmTqQ0FEHh7WR9KsNR3zEMOpCfzM
fxmsRp9agkl7Q1GHKaVbRwrCRRLH7rTxkzpd4kI1pDdWS9zL4AfTrvpfSXiIz4KB
kNYgt946+sCBesa/2ax0ndGUyRx9nedAButAymSdIui4VD7eP7wbuoMmvP7gdPKm
Y5V6TubZ6CUctQX7/Grm1guns/UCBPnMnWnPMf1QTG9sZYLmccKEw+0XazG2E2l+
FePCK6cSTqpSI3YARbsy9od8cwzlmx5FQjix04Kq07WPSg3l/l4tgA2h8/NUssLK
6nlWu5vMCIBs1iOEjqKD7d3GsB7/i+oRYefu0iW5g4R33hX7YwFaZFL1zZueQE4D
UlZzOCkqg3WEBW8WGRNIU43N2Os/0fTFMtyxRcGa6Bcc197nsumJEYbavU2rMcbe
1eZyFicTsezxZvoqRuEvDgnazl5QT+/v0023g/2MdWY9W9EknXbJRFdB5Wvh0x8+
C/ilL3HGpvvtwHUMe8YbaQDRgzeN53DMhTb8ZtrwUu2Ov32/rC0ReMrZAsbixK9K
mX5LKYM6ouKKeAC233QhvkmlQ93YR5rpg7M1rOv5nOGruN4Tkti2TROCMiNf3qPJ
u7sU8nhngrb7AK4xUWZf6NTXnd5UrbrmVi/O4Mc3Kh0rY+b/jfOf4UTHf49mT3g6
sw1D/HaKIeQHGFmVs8BBF8d0OWm1lUZ4gOIswgXs2ZJJMnQJy67KrwBS8967lYkw
V/J3pB7V1X5fwSfUsisJUdG+19DptgYiJJ8Oa8894UkmeQdKbScpeoc3Z5ooepwU
zEeL+4QjtXe9kn9DIICu0F8aDTlo3f/BiBu5dqgimtoRxR1OD/Wk6TBaCwOoFrP6
D5jL+O40TtS9WknIae2Vt7k+Ae0p9ILXhqFCZ1cB3SDnzPh7tN4DqykYNAf7GNOJ
jq/7xrT4N3NwS6TM5eqk5BeAYh1ryJBqJsDf9grh2JhfqGibZyql6gBLopH8UO+v
4cTahNXQlP0EEaQzN2RNre1wJhSkwy8vIsHQCBIIbT3orVLNGiPvOHRZI6fcATsz
OY/GxTASvei7duptAmFLcZePOUTtl2eM75dfVLBj3i9NoxLpCeIy2Aq40H0IGDpk
JgOQLu+qfTPK4+jWt9GebU16bZN0erVNyojmgZGSzM8ZQ/ZxttuICUJD3HjW1wCO
VoUV+3trxGQkYwwmSsRHlGCRYQDkvwkuQCaGO+gLRERO5m2rb+lHm1gWn3tufx5c
3aYk5gPkN0yOZKmx8jCowlzG8cN+kgdUQwvx/qTVK6kASOaPamxsrQpx/X7Kmyws
S5OdYhr7yX+4BqdKlj4B3Ge4Rn21SeB+MFft9i0WI3TJDbt4FGd4eojnXsvVqYf5
NMpA0b4EUhE1jgLc0Lz0YZAijqyZA8O1CzIUSIi1y8KPGvTL2M77jA3b90RqR7md
8lyXDdX8uDYCys6UygUyv1/htb34Oinb/4J2iTc3KOjPmq17IT1npfoicyDxggMP
5o2Pi1GUo73Q77DkMzT+DLoGmuv6Vj5MWpj1g/suAUG7tj75zPuK5eWAxA4ziAWm
k0EN3XTaotxTDlcfZQElp/7yN1DwtlT1jj/ORZPHobb4P/pamV8/0IFupObzeNwg
PVXIAZkWou8+v1DL4sMd0eVxl8gtAF9i9ZXE6CavouUdDkK9SzacPJYzXsJs5lRD
VQDrp3h5eXWXVvlAiylO6/OaPznpz/SUPeP54xIl09vtPqi4mqXskWNvrlHkRm0w
pyXMFQ6xAlTFYLJtsMNmjv6hvZZ/seMZhPNZDZcIXL6R6zwtHVpCPzIRQYGERjvP
R8qHf0JGb+AgUh2+RsDyctSkds6/VJqjcysA5rXnXwPmqh0jJyVLZF710xM3GfNn
9yUOzCGTUVfMFXFPRJJyUvn94ckY6riLjEdAtKhKle+TD0Zf+qweWK+HX3ULfqu7
Qo1oVq1n+nm2kYPV+gYOK8rAWdaxyDsQdFkdJDB+040CjjfGpe5cJocKtPCVqjwl
xB4QYJixxGnsg4Ek1L3XC0flsDSU8ZL6Y+EoS/C+LJc5bf/QPi0aqDeevf1J2FFi
LNbcyI4OmkrW43xm+in0tgWyJi9tA7W5KHfmn5xoddBEHydlhvXa7B/yhsIHbJbZ
e/KUH7cBYVRF/rp0CYL1mEDcJn56qwvtm3ZvWOqIbmdiyg0lIewq6LlBfzGgkKyu
MuZyrYsP4cfOLsJoJje5MD/IBmGjhIDT4TY0JCV4g9qEpiNU2GRQW88pwZGBmkAT
kwA1UGV/cZRYtcfptIcD3zNrEf3UjOw6W/sUkgc9MHKyqQWDDK/gpSqMaocEs6Co
1dwnY8SR5SzYC7OdI/aBw4JUM/KHtGG7vkq7dDFe3/YDArOA9Xbece3DVZIFvZru
IRN7zoWdUDkuoEKdK3FFNwnqXxW+fA5t5aO8HJiCdyU3xnusV5cEbewTyNQDIp7p
8zXk90vOhGP5nr5h7vhtGwZ25CSNTXkzLq4AX4s2k2NJL4RvvVlkD+Txk339hNp1
MZCAQ/LH4uh1nBl3Vmfbcw1+FkaFM003LS6b1if/fZTBWR+lIGvZRt3tjyxz5Dwj
+r0HXrtk71Dj62tVSFLyb3jN53o3PK7KbTtgc7Ab0AdYylx7/KL/7ZXENJ9vVe5Y
AIXpHX7/kIp0cjj2vACoEO3fDJGU7N7PfNmpicnLbGGZzivwRv247LSt4QSruY8v
6WdiXWiMPsDb7JDjAOYCHYs273YwEeB/BLd+q5wHOkNU28ADu24J6WMRAbAIN+7g
c+Q2j/yk5bolfRhZWAUqGuqvGVM7HF3T68SGbjfhNdoBQDe6/pfny1yp6cnIHOSc
nRmKMLFfaq6GCCsnJXWTJZqEp5z/bNgi4/y+TurD57Z8yABk+Wgv4re/dhgK5fjM
aljG0yxoih9a7z9fOD/j1Fq8Sl4Wx2JyMHzFcRAk8wsUTbZR6ij/QjSllE00zGEq
PSjTzkcyqVNKdLQr6cVKMGbSpOn0d6TDU/mMM8LX2Frlv7hx/QFcXws/xurALPD2
3nODHe4FpPmuJgMtuC1E2nkSxDE8VOb8GN+LH0Tp1gZmCl0iDeiRuvcld6uhot9V
KJmRct9n6KNIPgooC2CLDCUdxENDV2Lkid5yG024+oo7xaoIhXP5tS7kqVod4O7h
dBPjegB4i+4np+CQpkrz5RGJRSsGXSuN/ZV3FSItBf5ESlT76JNKSsEib//H430q
87bud/7EQRDEUm2jXT8hEzUgb5rCmyXA3xUiS4v3Jei5A60farBb1g229VEk4p/Q
b+eqYmBDysiCchWzP3KG0jXeelsuAFEcgiDWQ/FPR7oqYySTIUgGX72wnIRs33iI
5OnQPzadeQWpRSHFpb/V3DgeOt806wAvMPSOijsR0Qj83CdcKG6CBAan7z9z9wof
AUs2DLR+ePQ9thvExtwUGypXzBcg41jIuAR5qB91Gm32wk5yAWUgakq+iFAygE2d
nOaxtRXi3mX6AVNWjswDxse92K2Omd0h+/85mTGTvgFw/9jvxyPI/alNfeQP8C3I
lIXemBqA6+QFGuonpDk1OW9d5nOF+br4AgXkqM7y+/phNJeA3s/Ac19Dvkvsh2aI
fRBSGRGik0992Ges0/mRmYtHNvZgEJoy6KMHnrMIxNpLYK8B9Nm3/HLYhNuVEHaa
WccZH2L4si2cb50gARokCA46oMPjB/E99BAOY2iAB+odi07io/DVH3JRSM9zt808
IQSSB3Dryv1/ji58cjEvbU3ObRa/TmsueHUaj72/wWKND5zkCMYOYAHd71ZOvr9c
/Yu9veWjCoGLHFTjRdSOIqvNLgDJ9xERzKK86hFC9+cAmN0opdrABFldPNO92a8r
MRpuhQMG8amFyIUASvE3U1h+WpBVinnMpPIyLorV0xn08Sd/rXXR6fX7dTpZIGeS
bMe4Im5ea7sf7VyooFMMm3wkkXmqQ8YGrVMUrUjs7W1sCHqB9jQfQIavUIma1UpO
ybqOoEbsn0/Ai+vdhIoIG5RzCF5w4qnJAD/FgbichyenNmEGUubUTBiMY3T5L0rZ
JBqLVz3jpw5LTa00BT4C38lSzGEMcZdDavkNu/+0QSbCM3b7G2eaveKrE7kajAHr
vbsNv6bqFTOtbmFAISYu1JUzW4ey2N3nfh4BgfUcSKJPP5U0WmReLbBOTmHIPtSw
8lc/yaCGxMBjfFrJPLvpmhqFyMobJ7XMpGMeLKb5vvd7+LX1H7hLQCn/kYLGizQI
Z3OV5RNsj+8NTpvd7FQGCBrBpsn6RAkcNJdJ3k5N7B/f2B209HKjj+3euuYNpQ76
PAowv0ERXU5A6IQafGV2QS35fNIopx0DtaeKFO9DVy7syWNiV1rbWeuG17KPobmN
0+r7KVSSAOdYDJCVk+9g0D7Cks71rzqo2D0HC1B3Lzx3aJpOW0y5icOl0HCRvN7K
ak5NXI9J+GgFzKIHrP1792Gst5BmPAT1DVvDZxM6yYm8rr8R5yVSh2nKZbP5Jswp
b/EJXcjn1Icrl/xAD0IUIaJNDuwHwqig4YBNG6tPE0q2TwbkKfg+UoqTAYNCQQ1+
sf3JTW2ksZhMjfgTRA+HUWjRXhvSnzSnj+/JT7cDbFiDejpnIhEJRI3SlTXHmBfX
8JGvqiC31FIxFAyls1XBSR4RuzA0TTGs0HT6fNmyfZmDXBgTcRyxtoc1k4xCrfJ8
12Hc0IMaf+RN8IrVDjaIVeO1SB7Hp/4Cw+FcmW64Gqdr+685vLYeuwAHY+vlJIOR
AfLQJRMpoHnwVeIAGrjhkL78Ti8uFI8j1B2KL2V6UtDsDuME4pvj7fWxoVjT5/Vt
x1upNHXh13AtMEdjH4XOpABxD8f0bcTA6SZXRLPTAsRasmqTbq62ZevsOzYVIY0J
Zp8zn3yhnnodOG3boThz22m3mQThx9G+bWLVeBiqG03rMlX1Vd8mFE5AQKFZu1hk
E3LkgZzzfxNlcutQ8IppGt3bF0kdsxkJGvWVkVFuKYGtdMgCBMJhIpeW/DyPzCLq
s0ywxH3/C7ROUTptD6IxdhwoZVlLZDpTdZwpLQYDWW3A7nHIA23QlHm1tLBX3XPV
oid+YHVlsW/T/vhKwqM896APbOMENBRGEmqm01h+lXlKIP6zWm+heFyuQVObroZT
D6L+Iv/RLu5VgHDw9xUkS5wdWVRjJstIDaBnvTcDZ3kB2gVRhA/umObaFzHb3pYl
TCtURGcbkD2xbRLVP+QAlE+VOjoeOSynVmmdc1b4ge1HUnPW7sIz3tcoc9kY01nE
mKe4nv0cyOXmpNoapPCGu8Cg1TCO3Tz1pmsKRDbCBecU2ZWMvL0FQsmt7g4gmVsk
EZv9JDKumIoa8kqmlPSFWG7V4MvwrA4Qy5Qh7agJw4vgT1KVxqVihsk9z2uMQZf7
N5x/HJOVrE4G3AdHjw7QrbqcC1YE3ePvMZttL6bWuyNGtoZ5zfgEZGCqrtXWo3fR
4DlqrURyRAGOf8mSMPXXiT3bN/atNUmzKG86f/gHo0qG1dNuTy0oQaw6naLB5z0k
yXH9WiJVaPfngNPi8RJkbQKSmvSAss8DD1Fo33eCAGVxrDeoZ5IsejFw2WkA/qu/
tkQ9to/3nrTEcE9qF5OiX5pmNZWmLOnonFTr+OWOJsJ/6rpDI2ILttkRPswBubem
INmR52jXEEctCeoZmRZm0IdPtXwE638hxtF3MhlF1Y6zlBcNmkX1fhegW9UYKxh7
qIUDf7DiEAFZYLlPmyyuyEdvMWvT7leGdKTv4tEdv8P8fbv5JBptUH6uJmnUdtCO
gKwfMacygUiWWvtGgYOweX77BIvR7ZPiyercKDKf+9cwbQOxMeMaY7dcs+sLi32y
4vYPWAEQlHlNVQVEtCv4uyrXbCir51YYNUk6QsuGuW5RpbFUHvP9YUiholjMCSzI
IM/8DnIu1w+Gjpd2wS06qRGY4IwJLONXzJxkubqf8jUtB/6wRicI42pL1l/HM6Hn
97fGmNuGMJTDJQPQX9LgZn97oBuQenSVkUq3DcSRIQOrdko5bSR0/9xElpSS/w09
74AZpQspRYqD0dex+jZTG1h6UNaB34P+Ep5uxJf+ldA4N7ikYWt0cMN0UYV66Hjk
f1vc/p7tYIfakfkfSoRDhe+Iv78P2wtY8byOidd7RzVHYHhux/IkNBs3IPUV9OPp
fshzDeIEIUSnFDfG4HPS4DJ6wnMbSSxtcO3QUSj91vfxNBWPGsGd+wwxnP1WyJIh
iqihL4aYwkMvM4fE+yzNJj1NNFNHjY+zG/rLHipWydT6m72CRCM3uqqkRATAkEJe
UMRP+Gr7W1yhBr6hGhAySYLPW/2tP3Y5FdwKPZccoyoJRaqhP5xoj32FnZTPuUZs
TxrUgWCp9eH1iEKz0PNkMeqhMlGU4KzeZE4bFa8vp6olKtq1MNgJVpSpG5MYsb5h
oZrO+osXLLttZdu048S6saKXN3z3+1rI+vLMgg0wSKV2CPhJjsgjFALuocNtk8FO
588faRN3QibDSyAYdMI1skQLQskDy5b/V/MAi6sybSXwLqztM27LAgG2ZQ3JSVo7
Wu3Cvc5Vw4qJCutu7beWn7Ka8SQbKqtKfzwhKiUsNy/4QXWGycs/BrpFFDK/HfT1
aJmMsHjgHGv7n6fUafzLodIBgThhgX5z6tyY4Cytyj9ebrQv2VjXNJ+om/HgE2dS
gvmrLcpkQk1VAUzcg5x5WWrJVzqQoZRdYPZ4koX1c3bz0YOYBvV1ToHwqtYMm6ws
/qVZnzEnuV+8ln/JxZIXoQT7/UKp/El/IENuySu4L+Jc5egO4hOjbNr7cD70ywnc
XGz39UeqGrn2OdBXMDcJGzH5MZwSb3BX55XwCPSO6Y9fWYpi1ouqiA+GWvf/4GWV
9M4EqrjwSCjzZQql7egL3LWPUh2ne66X9lGar5Tbzo2kIkFwlzzlhRANENn3TKwy
Y2heOQ38e0sN4EoSoTmw2Vp6r3WB09gtZ5yMlkAGzESkPfsL+QaZGR8rzEQKAYH6
jFtdPou395Kw54Hz96GMjftlJyqiE/d9ibrFE06TQSDES/L8V2n8823xxSKD8KeH
XBtjT32D60RPmaO6a4X7v7XPDybgjR/EjwHjEibC+mMN7A03SrsUcFVgz3igxa5R
LeE86lKGqeB39U0ismu26JwGVzR8CgJ/12NJv9z7zk0kB7o25ldsQ0F0yXCCXRvT
YpblZX1roOUHXvsfh7JGG+pyzFeEDso9XKjZkkrMhfiJ8jisS3jsh1g/v12nnW0g
hcDdl3P+Lf8UGeJUdf+1UVgX26YRwG4lyZ0grVet9TOC3gAf+dhaBbhn2NzmB+Uj
QEAKvt3x/YRNk4sGUJvIz4gkmdp8ELG6pbxGZBH0t05f7QDQxfS7DpdxlTNf+T9r
9W69RQUFOMlVEkTiuIxZgPpRPW+7sIl0xW2ej970hqMPO8qmwjQo5UAFC/l9m0Ok
ro/LjepgTydSbORtgtGvvhGeIi0tLIupWsZW9UMgQv1BJo2cYfSrUBJP6+pXVtJe
G6YzyA3j7+1C3esFSqj4yd7kQlQqgweaN2SoleLQSJDg7fgvMgL0spB+Ocl5Y+lX
YSEYfZUGhF2SKEo1n8u0vKIK+zz2QO7Ftq2wVrasxn18yFLRrH9sM6w36H2dcX+t
svlFPsOqr7zsrSWRFQ7AeQMzMuoDpITP556vUnZVb4GdUyrf5EnNzH9/CM1VnSaZ
x7FrodpYd6uPRo9KBFb/el3ug01bVEKfs04XZFrNz4sWF4dHx+vfvDMdidZw/CV6
WxejQCIeiq2zBppJJlBG+GRj1Le9mnCkgnRWovpLrGZjXVU9PWOv/GkXWyx2TsU8
YFWXZisQagStmkMU5lyb5efFe2mWNcsTs/JkCzsfonG0ULTgJUGmEmMni6wIF2Ob
PPrUaJuOGkXFZAweMdT1gW5MEVln5+wN63lJlJHViVzj35xKvhKAvzUpB576CCcA
Qchm2VP9l48klPavZyCvgAaSuhFdQcU9SHO/CxbemmGiDXbqK4Se1PBCgES8hk7s
7CclTL+xyqdlwqqwdk6sbKlM5Bb6C7T6kFWDf0mVklIeC6a7/C8nekC3LSR4088u
S0ylxGXSU6uXHi8ACemTZPisYww87pVXGNLMyvj/m0TgIfp987nxYJ1FjGU+JWyR
L+sAXjxAfzAQ8QgtFqZ4WjN5XBblvuN27SOv2fATroKGyxoxmGRGyGPqLuiagJVD
wIG9+whwvgaDFFkxs8GqJcE9Zsl9VuJ74QiU/z9YvPQUlBFWgfyD0pudGlycdLp0
KkDIf0cfjU4Trpr/rRWiUZvvUlGGyxXm+Bz+6gAx/JeCX6i5oaHEq5XgJSZ0TmcK
ubxEdVhT4qHeePFsdwEGChCuT6Fs+PD04jQdUk6B0W36ywGkW8OLPsn7e1bO3PWe
u800l67pksByBnY3Fjng86HmnZXuzuOzPdqecc8QjkK3U7bAucxHsv8OUaofm29K
zjsrGmN6jJXOesiahVf5unw0HqzislFSpbEJLvwJiJmLLwKnkpPz8rCmHoU75KfK
bVRBNKvV6wV2aD4s3lmliJJWcTqmZadSsQWc1bhpzxSCRszC/EdYzuPsgbewtBBe
fvsQYPL/QdzAHBxGFU4vZZrKw4Pz5GCY3au7S31LbK39+aVq0yGpK6Bkqx/kNqVg
sgqP+Mh21yDrc3bPx1RZpiDbh6o+ejsblQ/rXFM2v/y/N/bCWr6NXRdgBOPCn+/r
PzfpItwDJs1YZyPbhy1eSUxxiyMxXKucESUOFXlIO8ctF/pMeKlsuelvG9cD3q6z
u9tat3kzChHHTF1niz/aM+qXA9HLbu9f5lUMeEkQuJukQfHkbaoAYPdKGyfsAR1S
gZxtVP9BkTPpO83gyXx28fz4o+YQIq0A629kHBUf5VXT/MLqU1Y3NdhLThye+mcb
mF5MYlet7OwmeNVWOPp32J0zVjbgfL6+J2e0bl4C6wf3Y5uceOxrk7kzGI6DsPPZ
j+ugJQ3U3mMcGXLZhSQFCpfbmX5eUzxmciQgHXHuvvO4xyG8o3GYKKRM9GTO2IfD
deG2f9HN4k4pAnRVho/qnx9E29665Q9O6keXOl9drgvpDfPhLAFapodKwW6MC4XH
WYH+JjWG659tS5k7tbwH7xZ0wtgktkJxiogPRYeX3uSQOUstQ/dWmivsY/2s1waZ
8iwGQbCjUiVW8WCl+V5454ncDTQf6eWfo1XXaYygbQtlXqdUkRGxTnjF43J94KTn
sGFaRn/F8YK9PYv5DFVDn1loJjk33pywmT6rfNr0rrO8uGjUfxsReLi1a9bYHmgd
ARcYT8oQwb5MjpzFjfAiLAti1Bwn/rJfw2bKP2h+D4JBFXBE3BoM7Mi4mrlda2Vz
HW/kbwT3fFRvX1XCQZVx3VQIJUocUEz7DeILqbgWMYJt5cZMgpZUnDI+uDpI7ysl
ferUB6MlHU+pps9QUvashKDTm7BLBmGRUlwhPNYFiXmM7Wwf8P0w9K0KwTTk1h2q
YrUZV+eKHMPqyU9898Wh82OI40Uo3X0zPhlJ98pVuG/H7f/aFJB1+9B6zo+nLbRd
OvGuB3cxyvOiDJhNT82FbI4fcs7fpxBOMaHSkeNvZ9dGQtiUDzX+S+lBc7yvBJEN
A4eTJUlI6gclR8gKZXDxvfHhWjH7zl9hBT01GEkW8DsuP+4sv4Qw1PvCalsPwPNg
3wH7qscfylQ7bXFX809MGb8tHT0/AY+rQBB/2slDOnR0HoZH+wca3bRWfpnQRcqA
beiRbMO4I5cpA2BDlS+oi4tpC0lJIj3Zsgd6vGGdgRU28FAsThKUQFac0uTfm3dr
IppVVqeH+dW3r2AdGlcnBL5dXB2PEOSZltj4+f33WZ4JYZU0wM/guN1iEaccddAg
/TxQQpkYyODBnFm3MGzARDTbh8OWmBPk0BB6c8VJii9fExplsOF68RgN1Knj1Z2p
xrpg3j3eYmb0pFrGLiWKwOppVTdYIXpJ7GSaaEhbgcVvDgfh0iS6CdrklCiKS8UT
Oqc+JQ32SNRX08shobwdGLf4OqOhPdd+/lBNZ8x+7eKUXWoKepZqvxhqj2HVcAve
BGp8ibJe4it4rLAexdtMsciEFEYhtEPScTxTQ4BQho/ePmWyQHPv1BKU9a0JgW25
w5SjsG2vYaZv2rYtsw/1FnQ6skQUMcKkni2IEAYdVnhuFuv56owXkunWf7+lYQSs
LGNt86FpMxqtwAKVLTCHFP0QrDYyPegvxxvUQ47pVRcVdjFA0YcSygB7vnMnVpRx
bDfmkku0nISdgEc1WhCsnEUuz3Hld7oDWdB0SDepiiQs2A4Os7UgJOfNbWzxfTdj
5HW6FlXLCaol4z17OEHvkbGsKdQ0FekrLAiZXnSUbyVf4N79XBScU4mfpNW2i56T
aB92nhyzziPhpBN9vWP7/S+WLbMhMjStdD6uAvm3ho1Cf0MXtTL+WPPoa5I5jz6k
SLh5T+oHYv1ZrzohcAbK4BSCrhQ+HVcBU7y3uNJ3TAxeq2hr16qFfkiHolAUHW6q
u8276dt226Hf/7VFaRRWJwjd8Iujqi0P8Dl7ETKNI6RgRKSAEEpahyBXJQ8RkmZ3
1/Dk0vUY8b/UrA5mMEFnLyyetEByeHUsE01P9Pcia5PjXpHTL3amr1P7clwjuNE5
Lf5WeZT0iIIa8YGG6pVadZbW4sCU1ERma46jsQ+qZyqMSflsoTiI48KFhY9E5e0A
0Q1Oa1pkBvvp0S/dXAx/EwybGoPFhC75HRJIXAUwglpPYiIYmIdmYSu1T52vZ5FS
VN65pWP+foY+Kk/NeQL3028ZSn/XI3ExAhXIfKaS0jKJPhh4sfDQXz/LnztN6GjL
ByiNsMwLQQbHMyJerkh+R38PyeXFggoW2Pp9ilMVy09dxYbK/jGgk8BkIyvTinKh
K5V+L4P+8Od8CFQgr0YpYr+LSharB0YZYG93D3F1aM8UNKUrG9qEhKsi28FBP73s
Qodv6NFYneitTOYlwFXzO+p+fLOOZHHMfTazXkNxeMgykH1Qrc0Oc/nD8QdlQcAZ
EsmGrI0vhmHZVGrsG3L/Xbpks40jkumF6+qJlttdNJITVGOy+Hlxa+KB+H+N4OSf
SUUJg6al6Lff4Z0m6BBysQYuzXPvmji7XONZFV5sHzx6zwDMSOwrqoLR8wLyOs4K
VFS4OlFOqHJr6xdibOmyOTjQ6Axo5R7RafU3QGYtQT8B+SKeWea34YX8BKMp9ExA
ycG41YGGBdc2oKEzpbeEITZYPJDgFrNOE0P4kQ0jeexCikpsCrxZ04BGLA7wRIUm
0TWf9Eo+rRwEtzNA7q/Hj05nUgTAN1HgOtv+L9YcuveGW929p+vGX+zjCl+ai/I2
IYjP+cZfCyFimwPoJ0Kx4xrnOP8qaEYfFbdTmpPM3MDl5rc36zK91GqgiXxiVOfb
omxO9cmZhV5KGHMJyZl35i4RefBEH8xMdQOwqaU9ufwfxFD0hwJfaXL1xRAPQ6Bw
8YEcPpvF/IAK+DpYBy/6kuQRhdIQQWbbtcg6upLRsxBEKo8h0vFMg822IWqNf8LM
DQg0RemIK8Fy5ly56V9aR0kQ0YT7sA1l310gFNJ8Ngkj07szX0vh/iGvqo/qpu/1
qUkbxQTYsYBeRjSOXHgqjXgs9hn22atTqx0GrEAEXLmUN59YSQ4mXH5sOdA16fy/
jKgq5cnYF3AZFyz512+iUxcKnmazMr7mB0/VLFpZwJlX8bldZT6gO8O9MhJJsQHj
sOsUhdAgXI9eJPEt/hiTmSDkCPB4Yx+2mXc9iRKGTKt8eNkFppVXfj/JfpPANcgm
89vS+/LGenV8MOUEaxX7C7bcBhvRFnAY5d6tY3128gFA0sJXof+NjloFODa/bRIA
j1rnj7PdZ3z1sK0gUaRq0owhVjcgqygIR8YJGesC53zv1PHlsj9ecbYMNZnDF8Ty
B4EgdhULNmnPWLHYHBb+w1thfo5P8OVWxOKIinjijAMEZFkGPmF0GLrxBG7PcJMR
iVK7zFsYw8GlFFsXQ2qK3XnHaOMhZYDzqtlQP8XayjhHCnSqrEbDZglf3byVU/oZ
HemImxinQ74w5tRGjxW60X/Cc+6k8UWfnad8g3rg/AfDmcQQ2UjWLBGW9RgxIXhl
rdcqXUX8Hm6wtItYsFfYvIBSt/oUBGWRNszeji9C3pqnasVyDTgRC8Hgj0y83Hk+
yq6mfpL9qMNm6PUU23DpYFXdUH3l7ujgXMicmTAGmf2f9CzVRGIMo5MHn9Ax3QA6
XSuXRT2T73siNV3Qwgmjn9jgz6TxKr/wSarljlbGOIayr2ST7OpDI1nBzo4tNLof
64tt6RjuRbJ2nHpG6DAHM0sB9tSSsyEiwMHgzK0+Cp9Cf4d0P1Hxls5EKxz3jHfx
5inBDoX5r4rW3czBM/7DUe7uZd/zcRVxdbV6Aish1thHXUOHovJhLH5gV3kBrTmJ
jP+1ayUJ7ryS1I5yH+9NzBCdo8f5EebltJPm4+sNnYDlNEHVNYxfG3tbXF0G+bpI
OjM1Q0cNlb2ZAmYMfuyWXOcsVAz0yJq99Phn13D0a2K2cTP38AidpYul9uZRwtBZ
QoNqlrHtiUunOKffc9wq9PhM5KVtoCsj4Y10VRBnvJXZRUAZ2+DqGhtgeWCXK7uL
LgPcXzVuxinPUfXEPbbkI2jDUF+jQk8MXDV0RAVwKbF8sqVmoTaog1a0QAeCPRhJ
DLVx9NLa//ptvyKJozhiup8zJVjxMPgzUgWCSR+SJcn78cqmm3mlApxly+Y73/D8
EAqrwhEvGyVV6l84xPGKipWSYakWMtfS0d88kf7kqifN1RM281U+3Qc7kXJcMCE+
+NaNhRmjgy/z5iieo5XDn1JxyDay7bd7Xp/fFBfWubfS3Av2egZVsVUlYiKmYWcw
t3pUDlJB5UUQJyKn+bFDl1jMEwLEq4bmTccw9Ko8r1GrruEH56FlHb4syKJEgptO
YQJKPZkqEo2M25mBPpjscROa/NPyP2m9mt6lmpjRWFF6i/ykLzOAKiWeEJ5T+V3V
56NRqxB4+JXaT/Rhx1eZp03ct2aumzr+V4i4SxBKo5ooJyBxSEkjmXysOwtRWaQ5
1pTrOfQbx0MZzLMOu3bCledS5vu5q+Ibs3wbeRJGGWQPWcTvYbZARAQyz7CpVlV2
XTT+npXqPvNM41QhBOd0yw7g91huE5C3Ot8IESZcsHPORG6CTTjzzkuetUSOMLTv
2nvvhbNkw2kcUywjxc8uaTlXOxnQJIrjVYPT1RegUZLZNfeytOJrBghwJ65gXu0u
HPN5wMYpGfI9PFKPPJHn8mkqzQp3oZja6tCGzNPmZ+7krUw+i27Dn0dGd7//buGG
1w36BGVztUQ3pLE9ZOaA7Gcc3ZwWT25wyBOgjxyxpNYj/8eDdUzWDYHDI/tmvNZe
HWfJyFwoKyGyP3Ztjio7pdyTX11VEopcT5nNbi3s0sYnfpdZwrpb3yDxyzQna2tZ
Qu/iAcHeoAjNzE0+coXlm+9VzsGZasO5IF6tXhuMPhI+Tgddc/nBRY6/XfddvJoG
dTQYn5apNYxdfEmg8rlFrNywutXGB+B2JryQqyHLAItkq0UDKRVuTVmEtYJCsrkD
DpX6MB038ngZxeYEsnaOATyaoo/2RQLuO2e+xd9k7MWgkZB4Pf2Uo8HT2MhBIKdJ
Myu6aPloUvSpROKRsuH9s+ttR7VfWLYw7+Hy9Wpe3kIT1GKI0vYulUr6I04PiSsh
1c514RyRgoJ6FNBR6A8vaRJWrw4AlXmnsKtaG8YHnO0UjW8Zcq2FHX/+mUa6tp5d
i+OOAjMsSkRFi3c5GscVpE6Viegi4Zl6CUROWdEBaY0DDo24Pp4o/48/BS4PqLn4
+o1MGNkizMSFvn5qUgz2GgECfE/+MseWdzFBY1Skr2eWI9YyI15Ki+z9e3/ru1Ks
Xnxq/fkvvUDBCRVLYmyWeVrm8ELlqNEvELDo8SllGv4WGn0vYGXhbSZp9y/TA/Kw
ZfEfYmtnA1I+L2Yb9j/KR1ZkSxQ6JgoJvlxkblb4eTXLL4cV27VbOlMzelhtfsYu
vn/YK82Uw30aFhgw6V82uilVHlDVBQJsPZiiN6fb/CefkHggacFdGBKcMwnLYuwZ
bzVeOZXShq1/D2A6/TMlFgtLelpE8h6qxyx3+HAOH2RUw4+FpDpWp3/xSwXykxPg
4HL3OrQaw8CPJkc1s9fmEwOMgBg35dKMH3s88s2ylSgSLKbdxJ/RLoMKUqR99tmi
KBHK5ij9pgQIi5zX0I9V7i9vfLSQ1EomQ3H4lKPxO0wm5+UAK7tyKPyhUWsFRcWZ
0EwpRg/36fpoLQ5TKlpY7Nj9s0nkIDbD80V802JzooRendjo/eDjKx3WVnoYhUMD
PQE8B5t+1isJphoGjpbH4ozOMy/GV9Fvn/UJXpPyPhPlGWB7G6UDaUtLSsUuqKIy
cEB+53OQ8Otuc911QUkh416ohLx8dE3dbf4B30x/BPSzv8H4ouz243JQNlEMHKsU
ipfyuZ2fZoN2rUp4QcbqMQm8GgoAcaOp2tHRJW4dC8u9FtS4eWmOfJn5N078JZqW
79AJkIFDMLhbQ5up3nEVP9Mvrk5ykTB3FIWPNI3NdfyPrj66IljxN1GQSjqfZolJ
rGqAvFNfviJ+OD+yxJUtkKmUQn0L6djGInJfxhd/XWtfMW8CwmafFlir8EbKgvDx
deQYjF7D1i98amhVkvbsGOz28Fjf2mvIaMXlM88Gyr/Oyf2HFGM8rptR5Kg4kT6l
ZqoVD84Qigfs53eaRmsf9ERzK1kmkNamU6gI5ZvPrkwkNYEYfGfPAOmV+5En53PW
nU2+yKdk9tXzWQwFWnEf40MrGaOvEDbExH9LiQNEGbBc57gHTkHihR/IGIKvtfIO
FDd2WwORijMkOFQ7K0J67HjCz3AfGTfeT+ATxNbZqzZUieO1fjWJtizOEUyTCPSy
bMTrncobwZyv21VeSi6ROyWk0XKrOuj3MIfB3yc9UVLRPfYTBkM9Kp02MMj0iM6/
+piIsdLFpaYiei0SyK9S75Qva82tRrZnliSBY/mpWyxSEHPej/h853cGY9qWimkR
+pQXhyvi2y+v+fjPKG3UYexcGINaxVYFFiebHl4DGmNWctWiY5Ko2wuYwVwRBMXD
J6XVYxT42VmGtOtln6xOTYqimq3KPI1/B9xY2JabeO+4wzE42lsURwj4J3RMVokJ
Lz8zS87SMlm7TJa7f2LpdFO51/hOH6WA/q0lLfYt5SojxwfnUOLYALO0voglBDtc
iaQje8Mg3zAu7SOuvB7OZKSY/5TChypG0MTNq99ZP3BtdXhuHHOP8xcS3hUBKbZx
ml0AvhGNOvd7nvCMXW7Y36zCLL2L3Hv3wB6gGbM5CInb7WkrvMEJCWuIssxn8vyy
jqxrWn5AjFufyN9nRN2m99T4loZ6Gp9ncYf3Z4RIGQL0zrNXb1RbGNUYDMfvYqJE
yfUisuizM3ZfwHudtY3LE4Kxabi2fsg8xfFtnIBfbWanNY6kZPT9+wb4Xg3OtJYH
yyxV3iKl0UuvpvNOnwn24q8btjXxR0ETIQ5ZnQPi5EYh1fK3e992HxwQmhz6qy8Y
V+GZ6OKosoEg19RZeO+f+j2tNMxSc9zKmnkg+nj02Eae0BdndQ7Ey8uzJH43gX/P
2k+IwIt2B8giOKTFmYRoR5TFhn7NW6GfqXEivBR8bKDNCIBPOBkrZWKWthZlmwHT
AZ0grWPdpcAMBn0ufFU3x6D7DPf0a1jihyWcCbhJ3ln8ff/v70Mr9/bEVr5uaskY
RMtIwe7FXqWsWIiyMqvY/amJQaEqekX07Y6fQWbGw1cae84BfC6hafEXjxDu7Hkx
5DKsj4A4nuJavwOL9SJ6AMJ/fQbVwfUrI1Iy9rkPp76SNz/k2Lp6+9+C7JjaXxLp
j9fFsHH9/X5KvwTH/X/dExW35v7U3iYlwBOzxnjozZmlGE0KuayCTF5rcCy8SccO
/9Xtu4QSmuQ+hAGLgAamW4bqeJHKVbaT/s60hqtzpaXEOP3/O8IzcYpXBTmSi8Gq
TKXmPHfmO7v/ZKpiyCibt+BBt/IuUC1wESVJY0eSui9CV0OmxFruYgb1okdN4wDD
uVy7bK1hN/lsoSMZ+CihsZ5EpYNqjHrJq+68MZIJ6AcJ8/wd8AfmHQw7MR8moE6Y
4CsCeKfIhpsikSolA3T+fht0vn0w4Crt9AObAOnagxFFQpAH4eQwqxVjlGr3cbQR
oYNgqvufb8y8gPiL9fCN0EwaDs2mlYknlNDm22N7M20lUtiFcmIbB0LP2qM/c39s
hyHd0F+YkZfYvVwMsGBeWYOlKERMFgNUY/mYJNm/xurNakpGOyM39yR9cJOWQSRa
rk1fdjYTB0c/cZ9JLvt6fQslzLEMVXsvAu4kXCOvVxPdiDBviBvXTypF10reU2Na
fV7lf9KsGCUbH1HkIRVASOibLxiqjlu+IfuekIaChpE8FKQpO2SdOuoexuht50kI
beJ9BiPUDiPftCtHdswNbwoPHy9ITcn0I620UgzuRYJLfjWA+NHH4oczgaMtDMtz
oXFSuQuzpsqmay8tOFCttfyJI5Q5W2EHuBrtW3UzFyibabfL95gTtuenCwSL7BpA
jHXds04drB9nX2dz8expsCrt7ufrUtLtcJqWW2CVVnjnZ2CUHn+Plsp/dF6TRB+z
WdLnehSbDlY1kXN4m5s0jZLePQdTZGKsF6CAF2BF8J30Jc8AqOtdc9kxiLW6Q57w
u4UQVohVnNDsOG2B/1cA+dE+U4MnMSIyexyw+9rqb63xEb6wMeIm3FFFm/08760H
TtmwBXXOYtKZKWT6h+aYFUQ26fgRik4pkYf827ZrxT7uaHpFWbZqN6pLGr9dZeVl
ybuOYL1au/5xlfrixB6fjWae3Oow2hQQEvY/E7onn7zvArlxSr8nMg2yATQHy1nT
eNZ3oiklNbDH4OXfSeGgcnGxKL+lUtZM9M/7GnEhJj8Piafy1KHURy3eKsQUmSln
VFqfbJV9MeAwcwFTahbqbP2Ekq3UTDt4pBD9aQ0ZsbMMtfQPrpVrbLB6BCSMu47M
9Pn3fyyyewzWJPon7/RBY0Ko1Sh360k2DxkIwc+2cvoqq1fwesA1TRlj4zrJN9X3
2XJm5cP7J+hZadojtgmMvXqmQ5faBHlDWaMHn0ndIS/LrfznCxIjo+1MfLsmuxuj
iCPE1qfNr2gdUAQkdV6YpRRmLxznu/57DpguVIrpp+RR24s//ZcZ/j+zMmeQDZHO
iuL7k5ysAOqIsb2gjzDBQop8WczMLWOtVfpREs52bLVpQnD/9MdDhvb6qJ5qWeMr
eACdD0H6QcoANo7zod+3+W07Qv9WT6mBffxFG38FRhwlVjU7UTapVbcBCTGnEBi0
n56cpe2T+hiDqHALOxXeilZrcPkitEiXdG9Anx5tlNnu5p5soymOnGhkn+Qf0L9I
t3DybCNBzyjm2EzcEWhY0BthAgf6jMvzCAJoj67ZFI70BOEvDiHx10XZD7qBo3yQ
COWB1LAQSdae9H2J9uw4xLiopWcMeyBiOXgp+k3d/JY41NW0cNdUvQeAWe6aVYGU
0463QoMlPberjlY45UCyJGZ23sbHdmmtR6F3LY/1L2ZSZHDQZSykIw+yYzAlNm4B
GuoyO4J1FxZMnzhxQQQSh6Wd+ZIycWqC/Lu9mTzL6SkL3vBeRMzipeuqiiCOZJrn
YqrR78DG8UfVPEMBwSpQpQlpz2nM1UmPbJ0DzumAHST8cSwvlmRUCYONqge2ZmDm
SepM6pACFT1/A8H1B+kpJMA0IDsJqG6NvPE/b2h+Vm5ZTNFiGR/NTDrJQwHYCnxI
7Z/YAW10XGVQrg4w9snW1antOrs4q+yDW+HN/n0esPzq9zgWHcIo5WlPaZeyfyJc
xYJ1YlwzJykiFtng2G0BYnuD30y/h2QpB0n2UfAJXrXbwpDljCX3JmhGpX/Nl7vp
L/SfdJ+c4abM/swiC+mtYuhYtE2ORGpZMG8zG1W30YPFdkIE+GpbFj4ixI2dtlKR
yUam0EX39DGMSeNpmzlCIbkp5b1SMSK0BEpkY6H/DaE+p5Cl8hKitluJkI37RJmo
dpaa7no5ebseBXEshOAWeVuId2u5wb/AeijOvDFR4RECmAUlorxeDu6OKciA1Wu8
Ype7VNKmKkUe82hP/ZL0dUqP/tlXN32VLUJomGLXorWMGSge9WI7ZcoLu64s/P2y
V7HY7NF5Cxkuf/4+vBC5etDkwKfV//6pvVOjY5sWTziW7Yo88r5sAQsVjjPtziCu
CKG4nz7w8D5POEb3tFHqLWnZp0cnikfTJoD0ex3maCM15BqVvxrHNGtsYuNkJ8dZ
UT08P7MUdXvSqdVx4wkhM8dGN734RuH8VTypF2vkB6LIpAqqWob7b3lYYz1zAOPw
XI0ve6jXWzSlBUmv67jkqeaqwqhkka1BGIHMwoxsCfasRbfeiY9aSpa2xU3SKgWy
bjBpasoDwutRMkPFHkKI5tyEKRaC05FlZzn/SzlGAuOEvPQ3YlkZaxMilsPS3664
9SPbb5NZ5f9/Q1CdSSfaYap8gVoTL3IdTsSp55kTBJDGg70ZK7D2dpBn115BPbFJ
3jXA41XlHkt99WP2BeUaNV6hzI7REfVVZp/VNPSnoY6NLtjYyrSrVhtnEHxJxgRU
zcTowb3dFl2Z7enwaMuBBcob8D4Bq9XxnuH2Eh/xTkubyoBESqL0Wbuxit5chaKv
Qh0GowUSrSjA/ASKi4kQARqmhXh5PDzU6FU3ZMNa8Y3yI+cgJ5dnm5/9+GCTycFn
UtYN8Nmb9SaUuPeOp6PDeNbZHQTea5XRKZef86/L23+WkVgUE7BfAoG8JYGQ0pwf
7hhJr4ocF+NJ9ZCQXYD+wUNI/LKAlS9mSJXW7gwtiW4aA+0XXzSsiHlB9ULSyJNH
K1iARytlCdN3SlxpJcOK5Q7QSy3DJDsQfWD4UNjbsa4Fhw3kJ86ipPRs1LWyHI1n
SqWldaDclh4ihiSjMc6yPOE9IQMwXQE34mvwR6TYiu7EJ3pfUvFyl6x6KBSOlm36
GWfhmGWzjz4uClWnPUG8VwQexpBZ33HSlCRTUhIHVMP4hrsvzK8u7EAgjyiL/+AO
x63586sfQuUyNlkVZSocXlBBOxzQLNFacNOwxuq8Z+k0LAiT09gYA9SUE/Zejsxo
pLHjzWVjQWn/Osy17KU0qxPwD9jq2wIKzqRgQQrG8H6tOfui1VXT1EmvIb2hFPW5
gOaSAPt6bGcZPBhDlGgFtlv7vpdfisBc15VHsm3/ngpPMUlLoFyYl38AJaKquCJD
ZsTVCU64zsEbuvtroW8ohN4NaGgAy6f2TtKlmzY0MvvMenJPmpqvjwS9pSgVmukF
MnityHFvz3xe7JtCX/UDRVIpGHk6zc+tlq98IgE5WRbRosMuGyxavta9XdoYT1SS
ChFiU8hohRtWx0rvxH0x/MmtlCrG3+0ii65mT2ui798fku+og/46DhAjmsCXhy4s
d+7Ee8GQmqEUkvFSMv5dbwS7jwo1+1QzKO88C5izY7/m5ptfkTjRvWEqLYQ0oHTI
wFf5vJbt7bztmLug95hMipTEMlubaaUc6kLwKReuol10psa4c47G0SfVZ9sSG2Gk
32P7eEWsMG2xhha/6hUMjptsOBPqpc1Z3JP0ZfPYUQO7u2YI9z39YZL89+6gWLft
I9pJYkVhH7sHdmiuXabFsnZVlydeYn1kyOmWEkApO1EBMmSiuaVHTksydwD8lOsH
eWGpXWZCtn67YAHSK/rEFtkxh3namHVtX8cklTkjCBy+NAE39JULInovt5rLER+M
WG+fPSEOrevK8Z0l9NUJxE6Qy/9Cmaft0z9uyZ+0WOQ6O4re+QGlTgOpVDQEftcM
mAYuyb2R71JamE1AIE+RaeqG/A/OreaBu9tCY7TlEYbvdlaWC8nf/FHq/KfpY0mZ
r0HBt6DLb6UW9as+KIbZYYxuKuPntquiBGujrFwach3Mn6NbgfFohBtPJdFOkAUX
SKC7jR9SSwQWm8eRC/ozFHWUVXe7uip0lnb1MqNLnLEWmQjPkAQQzmVBYNCrSkQo
TQ3xvZdMSyhdt0ln5bPjm3Ju+5CSinmKqxfWcJ1urXz2y3QtTBEIgt5tvEjq7+2n
Zmhp5txcDyVLWNS9hznDmtVwWQpCHj8kQ+TEb24+SrEsmJW3vcprBQwPRtslj6E4
FEFPDW+y+bg/tot5p3XZjsinx/PeLy1dh1bBPrFXzcc4dpR+7V9qJrT5TaOa//qH
ETXoVS3neWu5ev3HXHcao2G4mtZ0VAZt03hjDqsrR54OeUFy4CvRMQlSG8PHs4FU
Va7k3Zt2GRg3Ge7GO0T8/U+6VYWCxvXpCtWQDiUiOoiT8FHDaOsEC5kjsT0CZ1VR
PgM3m8z8msveJM+zD7Bfh1aGCXJjoI/pvX4BKz1q/twoE1gO3LBik9h+mOc9oiAS
hHL4aD+YJe8/RXXpRa6al6FwClACUSIlIp456Fq1cMwIt2IQ/gDnEkK0D6VKg/ss
zxmNYtd3qzMj7owoxAnR8ebDYlA5WdRnRxBryv0bC1IF+7kY4XpC2ta2gAmuyOSv
4WUe7KAwMDzUneAPL+2c9dDV5BU7U09m+MkJ5cPJ4ZPCegl32cxMqjEk8EuBXjZz
e3AWlBkp4jQhbLNe4ThGXx3KRS3ePnYamTNb93KaXO7Sv/f3dQztExJZEL0HXpcB
CYcI1hZa9kYK6wc1Ha7T/iMADpz20jRRKtgotxOcj9O6WcARW2CJiSstmdhWGQkG
1bSuLJBV6ILacixRgcuPP6S3C4hx613FWQY3E4sA9+GVwtIKuLPxlgTzFz2a3qDk
dwu7AUBXQp+1ixTrNIpL7TMg68qAqtchygfKin4z7nm2vXC6eBidHFSGpwoU7qiv
ZDqaa84QP7fIEm2iGgfYY86/euyuniOy3qtHNhPNdaGOclDItpvAW/J+R5HyH0lC
gW5tSdm4Cp22K9WlUjPtnEfAc5smFxy7Z/pmUTpgcZH2yE4bKmub7V6gOTs0HfKj
GxQtHniJc4e1cL6GcbXW1L2z7Bws/23Zz89KlQAyuYR1eHKnHXCWAzQvYmB/45KX
5oTMvjfK71jaSLVCqbecpzVommYmpEX4XwjZKEYS8Q8wEHnPNUoDpekoOta9EJjt
eB2CGLzcmzH3PY0Mu2zGvDM7hc8IEvj3ZW/uDVqvBfLD3HMwnRmgAi5vXNMwc9yl
anG81YJ6ePj5U5qS5b2zTFGkh1kNEZKN9bEH8bxzeNoYIdNfAdP7+WZPBOa6ic1W
cyFui1Kf7EHJKAK1IRyFPem/YtP/QDghc0eEUXUWnwEB1aDMqei2osVq9o79WSVL
N+y+kVulIsSf+KEEuB0IFGelZ06RyNnX/0MfasXpGREQzcRJ4EMCcAodF3AnwqxO
WAbH3EhwzB5296o2sG2BqAUQIu5On3tyrH6rA/EnCCafJCragfDEwwCmYCU3Lxfm
QuW7ValW80w4pFjN2GyrXry1iqlmNC2vpaTiJH7KHURmnAyxuZ64hf5FC8TQhAvG
ekhpGJMy+6QP7owH7bDj7zmlu12vCvCUZ+BZdGDWLpBugCyK68bEhduY1K5HKZan
gLQbMFkK0NRXFjTgNHU87k2M6p44ZEnWJcjhNKiBROnVNHD4HsqPXph33lRfuszS
uWZ24hqv53qwPdhwcTT8ejHKLadMDvesyKU4Ud3devtwv84aEDeDUSzQZUTFbK/L
QKgbET8DTG9jBAkrfZ9bzgy07St2Lb0H6cvzj0cybnoVb0ZxinUzT0UUseTAqllN
17UwO3bcika4uZAk0kAucdz5xSvNToDEimxjCqYhqjf9deWHuCQcsnipVK38IeZS
sfYJwr54EQgK0RZMom9DRIBGLwPeHnteWc+uDLLoTCngWRUfhFYBbSqqgcx0wYgm
2sMJCjbl+hy3AXlppyElRamI0POTrO8id+qZaaiwn/MLxsBayqcZQLLlXUTYxTb9
JlFHl67G68q2O4sniKBpzI25EJGgnJS+5vbsTn2x+b6U8Je7EtCYSHZyUcWZ4BqW
dqy4PQdc1naJ7MQ2aBgy+MzcpVf+ZAjP4bD/AE3p4SCbn9byoMzaDTNNGVb7ZlNx
in5qhQcAI48/EAxmHobsNZgpKB9MhYCauHIiIftpAuSAIgozo3ZzScL2QvgEkGXL
+fi3sm6r6e4ZtJ00IQ+MhlrUbqC006OeXa7BZIjQH6Z3TCOmih6qt4ru4eCb6hOG
KOA9WLD4BOSDYj1cKha4aw7mI/WFR2zttQSpOMJXMYtyqowBv3oo7r1o7Xd0owka
lbR+KFubExmUU39GEhE83XdcAr5SJrVN6dzUlMAzLZ8SxgzUcjMl5YJ7Wjr8wgmr
Do1siKvjWu4jSFcxnfHxnHRXGP7tOpey7lPeWU5mBn/rGnOm1FWUYp4y+jFQH+3g
EYvfIPHddwcf/Fp2rTRc/b2oGwKhC4PTVYOcZBWNPaBbgRXfWg87SXAkpmnfRnn9
EhVQ/o/BzZfcvCkaUOq2bCjIwZDrz06IyA9Zo3l33zb2sZjgvQELewAe3w4d2Df8
HbGjQ7h4vOEbyzPhJiD7GTgIbKqtMEiYo1c/Qwqn6Rv+b7tgudbCiZubv5xhmtle
YvAAfmVANe8H+XwVBpjtsC4ahffCPpVgoqurdc6kfFFZVEOJZ1eBwOadaMoAqBQf
VtXV6+w6uo1LOa+FHz/uLhdlX8VbpL6+DtIxoD8V/mwHQn/cq4j7S0M19sHTCHK/
dzFIL+ip57TkqtinBHvHPlyzd3NB02Ed6vV9MgysLZyWxg9n8A1b2rehpmMKpCh+
ctdloI4OugDD9DwSfn050aSQgkrxrYpkd5wdoylDyPWYOdOS66D5emwuupdGnJr7
vRVsnf/9go7t1ELXfnkMEYWVXHs8/gfpAXxLC1NFPtpU2ZC3f8MBFbuRfavht4az
hSNKFGC+0C9ZlTHAm/SAud5RxBw8OpZ1ZIaObXAt6S51TNbhhpjFf3Oqs1ryQB4v
RtitaMT+w0z57xAZsApXKh2TnoZULW70mo9/kKrHuUx6orAe8BdSl1IowPlD+qiy
FvoFmxOkonkz1+y3ySRIPvC8fH9G8WmJDm9a33yxe6Vqb+BNsDLCYHHvgZJzhePX
MyiL+7QQ5AO4ftsoJWtT6NBQ9Vo0R19Wo+zLwVv0sU6eYrfA8Jsx9WZAKX8J8KOg
Kc/z2bv3PdXjK8Wxc91RkmL4BPBSDqzDjP1QXIGZU9By47JuF9dCXs4cr5wdpt9S
IPGJH4y4Go9k2Hjcc5kOB/mqQrafVRGXvTFj0y1uupcBY2jE+48mAu58JSI7Q8pX
Rvf5ot1m0gaZmEAluCDkd8xmqJA/oPwvo2cTBIkkxNCNwNk0xnymbi9vc9Lgvvs9
5hQPHMzlz+lh3Gbpz8fTsCZzY6dFxXDqCj6FG1McIv5Fjy6qcN/cfPApv7zYqvIx
CbTuA9jB2jZMwbQWAW3Ocm8gOetJ0xh7Lp2dpdR9CpM8KUb+Ze65bxbReGrwKUT3
qeleZUsOa/jvPsyALrhqWEyBhaxhcNl9rc+VurPSBkYppvh6mNt3XuZH22EoV6Qf
+W2Tv+tUsN4IX4A8633TwCt9cqUu4AF7C1Ut1q4YhPhj+40J+9Y40hvZCSwK4Tmj
SWM2wZkJDF88dtSfPN+E/dVVTGqBMdog0IZLz4rlqFEP+h3ZtDHTR0OJvZVoZfVl
c7CDzRSKAtrdzmEfluc1hdruaePhyu4J3eTk4UQ41C30bhRG65FvKMybkmYG93fi
ib8fO2GvkciplzR+4kMS0VuoPAMKN4QpDBCwm6aJSHDNp3VofHqDzDHfWaZzBSDS
6YBBX6fKijetgFS94EwIS0DmRmrNTRLBvtnLjzWbru7ea3SmEjYwWrVP9ZQTud6M
Yc50yJShL8ySQZfp7W8HIkG2sQdaQ6/rkY7fbLHmGuKcC6T//OpTFkmeYukD93UV
gYq0di/YqHfIr5stfWS9aLoffaTlIWVQb4LppfQA0FMYFdpy3YooWmVYt0ry2bjB
mKmblwgjVOHhqgju9hMtCepzf3fwRi2ATp2+tLv6GuswEDXDIMhF8946OmG3rmuT
v93n9HzOkql4+Geek/Z6STTWwCKoSToRJ7/LoXUD8Yh/qW40RyFs3BOIwGVHLWw9
30+OyPUHxjPB/hMJ0SkuYEpjz07Sx6z+WKdYGrsSA41BkD7CSir6/lrpfP9tmYT5
2pWdzuCfoKHAGNv0jINU+0vuPTMhprzFup5sG7Fo9Xecf0zUnGKnIfzyx8EwCJUv
97Z4/CIbV+Z27BhVfUlZCAkkd4Q2EaLO9SmGp1Rk8rCI3Sk09Ikx8w6Zz6d1opd9
GKytXXi+M0Fa4Lk1mbwKYcOP2Z/cFw4+Vhv+e7U1CA6nApHj9MiRlMPjB9L6Mi8b
4IgKAV4ho1hXz04fFfzjVj1qwfir3UwbSyNt5Tt6mOjP08FtdIt3s9nSn70UnIEO
sK/uZw0M6sMecHvnaKOLWmG2uI9pBb77SsGKTBe76YGxLRW4RHf2aGBiHJyl6TLZ
LesAIvMu79sSvyQnKQSlo/M9gHn0z30yxoV+pWaM4MEbtwzVy28U4FlyL3ksRYFk
0PfiU87kdYI/GfDfbo8Zskl2UfhnECYNMKSsIROe0N29LbpMgCtQFxlzNY0wjLbU
jcNYLEXHyKp/B2kHniqw58+VKFSjtHUT0wLfZgDmNK5A4qUWJVDIy8Jvv1J51iWx
DGNzsTGUMqUWDrtJEzlc4ZtE0tEUBfm0vLwETBJyaaxmdb/cgqEepwC/sfDss8da
R8cyOuqD2DB2LrwwPHfyyVDLl2GOTO+rxMlGXY+aZD2Zz0ZcBBdN1ctXWt7hUkUS
s20pJrt0LhsdyXlio9YjGr1NGQzMhMQ1LyTjO9K71uxEZ1d1fgaYqOMD4XXJACXj
oSYD6Juw3NmpygznU7K/VrjEUHZTROj1dTSvJH3MZHeEEZD3MX8sABOhpF+Hj4Bn
vqvWzb+hH/Q9Sea8IHxokCLklx/fXWt6240jepnaKg6PXb6jjTv1GQ3B17v/7Rhm
gRUv63GTimal0c6D7jUzYROoHbxiU04Cypz0qQWMAixZ7/2U8JcCZbCIykutj7OK
fMtUr1RmfnseWeOmnOldtKazzb0fqX4zXlN80n+pobsAmvtkG2JJlCy8e76owWfc
XukD8aDrhfXQoO1fea4CPuqzkRF+VEYE1M9OjvWkXli0Bp0n4/nlK9x7Xex5L4HK
AnZQlM0fT4n+lFt37vXBMasiRiDRdvI6vKNlT8TdQwPHEp9tLSzSGH8HdG7ULzHC
0p4jScsRVvVBkydEjTFAh0qAC+mNZ3Cli4IdGdntBw+DPZILst0gZ87kaYAsU6kn
nY1GULwBB82ja1gOkdnpl/pc4DdzEoD91/KaA4eKRbQQWUP89CqJjqXXCEdMeHL3
Dg2jQTaLryLxpOaI5lzx3QPAY0QfXkpwsa6LN50hmmIYj5cjveezdx4Klt6JRpcz
2IoE3j2KLDGXDz+qHR4N//dYM//JAWejMjjp+WWCZm+kbNFvh8gLT2+wFnq+Yga3
wcttmqGQDdALevC63dJVLgTNvzdk1UcTnYuzZ8g6/RRrCw9LzxWU8Vu5gS35qZ3n
wzjkxJ9aE7p6swcmkQ/TOALQ8nnghSomkS50ecJ1pHniJi3Lihq3UME/IvpInWws
MCT3YMXfAu2JA11DudK06b2iZVuY2W+HQJZNAlQWptkjK2bHVA/ENwdgx9OKkrDR
IOCL/xWJY54qdXM/1CN+EQ5vxL0JSfVmHZEikHgftIZAvzCAae7oTtxpMZdClgjy
fKkWMc11jPOUydFVDlRcNE5DAHmN0OicgpqgtKhF0bVpF8CzeEvqs31vwCSbbBbS
JnBvZqge6RU/AtyTOObzyNvv23J/vTh+OWIQV1j5prgQXvNO1eF6n0cQmNe/++bE
/EZCbD4c08zwScfYW2lb+RQpUQNt3Skhnt4FSzTXLjfN5PRbTKjo2155g6f9D4Lv
EUWwnEi1GXAA9jozF9a0qauzg7EOl9TC5RnIYeMXQCDZz3x78OunPY7sZupTsc08
FkyiVZjlycxEZBMQJiYcsmZ7N6sZ/yD0y8rFBxLrIZu1tXJ76sEVI6VeqaU2cfIg
R1ilw0MU5Fc309lXg3VgAc6HGRu9d4p5s3KFKkTyZgiz44u2lZdYOG6EfzmytqH9
3ooEQ6gYxTPfJhyCwwDBCHFOFp7YN2VNObP6BkMpHGGRmUUUhspnNNzOQHGEnr20
qsCqqyskqi3OpK2hwhn7uzdo8p+EdyXlQlArOUU1d45ZfsfMgB4b76AhbTgcBseu
6mcWX4OMa451ADIDNlxJqGSz7M6T+CnbAaVUWFiKe4E/A10GtpY6B+pbdp+LcoXJ
UvRB21Lbnr7YHO7/+J+s8dlJ3OItEXMb6U9PhXzxwSB0zllfb0V5czNMZV+nFlnS
W147UN/o52wmc3Tm23+9LJTFXn5PCxakIKSPrVqSK/wcE1dsULGQ6O+0xF1WrGy1
5/RyJ/NaskNiueDZHx9jUI7I79Q+hz/IqHuttR/GElGqe/g9aGUR0hEFdtf4DnOX
wuvvf3zcbnVqRcXhKFDviMcqDyUJjbxI44wGdK+Bn3t+SPQMXYHQ1Zku6CDj5Lc1
rYueI8T1RZ3vEVBvZkW9QSxHL2S+HMWk5NoS9dX2brInfL3MFBa7r4n5fAqPf1Jz
L24FtViVxJWYf6JzlDDPxfh9LbO8n2d0+ohJBC/WuW1pvqTLkvQ9uXJJCMKNTTwB
dnpMeONvEZH3fGDL1Lo18qWeoP9CXwk2ZQfZZ7gT5HnuEXUMeFU3YTdlvUxAOCTk
PJVRrV8kxKqWIiLOv+0PqYsTNGo9drMvgt6/vqJ9w4klojyxiwkdNGWvg3uL5guK
PxSWcndexrqomSKUKbvouzkYMGJZxZ4GUYXHJawavImf4Um+ZoIgcP6XLBmCVclb
eV9C30v1JJ6zfdovEGnB/3FXayNx09QcPIsMwm3IoHOrpBx8RPTjmVtV2RBJHqWF
fJaxxwKUSyw8dCEcVilMveBvmjlyKbv9gMffU/G7gXxxedYZ5SjNmNI3u5jAOWvA
6HleFk9cWgVRaPLc7DtDpcX+H0/FkduphzjEcSlAefc88o5QVydSWD9+JsG+RYyT
2RFqJHmu49u/uaERC9qu0vArNoIxM2mR8uFMuRJPzk326hATDycrp+KKKkM03GeQ
radCCXOmOt1/A+g9fM3HvtMq+cbBZ8/gG42yIIym5sehGlzxQWz0FDVLZEoWhQtG
y8/HzOPWV5xeoQGjWM/4a5SgDpFQEvlbDnwDjNYYR2rqs5adtY8kcEW3Xk/F+oij
/uWNqbftOYOoXYZzU4iiDZcfo6kkMLJnSSVF1dZVZCKcV10J+LbvxmU22pUW9Xu3
9FDOU0z7D0nslTBredSiHzi6d1Xo/HPGOT9HI+4Ihn32s9mYZKkt0/9s72jhWevy
5ly86Oavl3lTzLTAUX2G7/Wx2w+ujAFNxb8ywEX0qKdLaQWcwfN9Y+NvjjjgQjb5
HEagMtmV09n1fCyaKkWdrrNZUX0TTcJteSlb/9wmHhVXkVU5q/e2elm3jpaPGGXJ
mg0Tgc20YDJn2VRKD9O1hDHbbc/Of62ebsq8qyWrDyG7iE0UIxMLre65VlRJhTLU
i/vqkiSk5NUZXNpobftGbbrapuYycuip/J8mRm/5mjBuwEqOsHkm2k2xjYnc59Tq
fHwXAf8icv/xFlGntC+vW0FMR2U/mDmVj9J6VufQcXht13EeNHs5LP1Fv+PGAVBM
uxY3nNPMYbQeanU8do+MDMQRGYZqQntYH9sZkAM791YN6Bzf2nen4csdX87FSo2T
X3v/peqQOEseiw+nQcmZRaVOmSVzSJQjPUrf6jJ0J0md8+gvRWF8W0ugQUga5Oxn
znYQJesYnYlYb+tVQZbD3CloJzBd9u4TFedEseNrsoTrbTJV/z2DP6cvKgGei0qm
44LeRm2pX6yPn8aq+AXU8e54HfrI+RQthtQC3bmFb2Oj/4/XxbpCL5BOSePwLMIE
NR/BYxtVIi9i5tIJfqRd+DnTc2ES8DRrZltHvIJ8BpK2fCN7Q/JP41tB7VOssD3T
tEuMOjay06wsGyaJNZSDeRgFAtQvawJy+BQNtvWQDqWceHynzAFydKuEc6Fcn9gQ
02ALmD4NiCZDQRW3/Alup2Id3qeat6uDhvIYIwL4yTwKSdQVCqwikdMldzqptPMi
xRNXJoO0fVwJ57VTw7s/eD/fv1S/KT5ktp6tQM6TR+lbhddX2ejBGgtPsZNe1ekn
Tz0Qmsk8r9iErvfNgCcBRPUdx1LVP1e0gNMXsfdISBN2Dg07q64un8Nw3PcFDmhS
pzSqcXwKmMMLRQHgqMXhPN37Qw0oOoyyctUZelQmT7dfOejkedysegx27Apflod7
/+Otkaqae1BylBeZcDF1HDIMV94i88ujkQ+ISpu86MjOEZF6ru3oATXL2SLJxO7H
gz7fmHQmHruV5MKKLc74yxRJSTblKJGcPmKxmGgx0zTycFYo87Yh7+Pbf6WzzS84
mV6kcxxWIStukXeEKHSvF8b+kjHv/RVrD4T1riJk7X7fr/Mo1iC8BQ45CkNX5rJ/
8M1rxHX4zl+8sLvWldoyBpyJptPHaUUGkLa2+j3KBeR4mxiobTHLVcikp/CLHckl
6qgC1bQhGLDtjaOs8jIFXgDbrI8w5mgNrTraD+3UErMxDuTDzpBJGmqJCVRgjSME
fyfR7LFLsdqApCHOxJSd77i68O9eQBjh1cVXRHSZrgq82t/nedksJbGo5b1swgON
oxSGR5U/I8prXGsFsjzE55GV0K0r26wdpX5JjveVJN22AXHw+mIQ8EvD5Z979mBr
uhOou7JvCnv6RTC+Ts/uHdYcPKTqX8nq7jxVuU2Ie/n98hb/JHbppbEGWEwj4Vd8
CwHdJfoXG8RP/yhRczQduwjRzEnsyOOPNfohayZyLJsYDL2Qvq+gJS0D2O8MqMSW
6UTc5N/zya9uyojnbF5EjJm8PxSVdbtxp3cmu/oXn3900JMSu+x1jXhJA1CxEQVU
Qq29st/Khgo/Xya8dIAc1XbTIYO0S07+sBh+Wiu5Pa1nk1gZxBipnhmfMgCY8SvX
ZSLfQYiygN6zypcnz4op0zfpbHpMUF/M9ffyyplLmhDqepqBRymkBC4vX/MmcGlo
3GIXzAxunFNC6XuBMps7dU1wZQmEJ379nVJePHIcYPrDcSAZ9bQWutsXX2DdFOxZ
+PSCIDv2qLEhVPCt1c/oKlDZFKvFexAmaFF2ny+T9niK5webZvoo733wrKnBXq7i
/foxV+vaH5u+MZPvKMK9Y3R7Z96txvAx1nR3xW3UdZxcFVxVmsXp3JasDgl0QuLX
R4AN1JF8JQ7RGKB9MDqexO2iG+nkypJgGTZKaU4BX6/jzen5sQZP6JbPwj3dE+iU
sWd1IeTlNqW/zlAfC82bMI8k/0kOGszgTwNpvIR/x8hgsQ70xBYPcox1Nz0zsYE4
C3Z2TzhWA/tJdgC/bcaS87XGPyDZX2Pe736jv1fbbxr30x46ZFhATzyiKWH8wl1C
AC/VUG5MaMKRoD5LULTdT8Qcb1Fl2LfaDZT+oreOPn8g4y33vIZuDdJxeMz0jXKO
ZhLXLdp0M84Bqi8jOGOO8UsOz2xom8Y9xd7CHT7LhgHV+DpAUJ5phWM1r8kQskf9
7XNMAUi27gDKdbfq5qhWIub7yCGikrzpai/wFw0hJqAMTf5xAFxTUqteuS22EhYN
8MohpjbOfNhuE/CCjhRqcHVUwtM1vK91y37dPfpytxE99oHYaCQVG1cEPAt1zoRc
E3L4QgRICIA16jBYtWzdvBVZzKNFGmDdra8ZycIeB+WndEI59tkxq4EUjEryAUX3
vwTsZ+1ykPxTIinQ2kEn2oFnnbtv/Xd4VIpZLo62fty4USznF487SGQ5OQXsE4ma
WltykyWEP882MykNmg0ehrDc5CTiI8OuxPtltq78Bgmw8pZdEJ+ShoVBs23Kk180
FmeAzAPZyFVygfZuksHWz3LZoPrQs0ACgYc7N3TCk2wj/pNp3a4lAT4gumgi0Axa
JakjJLgRSkij55B6sPHMai8Lo+JzY45L9C58avUFyVxwmp/wCBbKbrPMAlN0uouu
ekGpbuZVo+q+QURrkKNtwdRfSkEsdY8yy0dsnnxAr64jb5VPBfTbC3f2B/CHlyxM
T9r8v7cuxtqGmX5aCAtXPRjBxq7x76Cdne+YkRPyuNpBBiI4I+W3dnyTvC1j16JL
TNJEAQPzDQx9nWcX45EvYB23gt3ZeokC8jxOnnpaejrIpgYgvYYpUuBeKA5q5gHP
TaizrFwKgRAMm54SzMiWaJG9AvkP4X1GZhNT4L9zceWJ7+TwrwDgGx5DBtHn/6rW
knDSHeyc2o8Qtu3O+m2meTccIvtv5p9BATY3ELwXs4DCrXddMoc/auocL8la1K8m
Edcbkjj0OgILkaCi3VTv+1GcrpVS/yKiwDdLhqB+lf+D82GV3FJqPsQ+RN7kQDzE
YEo+m5vuphuW/DQ5xFfxpiTezsRrZdHph+6Xeaaasz5K6dytV9+GXjk2FHfwwmwg
OJdEHfAjNuATUZUhlgYnU4M5nLawgc7AB/D52u4N+MbtJuYXbMXyCVOfmY/Nijr1
Uyo51pguCEVAahh5CLr5rRHy4Zwysp+2asUel1i4qDjRtPeA4cBtu1pc+JzPaTtz
7KgDfJKWy+GRk2FYFl2/O25cdd1GtngyECDkhG3PGRuZHEVk3ux9Y4AOp59r+igC
7NjmRqbdYFeS4MQdEhVen7CZ+9IYrNieuCkwGSJFJWZHhkfAq22pLtdElDg9Oq/y
xs5ezrFoF4SEIAzObQuaBbuqxRudC+5gPBJ2tlYisxKmTEMWpr4EjQBkFp92medo
3hEnHZ22qtzNJolJtNmh0Hz4YpzUyvUnj2b+WvybGoHoJPSqMF/jvuhTcDnmbDBd
bPVSps51iFzEvkjQkvXGV0AAQrr1NGsexzpjmfCPDYJ5OoR04GZuSIbiHJSZS1LR
lblMZs1XEx2GwJI8ekuj21aVnOGDzmPkN7rzCAQ58TluPUGPpmJHHtqM2TmQbh97
o8oCINDEBwZ8RJml3BqgINRXENLrI6qKoxsG1xRZyVWh2KceJy0Ve4YDbzjcB87c
QEpvk/DvrMHs66R6RRBO1M+DjAvMjfG392PDdAVYj3A=
`pragma protect end_protected
