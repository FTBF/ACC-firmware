// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:40 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sN8493sYD/Zt6P8V6lCmniCfQlj2KFb8IPhnCVgziVhGrxoJ7y/Z+YZ20vIquspL
Bguinm+SH7bst3qdEWyQALqGDWwHQtt9OkSDN5RrOlWnbGqqeLw6k+mMFs0VT+Pb
BUj1bHJnyZL1ZhHkSPs+pgnMAoUqH5Yx5mcq4K+RYaw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7216)
tysU38B+C1jAc98E4VQ4R5TVuWTfNiKZdQe/ez6cVfXcosq+1agPDON0cymTATzB
0JxMgFp+JzOy057AoEvxwAC2QBuBX/lcElpxcB0xZpW/ShVS4HjdJGDW4jMoHiCG
uQi47bDdwkKnoOK0P41EfbVhVcyDoptwDUMkHNR2Ymsas2PKRNFBGrxeT00PYT+O
GhHQ6xTXeekKfpblefBx0Go0zcy3iz0PIJxLTWQF/vQOtstvTolaQhJnf5X3lhNh
4hlawMoM+tISEZWOfkDSQUxxHRKt0rK+Dr2v4s/kInIPdT2ERD1EKkZCSKDbY0Nd
WUD+Vf4kpFOj4NDNE0Ni9n9lC0xKZ9bzsjSTKdwZfjbFdtnD+IdYp+c1y3gNStSs
LUauLzTqPoyW5XmcVq40BZ6RDyzkM2p+ZDkmZgLvkv2Tp2GaFdeAA9qbSQSDzx4J
7BJFm+R7xR/7sHTEWTzHXKg/kz4sScgGeQeRWm2PDqGqbscXPwuhI3I8kzwRKkgP
GyjTPQFZ30eyAdxAZZkmOrT4TtxbA5uMxfD1AXV+BkXBi7ChqvYSNYSj4nuf5btS
usw01XjyvJbrwD8JufQoSMGTbDmfX5UoscbOTA+fNlpwqeLkJBnJTAe2hrbRmKtm
cIIp6la8BO75ZuasWNMATbDKLhCQ8tzuJvHmwfHtN/tzgzkUTpylmxO9TnWiEyFg
D7Nzt50ReV4QtKsKynwTW3kXFtMbTWFJ5s6RAyhh5Qsqxo2oiNaN0Z+dg6ontohU
VL4XY8F12NFq3Ko6VTEKgZa0PvxpHmTw9CZpQXaNGbz7a2SRXb0dtE3mb5fEaIXh
G0ZBmdZZJ3k9/gyhehYI/vAAky4ANrLYxam8JiByXmNkfdXBKmFHRambpv81hCkU
u1Y/h8gZvWdv+FMEv5/964HdWbLeOmFaZdIzox0c7HnVG92U3XUSTXl/lMPXce2V
ukEEEQn5actvY8R58nRlmZ0BG/Bclj1/sxBR0bvs2gFTa7OR8jge88W6OwNi1xof
IQKbZ5+tB/UJ9ry0Yh3+qC2rr3GcA7KiW1ndwSCd04xlTvt59XMnMn6Wp/+Ic/vd
4c2ITWOmQqT9ePbYkPK00V7MGHm7VjDCnwceXlCp2EATJqpwTSErnMtFWSoVFPhv
KyF5xstYbMK5aCbcYAgq4ANofBaLkAAuOILZnD6WdP+x2jZxgt3HitYC8X2eh4Fh
ZnD8gzRDd0d9+//FpMCObpDI8a1i9WNNb3UedPr91bGA78Gk3kUiwkQYI3NuLrBU
0dzKimuaTAYBAz3wcTijba62xZ6CkFvVWpLoCo4glewDE0W8f3cqB6TTAG0SxTbA
tQnlIue8Y4eeKAG11xE7kRfwtj7seRQKsmY1hnKZp/C10WbFyFkwNnTvMBfDrx+Y
PJeb0VE7homtDmlawg6+JV6bSBBKj85w1u713npe/9P4yPqFZQl20xWJzG1EJuMG
NXaZvgDyi2zs7EhAtLOrfo37xnSgveUiPRknMbf3ADFPmC0XaisG/tXAaizsgc21
mOaa3awzR0ZCgitre5cDZQmA1aUygHZRGiwTcQafifRv1++AzJVkI9xOfI2QPJOx
HuQqqr2KsZjfN1J6v6r8bnVitSr3gkt2utk/TEwkTf+KWjYRBT3ecFrKyaZfRAaD
1OBcSu6C0X+wUlf0iZFMLUyiVBnec1Ya5bJBp/t/vH1qXGwoxX+/zlRqrZBS7Rxm
qcBZMNIQY4m+wTLwAlBvYJx1gYcgDLo1XyLyjLiLXThO4HAa83XQM3Aew7lU3JZv
GXM3uNkOBkaWowdKlA/7WUuv9b1t9yENmAk61eoNJbixmf7L+g09TDBz3VP8o+Et
xbAbUAIepHq7CbKl7YvUI7T2J1WfYXp9sBckdgP+NkMJ3zEs12Kq+ciumDdIGZmm
f/rCSNHG3Ty3u+4iWU+Q46OQulQyUYDLplAeqYzOKBc9txWu7Draqtq3qK0qOA5G
lhjXVQitvyAF1mSpqjMYJqU9cbnx7cOsr26ygRphtr9FojOIYi6WO0gYsYna5unY
YBCVbKXwxnxA8Gbf5ulb4+GHIY+m1imo9MTGSJUTIRlj0+JaMW+gAxtatfajgPtO
XRUvUwR/CDqvkb3fH8iTDYLLXdsIzjc5UgXvN/6nT/UOYFdETRa/SNz3cROLveWB
thSdlhIKDF0dgX/h+Ocqv6PUvEY8CN+hnO3HqzsKCmGxmqA9gUx7fcbVLQH0PpoC
3FM8xx866Yf+rZovz89qN3C3TgLGyGCxVaY2G7Fm/UdRXnFhm80huS+5VTE78vws
xz4vkDXBimD+jZFMfm9CGcZEDwKpZdPEtacm/n1ZGtV0cD2m0g0HePHDoc6naAF0
9T4QbyV6yw9+HPG/1sDwd/iVP76L4C2fncOVwHuNXILjId6YD/UQzMTRYk1h9+KX
527iDMRTsZGaMxj9Cq6aMeGAXdbJGsoYXdlZCKzWwgkDocZy0hMqL6J7pr2WG1aq
khuT4pbZhbPCQv+aeKpoKpyPN8Xh3EUZEdErkeanPnS3Prwv5M7EaSyYYNo4L3J0
4PUYivC5CavrfuUUa3PyWmCXNa3VYztJaVlLmubGE9qvai0z8gSUeWzqV48U42u1
UYK+2xqs8obMP/h4KW9iWsvBnBWmN6e14PzxOLE44sISJbQ9M3iUxWIlWCvAudRu
7d/G6To3HJLBV1uCR/6zmdM+z0lUNdQQVxuusl7ig2Z4j5QFSdalla2uo9P9CfCj
fmwJBhuU2zictnv3WDA+2F0nnP1xjuJ4hAchTg5XzyNitOFqzY2kr8ljh+Sy7A2+
QsWdcKWbNWRvMwUo18OFnFuF4OtDndDEBDQKjhUyG9qsB6GoscNEyEKSWVwxTvYj
XClEcO/dkdhzGH+yuXczkeTr34HkErpsdUsn85t3qLHkcRKH7U7sId2GInAxxDKv
BCht6Y14X3INPfwFt4ApEdEYH3K01GCv6ZtnkD4h8RZmFbo0yKzhbJPpnqFn1+vK
B+Fer2GQY0urrWFI9PD1DK+Mg/CGAmFKQehrAz27U2qbvwNv1UTNPKnqFhS942Kh
b6s5xIdFyXGrhfBcaO8Tcu1SKR7tapbHMo851ai6n7QwciHHjU+OoB42yOiEVYK0
50WfNSWLx+otIQ20/BLiiUWIvUbrZi/BZJKBe7qildidekf+fnjHFwIVg7yq6UEh
9PA4ci92xd8a2JNch06L/x536qFwf44XlfDO6KOMceTH7bEJLVnX4mY7h5fA1lI9
knClOcTqJ2v6F3VpwuMYbvwoqgZSqQjAzf4zML+KPg7KhEtl+mcJ2XjA/MByQ9ve
VkpSAl3+T2AlNKqEJPiDn28V0T9P84BJQYHaookmBUS8vCqPqh6IEwTyHyT6ZD1V
DcE7iYjbK5zYA9O9xn0qKjy+6OfwwDocKhm7yzLwh4Nbxn7As2gIBPK/el4+PMZH
+LTRzgaXgUZjzAIvXnz8E0nH0tX4ITxUlVWugldcoU9UpR3W+QV3FOy32Zvn8hVP
qbv2pFPYtRYKoVKDInktfALqG/IeZX3d6Zh+R9CLGyjTFyvzi2/BxL819Ych5z0F
pXO8xe5OhQYgiGTuCRPilLGcBy2nPKBRaZVwgs6Z/DpOegkN4Oar4+gEqvmADwrB
SiVKners24d/J0FkmWIUGZW6O9eWeMuravJtVNNcHSUxCQSEZmEjiGdXDkEA3mIQ
H+QE9BF/b8DqflSc/uHLGGFW/kPZQh5Nb3oZvuPrqSmDqngIWHntoN3de1kEUfmy
yIrVd5YWPdvpLriIxVX+pEteWRnx4aa+pFGspZCCHNM39lHveH3q+CjisUFQNukE
4eomZ1f4T33y6KHYGBKBg8O9jKOR2ilhIUCLy3YfqHAscul0CbsZGaEFIynY2umC
W/bpFDKqXPD9A98hwKQRAm5Fdf1yVG+8h+7cMQxU/VNs9hdI7f3un2BubK/fVABE
FHRdU/JKteSVcxR+jsCkKpOjmkuScTk43knHCHfVB7YyUXKQhrM/GQQgxWAAewNb
yITjcXz2d6cTv/LWEC7gSNxoeAZMfeep4zp/x5vPW2Vh1zdW65UnE7FoiQfWtSlU
pYw+/GEvC3TRkYNn5a47icO+BnSMt4xejxpXtPM31XvVzq0BeJcbPYecxNHjc7Vx
YD7ZweNH3e0sqdx7lY6oBX+XySruRNtVAOIRT31FpSXO4kZPKY1/BFWCkJ/t9Zc+
9EkZMs9S2/kwQI0Fif/sF5wNs2fPZE3hsLO0QJFUjXZ1lFF0+6PrkYGH+/iECaO/
HHlUiaQY6AgEvmG0qJCkl1fy6/YvHD09V5u8v4n2EB2H1HY4L0NdVzX6PIoecj3z
jc8rsBAxnj7RQdlgMYNCvskUFpIobkDO3wJ1rZAfZlqincUEA8XP1i7eTQ27Bwbx
PUkGmO1ip7QtxxxcS1TSArWQ8j5HT48kmS87+Dovb6VqbJsfChiP1Bg5FhCY/FMf
sxGe4MrtQvNY7ag+52zT5uvOhzTaMYtKR0ZPmeIEUJ5HuYnW7z5ikjP5dr5I1qYA
2yCMNyPF7IUUj370LZpe29l09Tmxc/l0wJPi3o2KxLkJhbDvK6ssZs7b6HIkQf7D
D51fahBcEHXEhYUyw9dg3ZgdME8ZvoLNDNKcppug5Mefp8WElamOQehjH6cP2RXe
k1RDum0IIk4z9/tN91QZhAuYgKK0eX5OPCX5t6ojeSdgXjqCouWpd9sV01IonE+N
gx8za0u+OrwgVjt0q3cPjx1bb6Iovihhhu9LP9OfdEQD4lJFsl2ot2G6VAH0ayfZ
0OJEh4ik98GgC0keR6Qii3iULrK+NRjX6mAx5r/hp4lqRkwUWD/iv9KZBP4aDgn+
20sQ00tjflN+o2N/hZjSnyB4y/Bhj26VsOkfoWuG4Qq0xygxiAxly1LRc27aLMAs
sRXczq2juBnVQByP1ybymFQirE6B9uz0jCU54gOoZl24/BNAlxd88xB2gmGeZJeE
kptHa3KaGgXl/NfZOleBsnyZfZGACKocIjrO7q6ZmUiyGFOovAhIGiDP9SEjeuts
w8dXmq5pe/yu43XYgQtHwMIZmS0+BcBC4g1MfxxT+1X1c+5hJk6xAorcx5S7/StG
nQBRKC08XNP5phQ55GUlHJJ6SpL1ZM0pO4+2lgM0UqjbxLwmGzv4YKY4gZE4g3zW
FphLaSnuCDYILgAt8JS5rdpGCLUwqT3RYunVbXo9hgPrqHxwJTKTogddL+D9vVGq
b7V4SNgybLe+h6HZLz7/q+5NunDoVjeesKfcHNHeT278RVKt8e9Snr7z+hGT4k7/
TcDwFqOc6cdN6AUtqzSYeiYol0XVupbl3nAKAgi6D9WlrSZnE13RGEVp8s7xUDAW
vvIhGuWZmI9/WldFglzOnXbJI6qJW2qWkz0sHCs6JBJsfo85IXS0gaCurFF5aN/4
AtGFbISimGqnriYTMKyU/7T/DMY195PDlKZXU91U+9jlG++UXhXdKM9IVgikqTr4
Awpde2UGhJFE7s9Hm8AlnPkkzoGSdpei2g0dFwTbYaWLylQzV8EyYp5UaV2xOrMK
BpEe8AtNqaukxEeYzocr7paBp9kLcVwe8dqx9hxxLIsxxs6xx6BzCSMGkMuHo5h0
xKM3hhCjrHteqs+6AaMIDFqB9AZ/qT0Ut9ToVzLtGxGVKDaqgplnWlz0R2KIMXEY
bPt6hUWn9s0XoUv/VoW2WCFcHkZpe7PUwZeBHwwXcfXIKSc2d3fYi/9tzHQ8zLSg
GTUyqXu9zxA0LlpYnCX14PA1zN6N7a7bqY3TnHn3znsRzPbjcQFNjlB3zP4+xqc9
H8uh3PqX2w0JyKcRfa7xJfjQ3Kd6yjv/XML7LF5QGmm8XYIwPvpbpGqIrtSzye0g
0tXN5s0ZGsyVShNqShCWCw2jmyfh3o6hgKyeQZ04m/TOqmGT7JO1+8Cb+y2kF2nd
B/OZX3+whfvVg9Ivw9GkhrQpxkGOHX7a8XfYpnTmGaEMn1hKBDXhT8XtJ3iEHQZv
xULnpS1o0Rq8VSqpQRo4KczIN+7weINdDNcrqpl5hNQLm9zKfEE7dRsdZrUaZbcN
shbWDmxQt5lzqD6KqwoqpSAyZoLU020/3p7uY7PxK2HLi6FG9/lvSPV4U3Uv/U2o
sIiYvs7URShya+GrybcC4WtWB8amuv3arlHI0qLCTE5Ckl8LwvhRGl877rom+7h8
fZzPKgea6Tg6HvYhY+8H19lQiVcDQY/TfMLJJZEgmLPiTPkdewPAszJfs8J24KUJ
fsgl5TuMzzalccXXW62vyz7KCCoGAl+i9Qxv01k256uKRb5dbRidcxG9+Rbq7CKB
8etrwQ08OdoI31eckVtSnkkfv1pjotFYoCNUJev3LJh2wu2d1ae+/EsMYRO4ZYV9
hw2f6ye83TIFyv7UkKddIS3sOLSk1my5WypWoDgoN0fyaIvN4hDDv/jMKoX3BDpj
ReozZdwVh9ySsoqot0D6/89Hdsb4MyowBNQPZqOM8NQiR3KSuomPQG7nYlNMt2Cc
HElfaFR9VNYl61VP7ijRCEI/xlb7U/rAZzkvElHS7cVS6yoZ/oEri1BqW2k2EFGR
4dIaTf9wdE1Ag7RI1S2AZ76NyxGiFXg5PAl2e2ozAJk3lVdrnkIoXEuUReKgYrPd
ya3jpozQne9u8ruA1eit4ST1dQn2cQR119FNfrB+LK4s+i6hlly3r4yLX+kmAdVu
JDBqQUv1PjPTwK69P2PHQ/3QaaAgZw/8ap6WJS9E5Nw8oPA7GXIE0ElK3/orMSDB
xxJ8DATX42YWzexjffIN5XKiuTf80wpj1snjnbiC+QWCDsOABbh9RjHl8dmv48IW
FBwGH6s3/VQwT2+61m4pgF3j51WL53WUojrkF92+kMZdBEoJ/Mn2Mb685EO2Yjgd
hLks1dEshnGOEownnIMHGplTRQ41kosND7Md9xbTKehGjA2AVO4l9gWiQ4zdO1lV
HExJnh0S1BHkZzIqBzjFSgLHMX2LNuVkCrrtttmbA7SeZYAtupKTy7DPCgNvtQli
DNwc37wncqtlZVOZKkI9ebkKHBPREZYumJP86Y/lBDRPSD3HhzOhaqtYF/1Gzcb2
093Li7rW1O/3AOek2QoX5aNfxzLweVUwZU5iur4W6Do9uEoY4Z1Npk5i1fcbTWgI
sBCMg8a59PhpkcNR7/cQZ3+7kVngTf10vDqrcj78bFJ2FLi1svKQc1Vy1plx6Xc3
bQH+HJ5gctECjxKE+0VMSrhIw6IwRxotXrqgbaJE9hOjr8mZZDSx4pNVXRaP7Ktg
dwafmQsQTCYWN9WheyCjeThaMmUhhTlx7rdeccb0Je3NjAcWCjvcMa1NcnhYgpga
YCGsiYuZBgs+V9xyupHohVj+9aFx1dnkvVzp1Om0FBWH+xoJUcI5D9O+I7kskxi7
QLZaajFmEY+pskl9yeY2/IO/dIGgKyjmbKetP7DNxWAFWsoZsYB/4FtkyKCmdheP
nQvxDWXvjPZepm9wZh+bcgMvlBwlQx+ZdMGHAJfPb1HkFpuD103+aP1PaHghKHGj
5e8LYMsqABf3QXDanE5EzlJU/ykYYJaHn1+PhM087MN0VK9m0J9kdJ6+gl7NtGCK
QqhmrMOR9cR8ZkddBSoEhSmzYO6Mi0jm3fBY9PBLOJuPCij9jn4kwWFK9KjB3qwJ
JrCW/E5cmPksYqwLWZcvWa8K4Q7nCoFPUuuRsw8YZS2JaN8elnA2Rs7rsDg6V/HM
Z/19LkqGthSS8rF4qS0DyL6DD27X/FPsh9yNLhyOqA0SS6eyYy+dE2jsryODUrYp
QAVFQ6zpEbEveQ1ZZiPE0C2R1IvuRMSXZEjYFV12H0Y3ls/7idq9JuUHXVDezVHJ
PHMjs6isEI4u1lhjf7i6ROjBhvVHGVa7oR26hI5SXlrU4scX8GL/T3JFCPWfbRhi
Wiso2LD1fywabvB1STrx07g+HM/+bKzIt7siaGhehjnBJxrkOy3K3NORjJbRkGcy
y2vrSGmuTX5HmjMw4/u52IkpZyyDK7tam7axzC+42BVe3fdhJrvZ/p369RGGYqNE
ww7QtofRQaU42l4DkW0I8TJHstna4NCirgI8cyaF2S30CiO6MyNT1N3T79j1vBbW
wgAGKttOalin9Q1NPv3CvHGTc7RtU5xhI1yEUCrG+SRZN0l6Mt4vKCjTIyP5mAXx
gkqRPhhdRFhvWffl6NeDVlkLXu+tfqQlERr9te41CU8gKVxG9T/hYbls75kIN9jz
oB3dqixJUeDMoAOCOSaD9eTYM3MR2Zvxo2CkGfdMUlgigfT6m5OqBymlQcOMCKwI
CPNx1llWJqoGj7Cq3jM5BkiH3CXfHDfeIKXhIewfluuyLPyGP8EZJp32ByqVpqPI
P+npauGDCLUudKaTG8RidVQlZSdWiEVqnE8UOON9RWHm9Bjj7xX4uEWS3rbWOtmA
mHsantsDWW0YsPSyVlua9OLkTrpNSJn+PR0BQL2AWibdnPaZsZEQgywv9deSRLvh
6el8JSD3ANMIN0GwjOZSIXECAGWr/YThtUmuc8z3vjcLeHgh3DWunvidQMm4660m
NUR0JmptujJBvYZzY8OJNQha+XedXyTGt+aSQqAovOkMJam+J12IsqceW8zVQFaB
L7ASc1tJFsUY51p4FwLAqCV2IYzX9vupty+423K6fhS3rlTTlHUf8plr+jdfZgvT
gNieXJMj+AFACgSzkRt8MBZqga+Hj0wX2fIAvvHt1l1h30R8ti2rs9uRzm3weA4A
jIVNKjiYX1oeF7Wg+6UXcTtPOG5uI/p1AkOQbFxvtaJR3e2TYFN6S7Efgm4VRmSL
JxdxdKFCYYu5l7ct/VIt3tKlTVBVIGNhUaMHlms0Oi2Dt08mR0Bjw7ENH68yFWpk
d4hfJswtrmw7eNXrFjwpvO+2Fi0cfI8ppttfy5iEfmgdq5bkuy2KSvwLYiB9CFdf
MPRwo6izMc2VRlW/vRmlvnZRbyPSjPUHlcgSKrnOx6c0jfdAtiSyqQywjFKtH9G7
S0U3wxL7mHuHFPziHM8OIih7NlZLDisgZbdIoxz+DonQRe6M6BI6BEwxEvPy1tb2
UcOm32iDLiMlapZOIZUgdSDB76GwX0Fm1KUeBlAV6C8FNp9i2C02OEPQBcmCPzM0
54BIqXFJBmqDXWBxihBE6AASJD5CJel2vianRG/gdKMqsfwC0rWgyQQuXUBLhldB
2TWy+3NNByjusQCrKApn4+wEiDmk0YQ53YUQS3iBPbtHX35boTzOoqNDM0eCzDL3
KTvh5897nPY60Vr8ARU5B3bhB2+BYfQtqySdmQ+P+trOEAhqxD99DyGYdbUEOLMZ
pfYh/iF1Sw+lCDfNUpr4TRZ1pMPJxmhOiRuVV5t/VhJe091Y4ve9BnZQBBtQr6q4
R9LieGXpCVs+g3rEOHATHMUaBRLlg5q0DFjcbToaqrF+O69w1RE5cd7Ii/nxBcqE
DcxsfiNXIadgCemio0O/Gl9K90TD0vOGa6vr3c8IZeZJjKOc1qUTSauE/5KbWJM1
OepV3eg6MbuNvkhGJ/+AegjdpMsQ46+ziKOX5pjtW3IP3MZeXnx1El3fvP++SHU/
1/MMeiGc0zGvmZwb+SGTgQ==
`pragma protect end_protected
