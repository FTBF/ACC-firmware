// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:46 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ruFrDqchWcOkkdqaO/2YHSES6shDtnv2ReeX8UY/WwZUd1ePsoX1A4w7fIPcTRVb
ssTlcfKFXjvcsUSd3mxfc2vJa/NqJoXlISsHYJJnNFvpxv0iGIJslpjSlC0P+e1C
YPetBgJgeBpR8b2ZT+rwFRetMCabjvJO+GvqNC+MImw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25648)
0N3iZnHM3qZF4EHTP2t7Oia6FJ3I7khnjQ6c+KEc+zex2uI2wwL94hfGZ6RYfV0d
dYoSlxxXI+mKnTO27b6hxkXzAl4LVag0Z03Yw3/8jG+QU7S0Pkvfi1pbJnpgZ6C0
gd1qDWCGXB8fTT+b5Gl3rURXHe7J6i6rEO+q29nTpAPML10T1AdAXQpD+DlfZCSS
Kar5/WrsFINjGi2OHSHCMdc46XI0KCS2oNBA6ceJImUzgtG3/vRjjg8r8EvhetKQ
gv68Gp5pPs7Ndojyn6ZQVByf5eqFqnBb+oKiyY73653pXNvpYuqqc73D1mR36hkd
J2NbuWppXOIUkkBvkB2bwLe1q2y+vQk0pv/s55Hc/ERkO+aBL73udvAxwWzoaX0E
ZQQ/YTm0DWHmYpx4D1saIMRCFT5NIKTm/Y8KXAis0v5NDLRHc4TiFiITV68El/qy
Zx8jZKko8aFsK0rugM9hOyz4hlyCMZ4oQgOm6oNp/2YJ37EEKh42cxoTCZbObJ6y
VYoJGam3DJP8azm0/3PGxLJ3QTYx1exgJUBHBOvz02BS90532RR1xUbWuxiv6zMO
b63SVp9gUX8uZBf9UaubNrhgz2Za4V0wqtfz8FbELh17+rFzJvWKjBIWoXNmvz1s
z9pgrBe2Z3gO5f66KuPq6SkykNrNdwmUC06iSwmYMP39wBDRvwhP7cwnAkUdEdma
H42ViJOmQqRSIKIILL0LyDSG6W+Uwwf7fMfZFKlsBQz0RYLsmQ/jTBP3jOtqqpSW
1IM/TkISl+dgQxjvHNQ/yGjpQBZ3CEviJ2D565YTmpgbpInC0s7obudJyN/3rVRY
9O9bOkoE0VowcJChaL5THGDL4iTzkxQvJdcUqj69BfEaEnx3E0+prxqyEF3otI1O
KYvOkVQ5hG7wiNjG9j/oiEE6lZxod0gXe3BuTTD6il7V+kU/8DLOYgrX29rw2S3u
W8y5fnBweZonnWPn2VWm7Ih4ZYpjZd1M0zkqzh9H+k0yDQJwsSooKSPuu0s/B903
iPwcRhNaBomtNS1yQwh+/RrWl3LYTVyiZhzrvBDDsiHZHED6MtD5e6iVHCRkrpSw
9xxv2nu2Azn3lvjTnQGdJfXuFFyAooKqvONQjILiF69WuUgbjavgvzt6fmBCW3+U
nROoHGGedqaOPF/to0ZAXlsjfu37wIT/dy30HqRGlddwwNAjgvXRuk1EybyTd2D9
L9VUEMIrk2/fv1IdCIbJ3c3gzmpZBW5BhHVgpUYT8bOtIL6CTugKmbaeeMSol/qo
JnUlAqopp3kmJpDSrY7lg5vLAJo1w5mbHb2HsZDYPMDvQlgwZs7D7WnNgmm4F9TM
b+FJCmR0HHW6q0//yqi9QKvQXu4RpkS86rHNrAF4N1NuM2pJYQwnElRqQhSA4rxr
BdB8Y5T9cAon/pb1JWJ7xPRhrLB5OemKPZ1typ7R4h4r66rpzEgz3mQVASDJtxAp
cSXLBHSGBdIfbP/SLC+dXtthhZ6dJjZcJZ2Ue7zfSnKJcCCht6a7MoVTNg2E1aKq
s0PemzrXF0Pec6k+SxP001w/g0rR/V/I3RcM95X3AlgzSET+nJNOgtCMKIEWt65p
nkmyiGD6lPjpPG/3CtStLn5Vwxb1gNJYuW2J8BHqjigp9IJreFn3BuAgRc8mn2IT
14OGrrvqQk1iQVnUdImVq/PV7P0WTO/KdMJVGLLsfJFVfyo8nlkf9AN4cMVPMZhr
ARSq+YEecCw03i89NRId7cTLW2lQu0l3TTYbFFtNMw84t1B9t4NqYDCGZiv5GIHU
5twCO+IcZJtL7ujTbQYTw2vwrGs/LaC3ztvNU610W2td2K56RLe50ccp8SW0hGdZ
/4M1Onlr1fQQx1APjQuKTMoi4A2D4bbiluBEkA6CG0bblpBxw6vatiweMd81oNCi
0ll9NJ12XiUIZ5TJIr2s4iwm/kz8nL2ggIQ2EbOwiRi6CzCOmfj7ahja2yCFIQxD
PRHu0IJSIzjRcDEJ3r0uq+8QNl8/VhZ+aHhe4IdSgU8pTDy0G8kvl5srPkQWlonI
nNnsOqay1aJCLmdPhVvc2Ih6IHlCVkipyAeRHPMN7tf0TPOlbdo7x54MhL8nmQCy
1OiIWcRU5zRMtx6U8ERIaxLeyOnfXeymXYzYQK+JELF1qfiER+FcYeYOjNKrCtui
5PM31XmJdyc3NJ5rEwQKfQKUEOolOWCQKjj/ReIx1/uxapoa9uIZUnkbfqLbJ7IR
hJoznWJJrk+lVDGmwqY5e6EFIUN/vePDTIAiULd9BkiIR03kdjmyCWaAAvTsm50b
b2SYfUTBvIq55rfc3uvevRg9kyCZkhPFx67FfbjATLHMSjxebD2z20LdAvc/V9Mg
0WoabovUmJjLCCE2/JhWvBGfHQkVRUKxpD0IlttBO6Y5KNlryxN0tSkcfaME94mP
YlLr5nzFDsUC6ly6x5ZhLBdQ+XiynD5NAdtkFiw2EfEUmpiniXFTH4WrmmT2sa6o
gFe4thQEIl1E+Q1bUvsqP3E76vrOg6dGWFnLtG8G51fJ9fHPIeTcKpl9MmFHMnSF
dFNhMrUqHJYEBluSijGcNtxSjj2/aREyzn2sHXvzuU99Ysd+8RF478pdmKGfO02a
G7+FjBm1I1GKgKH3qhRgZyA7NYMMHEx7zBF2W38PtOiFJDr8ZOOT57DpsSKN58HN
qZQ3jQuSoX1BoCDUXsT3VOz3MqL452h44vy4gxA+e3FRGPCqzFqoqMcvUHec+Gop
oHxzgfOYmD6uZGh/2V1pySayP+1tidLzrvzp+HXxC66N63NA8xoysao99Lh7uDyM
fkIT+mQnamLakSDm3o94/1grewMn4ssp7I0KXyARIOE5kLwKfZl5MrPfP65xhY6I
mhZMshQLIcLdG34VA7h5GydlUPXloIGYAX3ck03UN6Q7qx3+4xvoZ4tt83EesnWo
mfwyNOUlWOJ4vlEFiwAJwvwkkurfm/aOcF8HTkh1QEIB1LyrGTSURDuxKAy2nfo9
okF+3ht6YX9A8PaKZQpAMsiuqbnzguiAWRjjAXDWOIQpgO1GcNpK9a6pWqYqE4DW
qZPYfm3wI0BdC+BbJ4keMtT87vEvcVhGN/SMmylXb9xRkw3mqOJLA6yRctq1kZKc
iyVMP6eLAxwoZUyUad7v6Q6vwuWO0fDfAlva/G+1zT32hFncHgiTuw/jefG+7nJW
LsRIj+FszPhuaTMNHhvshvKSt75dIpENSHAZ0c5OF9+5oJCWv0GfvwNa+6E4dLtt
Zui7BEY/m06TEHLayn2p2xlHWxNrID2TqUOSs/OoXKBed+bmqJbyMdGyO5wWKlwQ
oLZt0YqO9H5eCAV++x48wxVPuRvPIhZP9ejG43lq3Qz6K0c0njZxoKEQ2I8fzGuV
LxbX9ZuIGHQyu894FiF1rngiYqbRltKK6vMbVHiVDeQvnUDPVQ1b6BrGxCsUnlXk
/J9/FBvoJ0sNl3d4VoDMDBsS5Euix2QGhXAdhGppbY4FSywFoQxqED0n9MkgiqOt
BqBcqU9dxar51WiBUSkaYSvunrxEt+b3njNcIzjgC36FZZxJwC+eBMh6kn5krrxi
293k5joXUqhPXfIAT7uhXUtv86+DFHOO+DYGHz9PV3JyZXkNZmPCB32RpETqvmZt
xRhmMIZa+oFDTjLxFGwF0r3P755R3WNKMhguOpbNpqSl1dDrFzPYMnmvPqunVsuo
0hu9HRfAxJqYzmp0de6+6DURD2pkyCV2nwwoYem82XAiUfQNqhA4gqg9tZLyZQkf
iu8go2TZatShG1DBQ+B9qOlJd4NITDNpE9Pwx/h2p2XTGRY+qkesTlIlHotkNEuy
QDpyU8KiE2lLgRltE+x2Rj7QJ0HA7MT/aN4yrQ7xWJtK+Row7yeGHjN0yg3XGGS8
ZtSWNg6kzq87/kIUPIRN0YVp67BtfkwrgVyHF8rWosabHm6v11xUUOQ1v2DWNmho
zcEkkrkz0XdA2FAAsKNC3GKsX6sfo8Ny3kxYlKrjPJkw3OXoLtxpPR5NNBu0qDcy
oONpZ19pflXflYp5bpY8UApTXU/Epm6oWxFDl7Xf/m0AwA19Zh2xrMo/F4c/kRop
5I+KRwhO+i4dFzwoOvF+ysU9s/DekKQG7QgG0N31zAm+SvZECVrStbFTjOxBFvwO
NK3gU3cE8v6w8582y4Lc0dD3UfaLL42Q1ZVRn4fZWI1j2468/Bcdbmg/XgnxfRtB
IR1MnlAC0wvlUHsmuVzwPXESy1YalZ2gUvNhAJd4Ju0W5WXxNDAiTN8JG7/WskVs
FUI2gz/hq08NW/fo97nzqNSmQkMepZpyGU45B1+k1iWu8FUjaxl6al8hY8bvLt8h
qMZStweoCpZJOmQ4ouP3aj4RwKT0qvEh1HncWoXRAI18RR8XtT+9/kbIILLsZeUF
oZiX2h3ixbyZeFVfFchQ5vjX7HWKJtFZ74UnFF2cXni1dPfpUICjWwRbycDL23cS
iMqeNdqStXrSuRAIOepBqAoEEaSMp2uiQmCcV06l6a0Tp9GuDTWyQVvFW5iXk1Da
jVDG0My1feYtapaJwWc/06G29KZ+AAEhnGUr5Oy5vK1060ATHvywze5KBMALArL1
J/qspeQ5RVE5jqSikW0VXoD5bcKGtYU8lQ1gOjmoB45hXeKOg7ke79K3NaBT/C/l
KJufsh1+nfqDXO5xtFfqJsRg19J/DUCQe4dDv5ZXLkFLV/so2l4o7lGFQns4Jidu
kLwMvgFD6TH311U/8/3m3zHnsDkrUTSaWDF76qqE6VzUjtq55xlUyhZrsGpgNQxv
BLvsvIvhbHbCjRHn2IhJhnaINXfIn4JY7mmjbVFaGwqxJJ3tSUjYQP9kc+p0bjxj
62K/dFXfTc1Cdc4BNilggNnEUaSCI0elc/LgXoT/pF+g+i1K20AvlkL0VFkvFJmj
zatOIfhpspwZP1+h+UI405/jWzwgWi+Gj0dN0JjqM2+ONfrSEqIeo7wKCZfBzVcQ
FVhbveY/r8GK5Tm8Cqdomgtuh2pVYE8kxY/f+W9rvpH+9P2CT8JlEqGHqEVpX/ck
3/VJ4mQtuiYktpjPSZDuXpnhdJTOu4me9GZJW0mw/+Osmida+tnjdOtwn+HlCF53
aHEgA03S9GAYAwrrVxJVa7OfRolowCbZdLwgELtPbmeIzpVEiyLk2wqRHxNv43bu
jN5E1wvoJX90LHpaQfS4GWeNmVodfLhNGNIHAMImhdSP6czTLLhCLpwu8nt7F9Se
MiRTdMoHR4E9NGoDfmaZdciQI4MKzJWe3GiR+co77Bvm+sRhiwTEvudWkdkmeafL
1znE/NAm72Hrov8xLiAfKbh+RAetTuu9NLhZoxZjhvz8d61pxMIRAmbfdefYJzLZ
wPYFtBILXkgTomCoiZJmtnoU0+3+CLVcCGKlavPE7C3QbsKm39Qb2yfSwGm+Roy6
zgXg5SRn6vuE25TZ1qSJRtvmn/oiVCK4dn/FDo28+2zYIn+jxkJa9ggbzNeknRyb
6UIHuuOjf3oeSKzlhjsBVXRCv/boCbvSfd7OIkPwvwmDvUokniuzq3zGTt4E9b8n
CjHKqyhB2e8m2lJ5hjD8qeJzDkn8UfyigO/Zv6CLp+Zq+q6+SDxsGD74FlLiOqx5
iC7SvT/EcMrgdxNWuRZyxvqWYaKFlKLfZb6lvulCTFD8WbJJA3FstfIGNAWuQAFe
1y4Kf0re4JqkeKuHaDFveDWsaCC/uvEe37AzyOV+PyYPXhI24aboSi97sW3pciK/
DoCtYkTCXnEEZTaNzJNB7d7zDC/P7gFmLb+ZOqurQ/RjleV7vlnx7h91i3FzbBuG
h1bud4joM0GA4fa6RR8KCwjyFvdzNBvkbch4wMx7q4jT1bL56wPl/PJnc7EhLY+0
dy983mYWzEDqQmXKPrXP9HHBOLxshu94CGv/H5vynGzmo926vIv1hbr85hAX+fmI
6Cpecp2Nd6BT6vn3yYOfGNRRPdCKlN1eSnLcNnB8gRgjuKQCSR8y+5bb8dz67NhG
tJ9rwbwoB02ctV7891oruXKmNMl6RPpMsZHMBZX6iVhqUBuSlno1RCfYay7FCJHy
gjwZmItr1DzVA7PoM7IiSCt+zSJHRfxmZULgqZiwfJ+1IuU4TFThcA+xmQKT2W9K
e1cVisvXf+FmdTPXdUMPkwEFb2lUfDW+4rHbDpCJw1NpJ1EggGd+bwahXWrVM0qa
QTQT8YM9BIfHjNcBNUb0srEff11itcvBRr3Tm1VHEb/QqvpSAwT8NHAHC+wbwK7h
nPyG5ottyz4EL13Y+ob2tCT0zr1o5FX6E7kHJQ8DNvVwa5+2+oq/gddxWAL3EKBW
K8CrFS1DN3LkD+84n2mc90EKzUXuXiB4ST/SS3/KaYqJJZrcav7YDGLBpY66vF1q
rz01TJPH/CbvMINILOnacLh0C6fPmACAVfjorP6VjqZ+8/9HAOEVkOBYLyc9q0gv
Dnis/YEM76t6N0t8bO8dwcaXoYkP24Q1sCBtFpNokYrwGNkdJ6T4K9VLaS9KbtZ9
SnyNHV5Ww6r9OONLATEi6jnAIoq2BjOy2EpCUxmoWuYdyUDMMWQiWu/57dH7Mf6h
jxjxb5Bmdno4X/CutAkFFMmb6SSn2fEgw/SnWgivpLN4UpkQVSfKmrCaA8lSVULz
e5qefo6GCzIp0bA2uylg/MvsjhYz1vS25csiJ1v7RZ4NMM5aC4ENRTn4DophnwIa
VFdZcnbv4qcpcdA5VO0gDyY3slCuWlgRv4VohGRw8Pjh4yOhEfrd9sWx3PmIbCZ0
C330UGFczvqchq+CEcxQ0PjnfJsmG3jkHDOm1UpqeP7mDDxosacbQH2DHXIqxXq6
9gaSKWGkS7ZOX8QagB8Le3vMJDKsRvM5vh0TTyCOxP1YHrwSD8Hdwa0cBtB6i0Ku
VoUJhQ6DvTLBlq5JVA1jCq6IG6xUfO2D1iom/ZRykd8mYnE8my6wqduN/yDGvg76
bGnPjuGcLraiqaW5JwP2/7kKWGluS+i2dSaeXSlvB5YSYYg1Jlf0XQ1zYsMTvcJJ
T7LkHMMchiAdf7jbl5CrbXJHcnm+ulbHKzTQM9FoUTptSnUjzzzGDl5WIq4w5yBr
IPhwQYDVWYJZzLz2wVfeRbI9Dt91QwsQhsh2W7yeYtIaqCh5yManvejKtGwwLDgN
2DdwJjI6MHSqfKCwF1/QjP1LlzP/afmOiOMcMOM0ORytjDt56nIN2ivP1enQItEW
Zcu4F/jeBRIZZ6kgjrfzvd08kopysmtvdUTCzkU54FNhFvXTGrlgec7k0wh2mcO/
7LfI1IuE/K9IOq/NBAU4+MNPY9ByAJ6/tDensCg6B9mH4MJ+IHxLKegktNUMoeCL
RjHBnwRC1ado4qf4fcILjhzrvH0AkiCGPv3hXSS9cxG3O2lyIGI/H6Dh56GCKYFS
JnDcdU0SDMW9N5Ji8FKyHxxAHExB3M0ts7EL1L/9MK6/kEGm0JQvtKPvjPKYULK9
80fl6p3OAwrFYR82QH04Z1F5ZqUMEwK7q9P1lWcupaDdifHCB8L7SkwxqXDOgW/G
j4Uo/zFomidbA2BYVrfFYbs5MwHC/QxfQaIjeLOSZpkf3eWaWrhZWqpsGvCi2tS4
VP2T1hs/m60BAzeGX9KfpzFQqUiFlbb+RZTnz7IJN5vizBl6LXvPbY7MI1sG50eC
ktq77h6rpMP2mfADmzWitx5Iyfhs79NepMF12+PGLuM0BQLBvKc75CLjh/qxzRj3
f7XcBgBv2HfoQm/pXaMsukf65+8sZTCb0Rl+dwIX5IUoMJBks8ZBpQp/g5z5atQN
WLYfdciVO9UFZ1tj0tYcuFEYsGgMghBeGr7YzKf5+l9kS5uPtKI9gQG24jhPm9qF
WdHnBTsT4fxvnhFjp8YMs84bU4ZnZsjg7ajQKy6BZeaLPfg9agWBBHpSl9M/FYrn
tCrF8dkt25bNE3AkO9STqgfNnnMsYCFycT2NE2TRC5Nyn2au28tPmvxXdBZNEP4K
0AZFjUD84GDaJd6dJ6gCpdHRPHM61rC8wxx1m4qeJvnGCR08RSP9e3U4dwc2G8wg
5AKvz9KJAvIwfB4bXgPFHc6Cklf6Xa26o90P5GHGx1OONy+jmIo7MiyQLPLPqQCp
HVMEEgVFqrDsTfbDRMsQcnms5RgUr5ErlMMzA7h+OCfIU0Pjdc6NvJ7hAGfeRpey
psP81WRy5PddOtHGprysprfZ+bAUYwUabF0ELX1RT0h467i3d5zv7WIrOYnCIuSP
AjJYiB50bMekcSYFrNMsXQG7gCQMuFE6qNJP8+eaa6wPDmIEKnag/8sZEPWrgTaH
zh8I51OM0XzvYqG6GU7bsHSxSHJxNjbGZ+OONvhfJfW6OUrBnRAJSmrOjMkvyqv1
awwQ2SH5pms/q96Pfu8Gzh12/8SerM+P6VwHOrszPkES3S3IkBB6dT69z391XaUT
PB9dU6MCzPNxanyvjangFS3F8/G6VeNnRpX2leoHyQRsxdZTmJomzB4dV3MDGFgp
NkWdHM+dB8dQyS77ufePuFUZylpKCMFqChY8/djz2/V2g6ec72pE3dzrMtTxR+/E
16mwXf3YNxh5sDDAycyKhdboZzltznbUy7BZxiQO2Y1kn+H9TYuGlQiTjqFXYsAx
vi082Ydb4qZMdrp6jSqOxtcEXfs6OUYn17lCL8nHNNjqGJ5cH18gnwVjq9v8+PZK
OJLVaqE+3Dp0RkfBspEEBZ3G/dnP3OqCD0b8yTflvTxO36RyrP7DjqfLcyjMxyiC
rq4bmhJ/CxitbtFqdaGlwXB904P/9OmT/EaB7EJvhUHknVb0GZXCYtmXj7EREeLw
Y2XymOdjKQ6mL8EOxin9VPM0JM9QdZdBsAZsaeyiEp1EgUSvwQH17LwGEfN6MXzj
Py1NRrxM67r9wqA955a0mjysm1fCo9iO2fvy0qb/Dx/+lQa5Nu1S7aRl3tvbLZgX
rzRoKw1cRse6HuCC15pzmTOqJ3LiYJZVsLAjaYgL8FtdTY4UOepxg3ZvfOTc6uhP
CN2GWZHu1p/eZ0mRfl3n8rRV2HUkWPIl12ca5YgsQ7M6TxirLGq2t5xOyQ1bVxrI
klDcHI3eCS0HSdv45YCZe8bfZJPJDTK1+r+U1fBhEzN/Qs9vH3jQ/QCSKyUSVN8t
RJsDQY6ARDLLEgt/TihcRlvax/xh1y0WMHCHpofNYVrYLXWFEY8klVx+arGwZ+PD
TJJAkVG1+ehzfehTdnJTlXAvpoalzIZSjPPv6bGD0o9+tbUMhnhXaxEPuxGX3i48
lITKHMMgeeagePX9GLSlu9CgdsC3R98FhRpmt3QVQeZOCVtQ8pdu6RvJX6YMYhnU
Jy8uP2cI04lQe8CHoLuouHE1n5QVG/0FF4o7MPgRnIA7N476Z5GlwB6Mnylx30U/
ahS8PCjFXkKaSb8rj8lpgOkH6oaeibzKMogLAQwoxYS1MBJekr9vIUWZZlZVKWzn
SwDwC1PYu5z767JmmR4V0XipGP3RxVCoQThjlBB/y0Nz7RKR2QOfByg8yRn1OzXQ
F29iY7FKR0/IALONytkreF9JhxMKFFbhRBGtvLS9WGA6OWZyeq6wjsxd1Nfklx62
tWOSiMkB15WOX3i9sQ5kQsecHlDR6BnE17q47/Kcda42cwHPUJD9MdAp34ZFnrS/
mpKCOyG6gZUXGBtgkqkdUbduNkPSXC+FMmAdwEFrWuAm6n7qNw1aCPQW/fdaJBjY
PZkW1Ea84oDNx3vMRw7s65+NSMuacqZuqBEOLJSSz1W6J3x2BD5/AraahIp67NZ3
eERoPbvCJ0I9+8W4PLqF0bobOwc4FVsjmMfwhhrSW0dtRYnow+EXF4m0aqMEG+kc
Ed+kIimqcxD/L09Vqpbuic3Ojxo0WQHXtmwR1QPdkqQ7HSbYE85y9sQGmWQU6diy
3CK8rWgL2X5xe6cje6pTLfYw4YCjMHF8lXtEEGus6cAl+B0y8OwFOrOVitoyaQES
bYiKBkFuBlCjCSglSw1sYsKKjmp5F6H77dM59POmW4qtdgvy8t0Y0IhbSqH7OqWP
PuwYxsRytwAc5XbIvP49QEO7XDV92t6xLYs/aU9rntGQn6DKBni97DVK22CWVFOS
vjNYBHbQ72T04cMeAswJbdSZVNv9+N4M6vAI+gH645aTEwEepUDA0lldy4Ry6+1p
lsUlLMQGMm/VKP+IfjBP+aQosvm7elnG2yl6La4i5B4oNzubRPuLOGYaocT6TlqZ
OM1Lv3EWlvptdFjU3xgLt6gnGv2mLBrDwpr/5PAXbJXHeaZ9l/kR5HlzDXw6yZ2X
yzqEtc6pBvvlhGvhOdTzoXhhiy6pxcnF7PTYjC9Tmcn9ZXO3Ke4UhIwr5WzayC+g
ECVpv+WmQ+Ug0Y1F6PMj2ZWF7XAncFir3Pvf3RgwiLzaZEctseOOvDoBFQwbErEr
6g4kAd9Jlvj853BKXfy5sh7wmX+vqdxO2VySm/mA0vYJsbnLZtpub9Er7MaHaZJw
ISgdbmh/ZAj4OameBVdYJjfHU6IuXK/JrIRk2cbfQGVfWeAVKVlaOVgtr5fInLU1
woUjqeJsOvj2brPrUd9mzwT4gtSDAiG0w+VhLgMz+klPKYyXv3+5iwdF40CSkJ0B
fRmJUBis0YgMPRBiRr6m6iw1DbyEDVxmKx2eSz0cjnGdVbTEqaBxd9iFEhPL6Jtd
LjlHPXN3uxPRRlDluKY/JDxU4nU11G+1Lgnh8MYnFquHLZu6qoSLUzvHH8hnvVK4
tepioQTHLfBOJQ4MbEyQql80NV6c816ATvtRoeHRqfQE7E6BjHI5b9tOUpXjPQw3
seFyxb2hCzNRnHlKP+s2t13AglisVDEi7EdnDe3IBHk66txQQWA9HE2CU0ZTrMgf
X9xQ1wYE6UE4XTCd+ny6//0XAn0Wzc96RSgjW+3NAnUgNDwdxVOA8pxvbxWIOG9x
/1Q7+JKnCLTt6BRgeerpXCgn+evrFvGZ1zD2EPPo4SPtLEOMVNVPgMCsgfkFV6o9
N1NP9vXgtwKKbzsDxYo1gGFOyORZsSJ2xuU9zteDylrSLrwtrOwgjShibOaIWj/h
JOCqWOW8zTTOeMmSqhJyQUjRYWXnjMhfoUFdtQ5zGo9nYW7CyY90w6CrnwpHhTfe
pcNb3zMJAt3TuFe+NkHBmrNYNjoqlebMQOkHCRvtufNAgYebYD5viicWfo7NInSc
3/8ZC57DvNdNoIoVYsZqWFDPm6jL7UM7+zzilH0Jtgqm/TUm59HA1NDUWacIdQ07
k6mOWaB9k/RgENVqJPo9jufoDVXTZ3fnP4YHx177L1YsOfH9ywB41PyIm9GrIHBA
DTLq1tnOpKVANbBzndrSQZR0E7Bzky5dqXX1SS8edco2st87Sr/2qUJvBiI1pz1B
XZwxWV2u8BM1M1B3kaZ8wt+nEnQU3kN7uNtx7TNOlYjh9ZWhAwIWGFsuENyJAkuS
6g7E8VWov3yZPGS+JfpujEZC2DJ0RSd6VIeNLClP8hKyGCgQcQ//jzXoEDYqZfCk
BNSLuEotpfRildm0Jt/E/5AipOntfiFODsu7a2kPF3d1mGbteg86IJZHHJWQhVng
lcTRS8SveDhoAGY7BdzzRuHN+6M5kyY6GmfBPtRv/nFWx1W25WkUdCIJHhwRHS8X
QWacB3IkOyXh/GfyDDg/Rjeyv/RVj+gBBllLzMUgdIB+qeJx7YnVG7iLv8MBh+PZ
UUqWbdoNN/ek68GcMwKlLc8MHdtSOstKMVnUUj6iusmRcQ2w9+P0yuYwagXaz86R
8YOrdFSaLFua7JZbprhpJhBKMqz8GqKJzWxg6kbCPeLSKhwhNSd2nMdPadaKpryZ
bqZkI/L/4FJhTMHigrYHUDxwChfPwAR6bPLonvHE3vh1NeJ1YCuw/yoC76KwS57m
cwqJYLHufkHFnbeZbH9XM3aKbsBvgTBP49iP7SL1r2UBP1cVaV+9V+nyWjRcrP0l
M8vI+09F5B7tbmXJOMj8TiNxCzpMGg570qmiDvJr8xdTnjXubyyrsTgzcJ6hKV6z
4oPBikyz6F4NII7NRWb7GPlnwcQTKoO2QTauO3K9Gk86GIIAWxuhin60fPd/dfpG
Ryl/aNOUYIQsN7z09TPza2xCUTPsbuDFuQapScUqczXMychPE8Uk+J4d2Qp7d3B0
eCFnm3B2vxX8yOkYInu+ucwNk12eZ6Xs6Qre2eLYN0c175no3MT9JfNNupuhMa7+
Yb2xDN8VJjL4dIkbYfbEkwBkz0IkqTrcdbPOM21jZfNf0Ger6QG7aILcdziTlOMh
hNMkV/2QyDbEUXV7aRG1g45jVY6FdhjcrBYeyRZNE2mJRQz02YOyNMUUjmBzfCoq
jCJEtICOrLA4nipDxbmkC7ZJy6YfgMMb/gCTWj5rEezYPft2yhOo7KzcjBH/EgMw
4j4ZVgnS0UUve8rB/McBZ2xUNFG0DkoNmvmFgG58/ed2hvQwvJ46G0cg9W64mvCJ
u9zgxTTsuduMjbvf6/gvsBJXquMTddo2wIZ+y4j9MbhoE24Qv9Zu+lOCV03EOkkj
F7ADyt/vx+uZgnAnkfIfDJN+BHvaHRmGnBrixA3y73KZKkSQFWeWy3mX/kZHaFJj
VOFL9Xm3M1t1/QenBmP+Su3lRz8N0X3/fz5CVU2wJFp8SqOl3mVb5Eo+l+biQbf/
NPbpT7UI3nOp867x+ugPDhS2TodPZqP8Nc5e6wDmWcDmfwTE5nC9pvokrGl7ItCb
/Cac6+xNtpyVIAgLASxAAxN1dhVCwM3Ba029DanP8fU2XT6LYp5Jk+/u3ZMbyj4h
SCV/NRGlkDLskjac66ZSGcFd51xhwknMVGiKkJCVoCHjaujoa8akEWM60V4td9Kj
yyp27s+uj4lRcjI01LRAKOvqtfwAlAuB2d9NBgz2cCKfyQ2n2rYfrkmBmHHOwAmU
hq1kCaQVRqmGhV3W4Ns4Mp1QXISAjhCruTK2E7yxg8xS4Gxz/87MTREu9W+xoXha
YXXtKQXiniRag2QgwrbrdSaZo1B3YSRB1t2TbM6l7Ay0poGdXLdSdPf1d5lYdPhP
lyZrKTw8oZDxZDu5eoxibeCXtMLZzsRLeUXm1b+7+ibIKsEBVU7npedZggsHAiaK
9cCWOvxQYEE6h6qjPZxwTETxf/yjTJnS100i3DqybZ4HahIob6sw7XqPpFfwQd5B
SUuxfDh9m2N7GFUE9aT2Zwlwtt8rxR1Bx62VkUIrU8L27Cp6ZxzY3ay0/AZ/zgOA
tzETXPD0jZ0xyAJT+jbkAStIsIgd9B+97NI++BKCbspmWR9j2VMwbKdvQNfmVUwM
vWPMvQN7GzI+Qq62xY0/3l2eQKoJBLr1CPIclODjmgrtyO6w4m0YDE/WAfTbBcbs
/7mCLd4t+cgu+PUCkSMVuZHhwIbDenTIUHoXPf9eZ7SQjB1GE/slAw75gw/nBcs+
0Jpeq+KKLtDBdH83jTLVr3EJ2cFvP46KRGyZMW2G/r26KOkP1iDTIE8MZHtlV0br
1Dy3LvfQat/aKugzPP5FvnaFeSq/1hGHOykiP5ElM1P0CZvzTtBiQKJScsHSUJdF
YJ/vsVLG0vtppWBIPZbJVLA8s7XRfpHAeXhAwV9jVbJ4EwYTM3HFEhc/usSqxXXX
c08VwkZ9G3gFS0I+hag/8KqXhZftoAQv7mkKUEaYyKDZ6reoBHHwl8umGwSn+mPF
YZN51MW+MWxbLjQfeKqy1g3D8jvhUjtFn1IwK30tT4uqXqZ4hlqGewPZ9NCT+9Mt
jWKaWwHXr0MC7cJG3ltM3Phtx+DokCoPsWZl3OQ5f2rD5oy4EIz0opzpDVEQbkUx
EIIQGj5bmARQFyD/fLXc6JmEd5B8UbvL2xMEKQeyTCwJP+NuPaX+aJoQwmTl2PDm
6Q3YLpPAq0oG6zZiMV8gpzjNYbj2htwW9heyTsbvE6qydaKum1xfc79ofhbuYxqb
QQbO4Kl8dwgopzDouIw8u7VWNcCkegW/u7oMWmb0dT6j4CEvpO29TYc4uaFcNj2E
jRNOdrhHP/r+tG4nNer5v2wWBuPkvvY7n5vEotLNFOcpb2CkWS84QlzFWMkwf2vD
i3bzzREw6+NQw98ReOrcuLttAmb1fKcROdSDg9A+t2kUDOtyo3rX354iecTLUCRM
/vkoHoIT5+/2EEPWf33ixsWf4DY4QWhqrciht/ccspoO/F/HZgQilngdTJpa0xfx
/x8XvZH91Kcd41UeBR6kOWIf/Bt3/4Ta+FweGtEI1Wz9ZVjj73SoXVzoZR9Suwbk
g3dU1WiTax4gdP+CyK8wEJYiV/u9uU8eenfWLtba2pRQKy76E0BpFKuv3GuQE4aQ
kNeRnZ76AyQ7+RB09lAYyO6VWLt3KjWxLRWcm6POy6yIW+Cf1FwlLDTywprRNULq
ctLOWQiEqeBns/VRlWve8x5831HWChpQra+P7ydWORps3ibYgWG2uIzX8SgDvAs9
VBFtlYwOehESX+4v0XA2CBzihZnOTsQoGUhcKvOnjnpFses98raJ/qmiz/tiNyz7
8xkzk/WrnTmHuR4ETwLTESExgAzTxjSwKdUK2t85mEsKBrjgPx0NVX6/lYGKQCR9
40kf3u/t5TmEUqE/MbTBoKjU0hRrooagHpt7RURZewhTcWjFjvrKpodFwf3hLDKS
0ocbGKwClS3AtvvT4SERWzw7jr4cAYIxmipc37/6iLyQ23Of2+LPAhkkkEWqiGbN
ysiZ17Qf9w2n5O57YX8yXx2VlXg5lQFL0vV9ZxukMit1rfVugbVWdkF4rYQQGxuT
rR0hBthdWmdPli1wa9kpY5BpFXSWeute0zBhCWG1bvTTk+iy9077AUzyw+WhmwoE
pKvGKX0tIwOiY8M1BIQ5Y10+PE8zCdquPFJA/bWg1+9h1cTGfy/z32CjH9ldzzII
rGIp6gO4FSkkfWO4fgsh0l2/WDDKIi5chABc99Sj6Ct2u6/zGl9TRdQ5tuDKN5XU
gBv8KezYpvOnhE/6RUG1XilbVe1dKEfG+f+A9Ynjmmq3a3tW4uXxkcuk3KjPZnDG
n3lFpMqFr05s/auBpsCjtITTnB5dn7NL3tEXm8bm8jz6CbjPsuexUzPzNE3EU1it
XtPENw+iflEUBzdfBnfzK/Pesm/lkQIyrk1LDZ/huqKP1/GtgGSQxGDlFTaZ5yEn
w9eC88rsGr7gGrI25tyBTdJBLcL3tglMzIswcCN5CZtKPjxfi5iAtUsQQ0+sk44r
0AnJilgrCupPwK4y3BWZmKB/KSB9rX6F9hTKv3hIVESO8SHl82oEP6BLv9LP8Xvq
dgRrUn4It3aeOZNt1jsKtT8WsJmMxrPvzkPDWcs+kqVTMPNSguhvdoROm5QPDnlt
SS14EFCcBCgXaf7SopK0LGHre50iyO8L/yCxnbkKeBYIY603iQYXFuPP2b4Z8bpL
BUV+Hq4Dus5e+K++69qBnlWje33Q/FwWBX1mDsMnvzC+VDG7rzeXyg6R1Gvq+2MO
sGIZ9B8xtupox153Kik92G1hj6OQtttGg7hUxdRiopfyvbuFMyBDkJ8sfj67pepk
SG/VpvehNS4lXd6o7QInYzf4i5biTRNQIdd91CBtyKM7Hmv846P2y8DiAgXpgj9E
eKfjj1rtRlwHLqUn1AG3nvOgmI33OEpL05l863/uBdHuKV9KLYsOKL/ocn++7+bG
uwDY7QgfpTW2QZJ8vFVE4XPo3ecdEjwatts5/CXoJ68pyDMUYluz9kPAE/PuM4G3
NvUw+tfZPdRRPfYNl4jh0XUylqY17gsXqTOiihGaW2cySCwZKG9GXLRQBTg/xCtJ
hl5uvUAdO4CC2ACPA2uJcQfLQruglH3o3dEX9IvDiaO2F1D79pz3FdDsvPwFydwZ
D0LlURgvjUbyTmgot4WGy+ZR7Of5++EJxv7ufvog4qPbDuXzZsEhkyA+DnpjzFBw
QZDIimWf4wNhKnc9le4j090GiozmNoPf25FKnRNKdY06zQ8WuEJAbu6kej1TYpOF
hy55PeEhAKt1+WwGS4YYhFpcSuVw8R5hVnPohM78ECQVFhfgJnyxx1PXT65cF7V+
voUSL9is5jsVZVqWScqpP78+ivxNqrQeaJeZQH5w9quu/DusPI7XrYiYuQsarMeY
Ud+wJsADR1lK2/meEcOyAnbyOu2Hle3/3pBBTkgVEfHcsXJdEOxxw+QiWTHYt124
WJi6wb155w5F7Xt3r8PktkEjDYKGdpEpIXc4BuXRwgDzZD+s01D5RbRTOETD0kl1
zv6ZE1NB6SG5OmD7UN+ods7ROHG7RwbotFDmj9s0jfA6HeRhrAtDUWJ6QTVENphe
0h6VrOeNcLLhRsgZYbWj9XsTeb4ELrouXywZMBBQr/cOiABuBkH4dveq14l+B6YC
slJUb9RVzBS6c5QM8XVqP9lK7h8KtObNpBXgVkvyUxc2mw/XPmPuUPpB0AlDhUGD
XwXMHFVCaeEWgklABkV8kKYWVST0HeXNloG8dEoZxe8YVlrsMETW4P0AlFOS7IWV
VptPyZ+p6MxfILNKhTcblDoI6yyl8pd5DfJnslql+b0pvDK7ZTpawIaTjEA89SMS
SjkPBpuKfUSvLIynrEHZt4ne6Ubcbm91rwknrRNDmzY9DnT8drDoSeuClH9WoFMK
3lCAhOuKQOT7+7MLyHC5LK0TlBSWWXaZUqkpzXdECgzgtz8PBYFagpGb506v8Ii3
sE/XkhRwRUKGlqeeseaItD/bZSrN7Ru5H+dRC4HUPimKsvKOLLKcBdVLyOdU1ZOy
+hNtjoLHpsF2ekXjJ7S4Uvu8MDnQIF5y899WuYBmDBNWe3o2MdsX/wY7euErP1YH
tx6JvoO7EW/9/NCnxPQCy8q1CW8T6wfrV2thf40pC2PYurW+UJsVrJV9v62s1KO8
thVetlI5q5ZBn37avA0Vy5EtCGkt0wKey/SfpLyYU3dXDpPQ8Jl8pM0/MDSWen29
HdwZr54Nw65wLjPA04NFR8b3/ZATQIvD8fJuITtaiMQxJPeRS44kZ7121yk6eAr3
j3cHeqN7bLpLmKOknOdtWQYrPRpazhH2d6N7dYFp4zUHltSnepMjUzGMq+WrL42G
9waNETZTZ2L58WnFKqZFPaVHsd1w+7TusQgJ60DBPkwOdKgH+gQU92lmgft4gphi
H0cNM26IxWMlir819FVkb//q9wHqtDMN/RXBSghEB9cXAglmlE6dIPCCC60Y5MNF
cDNUphiED32+7atlT1vejCdfPDZAUOlphwUTZAf+uvES6RjKRwTuyOnLnSg/yD8J
MCuUh9qKtBsflgeVCAoAvdvgnm0QN2u7AfSoWnU7CRZHZv/U4+tp77SllE0H3P7f
MyOqBOHLpoP04DJb9t02oHE6jtXIwgS/os+V20vCHHd992a2PmKmT1z2vVRgC9VR
99yf00lFGOCMnRohAxE27RleM7O5Dqngw80WaJFDeB4htsXMa08Lx/LC57GKuU7s
bxRlFPE10l0wshBsiP2L3FN4nFLyEc9R9+CV993mvGNFBkmrF2t0VH+iu6Qivb8m
28F+UsdMyvjSSbi8lSOmdfKoUnd9VAZyiRbJMrYYB9mpxKJbZ7xxzjEcqjHhHDNh
TRRmMw8ogEER7Mn+NqlmnD5yVLULPHCieXS9hbwnKzxspP/tC1oddvLZw6OYjsvD
iE1rYjB4uWKgOsMIBZLA5cfM5UvclVh+g5ZRnqw803fY8rpJipY7wIhYpBFbStKk
/lkdLwP2TsD4MWaMvbWYBEZRFXFcw0fn3alEMeU5UibierPwZtgrABmIj4lGPY4X
3MyaqGHxJWbWlNNe0hZW9w20/oR4K//JoBScFK4p4g8XOJpz+yx/ACozqQOY67ig
2UvKv5RHy01A5pYAp58e5sFBOPBJ4VhQU28iR3XpNiTCDgpOXgVvMySKOG/12fuT
HlhOaYzEYAWes37Vn7ZaF7xuc7pCs0EtRMpoNQ6dNGj7ao61DPdbY66BV30XqrXD
TRI84jswT5cdflxJZJggdNjcqLJGEcoiKps964lKhy0er99ffz23q3xLmrIvEuU5
ZbsRSRkdCNT2+8enyYHSl63+xe5xJYw220RRdk7ulfF3o1RrW2y95EQ4FDVkZylT
a8tVTpze6vxtiWXYlLBfgpvp6jyitbFmw4yLuoXDOdM8MoOcSt6qQgpYT1b8Lq5S
aAtLr+dYaWSsfsYwXHQhYlp3XooeWOloq2ZwtIPnqa9cMCnp4GH3kOWhp3zIxpI0
byJXQE6xYeBoWuTTyyrgCb5xxm4JD+qPQhZLnFgY0Ad4etzoTogqyLyupt1isD1H
6Wmf485jID/4krnXHP6dOcWgEdfEdM3O1w9kH/yCNDSXmN2f+whUN+ez0OP3L29F
Cv+aPLLO4iUn/DKQhzawVBzhdWUmHkcPooQI3/rFraqBuP0ZmqImBBC8PjMhfnX1
/UuikwqBGn5Kzr5eYKwbUI+Y0UTOaI+qhzb5/V/0sri3twmwTI5BmLs/tTGWqUv2
vORYer5q4UC2btPlFLF3p8lw39HHZWt7gVt9tW7E5YKiTMSVOVRsf5mw0s9cKwqO
h4L/LunD6Re0yiiI7Ql0RY+Z3TBSc/Ye8ulnRZIbmGn5CbrjbhK3z+2LSQEZ77BM
IVeEw7rkzsUISL733BxMKiVRC2Edi2+ijFtQzm/GMxrPeMNv8itCuNZVO+r5jDZC
/zUNm/A+wwqN6mIXUYkn6sedFBFtk0cXjnYGknFiVJEv0FexsEoo1W7nDj8pM2Az
cmYWuRhqb9igUdqcTgrYmEPS4eTJrycXLnqPAtRAtj96444/w6juuz2pO4xplNLb
saMXCU8HDHahltaQIuyuCjax4BBMVvKYRZSy8uj3QVToSxRukW53IjTfzrml65Fe
GEIlIf+ioo8siTT/57RIM3DOvYV1ymGg494eLrRDkcfsx7Fesrm5x9F9BpF/jhqI
Hf+JFQ4cnnjEgD1vgKari2nDThc+LD5eYx2oejFF7uBKOpVFNr30GOy0OeVkvGIB
MDKcuY9YLu7yndXdriNt6qpciTeP5j8QxYY/85ZVRAVGyc7RLwKv8mC9tlXQ4CZ5
hTTsDCM0Dg/80xQoYF2+ZEcSq5fRnUZa2Pp+cq37GkSByxCNNcvv6vTD7FiwS0MP
NaGsgWKrNpLoYvWAGt+5pE77l9+zFJnkT5BIwbkTT8SLu5+InfoAeRRXFNgkqhqy
oXlD7RL/TKwC8fAoG3BOW634sbVDmLlvMgap4cm8NGOsNR2H8l0SgrVLjqlmLE/A
07F9fDZPmCQaqaISPZNuPdIJp0zTXn1FEhefzyyMR1MurHG2hbGrX5z1s4cE7zpY
HKj09xqpxSsYElAZFJ1MZ8PZco01VNw2kEiliImjShkzzVNLZoKKIOLUtw4Z6za1
CDv/Eb5gO66ePl+FvH5LqrfDDujFtaviSjmK/On0g++VuT2ufAweIYt5lagoMkO5
tQp73CKMR5gzfLi1uGRvWQIy6EK9TOWGwvL4OFDe86QTXay7ZkilgX9wQ4VuMtEI
xDWhRCwfSPgpL5biC2eDa4etFdiPGrz+reqA+VqAiEKYD9Y5hceTNrNpNraX9ffb
3bbjc7/Yj5vRqf1TM+KO176H4WrwmvtzrF6oY+UjoWmaHZql0f7uBt348GMMyy5r
r6nvwskDcaCKhChUQuKDM6MApYPjKWZrUwh6xRDmB5o3EKJYrO16T3g2ShB5+m7n
gj0oF2skYKQBwwAmj90i7ayPwRWVUnG7+MiAJLOCtf31QwxeltGCJeNeKDHbtvgx
iJc98f3GrRda7Rwi4MeqzT/hh/PQZC8zQjjxYaCj92zxElEO9CVccs1HfMHQXxs4
6NWHjmSfXp21keRxJ8knKioe9zAWX9QkN+eDAaUbmgEraCEYv9+45TXeHehNTcsS
ZEtuC83apejtgEn4s2KxucZiPLyhlD2g1nRqpX37TZYKj/T8raBh2pyICd3SrCOn
x7OtVJgjCFwHTrVet5tD0nwMXwIL5QpSwWxRIOzJT9RDmDYNHlGYVSP9GC2HK7t4
mLZAJhltC8rifv7aZJGjkDOyOrWJg1gKMUB7xoS+9M9B0LXdZgl2ImZ0W7bujGYs
TbExSU0hQdjb8evHJn8Q4NqZhPwaAnB2x4L3y80p7NQZJNwoQk6UF0/hgHLdDsr7
twvmK2o/jnt6gM4XzUwIo9LPzJC50pOm4M/2WnPHZkBd9CzsUE4qNRTDSqQ8gPaI
t7uw84Zfgn5Z1A94wKGUeyiHg2wE3fb77GaBhc4btfEVgyj7pSjGzk9lj1Iipfj1
Fl9xdsWmgf9hkImAm+5eIJ4JgRHxrW4pFEKsXOfplA9aK6ImUs70qAsOzwwy61GD
ByLW1pCwWZ9xMWDS+J/gb6qjhl/xtMDN9AFR3zLPZ4I3qNYOEyyuDMBcbUOOPnXP
WmhV4YasxCps76FsxvSp9tVspaE6hqxzdbm9yligcdzNw3HSDfarIWaYGICEFgXb
QAa8N2O5jxbGRcrMqe2eHTSu8YNaSKpKHbS9yY92FG/gHCl5mzT0F6OvAAvz0TgQ
HhYaGWKAsInUd7EBI9UodPOu3Xh2lIGl/6V2OUkkP7zm68xj+CIEESMqf9W2WgWS
DlX9o+mDSSXRJPPe0El5IW3JAHOIisoy8Ied8Ko3ctpFiZNNbdoMM1yNRvGDQq2y
ZMverz/tg3oQ33uNllBLPYYOP3fHC1IS1/Sjc4atQ9YaSu21i4poW/VP+mfKTurl
cdlU+gX4txBT/5Vmui9AeqxXFEksedM4xVYQ9yx0wZrcejYUTGchHD1NWSU9gBuo
p+tFOuK6eVTzQxGgFYNvupFQsH268FQWl0hmklGCe8xYkIOMBqILKy6l8tw5uAen
SjOurDmxXM9guZE2j7xwcNESbfr0x/7CTDb+waGg3PhTB2RH20N1dO9FtiU/Dqa0
xNEPWOFt470lshvUYIATEzYEAdArsgBl1MKMLKFUIP2tYLkD3Q2zQAEvhyXqo1Av
KKHyC1I6rjBZSc4Qm0Fji7oGnUAZZd7CR2t6SN0Mr2KsuLTCAxH0pyuVReDVUZA0
o6TJ1sJJCZemYwqmAOZV7g85191f9sw3zCMDkeLeXyG3x+OA3jocG6FVbcrs/prD
FB6FuSg6tQk96dUfM5aSAzdfY1yDHMWmaGgiUxOsURxC1hsF01KSWOY8h2F87Mnd
6hhv9xpDcimuE/Xw2ljTDO/JsYJxq0Y8hiL4f+uXqw+QFIk3qyXQmK+2eGybldqQ
H/yWTY/GzaQD6/yFh1eSGEPfoq5Uu3kvxgTlAtF48tm/AYNwreFC3I5FbO7S3Zf6
H34L3HdjhNTevx2MPMu/oxYTaHHpTMOkX2QXaDBI02cj46a3pIKVbMAaG/0BVGca
FxDJHU/rZpLVkihSFxTtAoQJc7lIASw9thg4LjO2qir9OXmwqSSdqtfa3jagnuhu
t7xx9vUE087oUoJyoZVWQFozs4BuJrEalmV1c45pOilbCEQlR3aKrIbmCgBk13ud
UIg+oKukSt5TRPzTf2qiNc8hz1ZbYdLlfplSelOB93kshWP6xhxJBtpJFGVBcRbv
BbMdcktMTGOUaYamqqvN/7NbFFGJP8ky2dyByzEBUNkiyR/kipqkKGQSyxAgFyiw
Fk/jiALTkqrkWqBLk0BvWWWRWqW6XTxVQBrumy4/u64pzjnyGMOx167hcOjtf44P
d+YxkG6YAkLdB3GHxKA6PxlMPwDagmvrTgUGgR/l93DO4lBU3ZaQjxIwC7Fkj3/S
4gTdTN1PNx/kdOBvUytLfcUVWNUaX5cEwhXd/OmjZV02DkJ3c9EEcDJvCC9kRV/z
Zm4ZP7IyjjpcK+gor/3Q3tsxVALiJwlUPMGNdoF/ISdZlulJBuWVmLTbRkTiMvgD
GMakoTieomfqSxDJQg4XR/tfzcjz5TILIPJwBxAV/POFR0zhc3OQPNrBgyhEIvnx
8+EjWNpfWjojzJmH/uMNbtwmfkcZwGseGRjG0/+RbM3DzpM7qssFSDwMUfh36gRK
xZ9Fn8WcKPmJBdT36g5KqRc78IrdX8HQme6yLBEzUBhzdz5alDolSvyN7BBTbwhF
3hc8w7BLMof/Q7BZPQFF3wioxPJUD/sLB98e+N25WhgytuWpegNLfeuG9ktiLhJc
fMDhP85ogvCIBcvwwh63Ue/co3rmgiG539niYXN24JVbfnTvY99eidayI5yXYBX0
BUImawMgtKC0s+L9UV0V7HnH9cTYP9nvoMG6Qf84xhJuqT6O/hnpmo5vdrBq7W4w
h65JaPglBX8OJyPo/1xh5AceYnpImpu77UoDfAjAMgRwFAZTWA+GyH+o5D2SrEgs
xYaNAAthJYLtD3rScip+G8Q3vNv3k61zLVUl+FqX6c9JeX9/1mUFAQhTSurEK+Fw
gYlDZDE+4riKzTAEsKHRzXjBV8OkAvP1LZ09PiFaQqA24IMBn822XA0n65Fpq886
lSYVXijWvch5wP9xFi/iB8XEqKp497UU25ESwzK/f7EQ7Z8pJ3JxEIzlftjrDuYL
23siYWWCdmTuRETH1r04Al9hZgpCyZnr1pyxqi2lj5hukhCgub69HTWn9/LQzicd
7a0OVtADLkYff1Rqsf6mCJpz2OnQxTROkNKbfnWimL6vp3OjDjwsA6mQRxEbW7/X
oHRB5Br37pnTKPBb7UbSzsAcV4/3rl0z40UTVqPL/AoFHZKqGw0rcDNRmmaoif6l
jye+11YzCSi5b5xLfz4QW4c/AQJdPhRRPgWvJbFVi6rmYyoHiGHUnoNxdBnOSJS9
DWsoKekqjZ7s4Lrcff92L45N874b9zwXa7kNLQV2DPkURUXaTCW9/NxFvIFwiPbI
XWWCesYZlWB7t7cK+8vENJBTENfuLsfpBhiZTWHl5SYFvgV0WfxFdsv3ID60wcIN
OxGJ7RtvDxgD4M3SurE1Nv7abHcIouhB/ZqxqjZ1P4+rYvmJQg5AOMHACBxFVfII
4BnoeaoQyQ7m0Oj4HEKmUtCWi1nDteh3DU7uhYyrf65DgkNScLLDChZ8kOklR05B
a34qtWFtHjlM86lIb5o0pUjU6yAzwNQHZP3pAgZNw4yPzFhgCwjklzFMewqCQHbg
7+PQaTEYzeGMrsqkYrmjQUkHd2quoOHN30qqaDOwXTTl+HJldjh33wwY9ZYYDUrO
VmuRxCYC6xMByw1PU5IpkUEc/vJYaumP0P3CnZJ/usTkCE8teSnQS0bd1ttUreaT
L73gUE9fzVL2CCmujVtVMKoCcU35YJxqP+/8q1npn5ASnvS7iZaeAvMhUJk09Pva
Q5h1aNWGud5bK3oF67Fe1GFvfejPEgy4/h3cEaGzgDab1qq6mq/7faNkUPpcpUNp
J8nvuRC+BSPB/KAUfTJsrEjvOWFaqqiCJ/emmC1EAWxMrFFHck9dISYHbiWyXz/m
bYe+e0/hADBoDslA+s8FOPKA6Ehw326GX4hMMkbuavSyAqWsLNjxFGXXPJmt3YBo
ATz71F/zcHLzU60rC+WHm8kY1lKPLRqFD3yBhR5V6YKCieZYCM2LazulrPRM9GQP
fF6Jj+oM4Gf66GGuut1OjBH8QtDrWk2yA4EOJE++pGi7CCoyJLwvrSaFcxCfknfK
rbpQprIc+XKdnswYQKabkr67lBu0S0gCN7w9Gj6yEE5H6/iJbfZdNq10VluTw/Xq
N0iWjz/UVM9v0WdG2ZfnjyOUjq/DHOwogcklIKbgoFxe5QPNW1Zfvx/xbaHMDzIh
rJ1r6utfYH+5s/6xAttAE2YXYjsU8gk4xdipUzwlLdHPv/qR3ims2BTj/obw2H15
CK6CLMYOinpdVem9ZM9YxmXEMlxgQtOO9l3U49dt92CbncHJ4bpXSFHhvqjFcGLe
+tBzuq0U4DBcBEWs0KqpY6NCt9ynnoohe8uQbp9/9lXbKdO59FUSdMcaxbYG3yxf
LBn9NSR1u7o+d6KVIJRtoQtQ+xFRjf1W9gBXjMHPtguRUTLahGpnuql6ri31+M7I
5N81S406dxUG0LZIJynfvwu2xlQw9oIUZOB3YclLxVhVEr1bt46dG3/s7P5dwLW6
QqtatvPfvwXuqDOAXsibISHwmnK8shty8qgZQv4Owg4upgj/WL+VKDr75S9SMBjA
J+TLZy6EWsEBW7nOHPTUnNP27u39l0dTvbt6PBCTeK7gpyPbLHSeOXj3qOCWsqpz
GaPel1pudm+2a2CnJJ8K4XczH6zaKDsrkj0KRGsVa0Ew8p95klJKeXVgFfOQ1cs8
7rkx2JKkv7rznylKwa5hjzUBQpP3it3lkDZf40admz++jn0EPCy/jC3H7behdQTk
7nfo1N0TwztkjG8R013Ti2f+ISy0ZH+jYHc9qsKlM4LwxuYCA7RqWQJVbKqcWLCR
mFnbbsH5odOIQf4MD/AYj0VkUNStWicvpG89lr5DIyHVu+v5MpPeP4ZvOIpLT6ds
zPnJ7sfRQmBJ0bGDYTC6HmBBn92fcRup4rP76vmdWEvAHZ4tIa1a8C9kppQhKbe7
JCO38qCIw/cANzEwOCdYUtTqW8hJHo0WwHL12hqQu8EZgZqOacukU/70hJX5h/EV
KTaYPyUrlUlNzUXZ/hyF2ZkZlK4m5Lnh2LCuFNOVD8SAY7h0VqELzp96561CMxF6
qnoY/3bd18VglbfF8oa2KXglo+pwLmXd+YHz0vV81RvVGoZhrRtJLMJFm+VObqZs
hyjNdKefMahGHr1qkGwpREyQ/e3FZHvzU808/1FVF86T8EcEHqILMhy1Udu06mK2
cUnMCMShUIB8ZiU/KNI4NLO3o7R9xL0RG0UgSLnCcvE7yaq3Fbxw7hxDTIiDJSx6
EV8gU/6xA82THcCPolhWb8du2YGem6Rtm39mTj39DCA7D5Y3Zj4NFXZOHQIRLhQs
rhFmAAh8gPJ9Suym2/hrseE4NDiNOmnrVvN7IlLdldHUK5X3CLQwgI+Viplz2a9l
3uoAzYfWAWn+jvYgbysnQC2UWSAR3xnvGlB6QFLZ5Z1qEKNl5dNgCE80cUcQztje
MZTNPmQK8dxF/mFdFbUxxw0rppaa0pP+gURh/xnxvKASEli1Y2Z6fqmc6l2kc9gA
ztUjSUdRGMxUDZ/j4hYXvbmD1XpGpoN3OpGyG2BFpTLbvIBgsVpm/cQhR1flvlhi
MrJ3q4TBa8A7lt+wGg5KqgIiga5yoLCYfAtZtOLr1XeVBMo9y+C5ZPs+ndRc7an5
GYf+VH534ZE+lrhAa/mC+vQW2WDwuSruuJtX76AconfPdFgdmiNb5NEypAjXNnTc
4nFnh+0eYy8qZfFGVyUMgSL/cdXxHurPc5yPMo7LN7m1Zs3WNF9U2FuPhXgy8e+s
n46Fy11xCNKCYMa9305RpH7HsLcHXxE0P2O5iILOoxc9Fsfz94cdCHS/PdjNYVrR
Xy5wpdCD0IGlGmggtf74fKDCREARpu1EF7+0hOiKqmpuPlelI9vr7zbudnQsIGzp
eFcuzg1J0Psu0jgwSNKiN6xoOtY2oGRwaq8mTkjObMMHqWuqoLzGgjC3yDKOhn0C
kFhQjnn1JE3fsHkGaBGvwUPWGojY00PFPP8vlI2nmKJuqj2tA3QFo8wh4Jm8yKsD
vcP+1FQQrBWHWin2wuTVn9V/oEZm1qSYCjZ14ecZM+Xky7Pow8Kc8wdWa0yCOxFH
jkHuHZbrkpIojP61KkGzYaLXSxbuRlFuXFdo1VUEbjklAg/YUuoc7C7PW3du3NfC
RPq4W/lHslNRbkOWpTDOicZZoJv3LFzC65a18V6EVwPtqcPJTOHG3r9NiL1FfPF8
/He/piS9cTRMyDZL2u4GwzhjEXvx/hkBANvCo1yaaCG74DcYsXEIKAVivEP93n1+
EaSFdTWccIB9xZAvcp46c7rkkAyKbKfr1Nh6N3mHqkda8x6LCwrXhOzc8B6tq76B
WETyTCPw7R4TrY7/w4XzV+8LOlknx2x4voKDdM3qhg0c8/rVGCG5baTZwC1Vcf6n
BjULBRJDOFUBK2nUeYfVYlpyMeSOUqLA030X1Xw1vHXdIBCR8R3CE0JfDdGtybUv
oZQ06wxKiAcIVrUobZOjS/0St1EcqiUqdTFXZmmdB/9vWiDldCY+c8lIWvxz6hsL
tYD2pKUBE3+WkJE3CC+xYGEnW/k630YVscnw4WT6OMyeeQj8+tct24gNrTUEXVsg
3QZj7OfcO1Rh1Ab+TVeCDNBc4S8DRoBGq3k3znG5rmOj7Rmd/XHFlozjTOz1tVtN
ydp1Z6ex4l1mkhiVgXQqfGASqk2MO5hqxcRJL2b/6SUFoevbRS2EqB4qHVhlL3bc
n+e9pTAVb0hniVwryXX0+bcsA3Iu1sT2VYnhPJefLGqbRnlDInGquReh5cfTtTkC
Ewszv9wGbJqDZryau8+sbm61tiBfdqtCstgiAIraOh5vpZ+vcAK/MocaTkKBQNmG
rOzgSAuLkTp2D4G+U3JtyuBdhrJoOvEIFobS9vC+2kvRzlGoHyG4b1ERUfEahWdy
Rm1JqiQ5lldHUCZDlVl3ai/PglgHoLds6BFJqsGXT7GEyuByC+5alV0ujOPTOKJo
uc7zntEiLU0bmS5CxljcM061wROHuyxeo5knqU7cFVIL1OH3e7MEnC/AesM0GXUp
ajnhx5aJluyc2s7y9P3Iq8M/Lq40mO1Htpc83UwIJ86uQ9Ybk3zdHMFT/JWEO4KQ
2vRmh2iGRIA6LupTSqsqdxLf1ZQuQvVjI2x89XmHcgKsvS0y+7477deaB3dW7O+M
XM3E+7sFuEXKv6CMMm7ttpVNYM/pLu1vbDoCCkRkdGwFvw1G5jfa3brtIlTu/mLM
rldSzLCoazO1XVcZJyOnKswO+KBCVCcsW0rdyal4UaaaXLsXI9c9w5rMlnyogvI3
ceCdhSelkmFKdiF8h85KRzw0RvKObIMNFrXOnv6dx4ZwDqgpzwAfiZFdYj2qWnBN
rUArOzi4Fc1Fo6+K2Ay1R1ICms/iI0sZiUt8VgHqpcnAVbeBnL62nBFXWMrgOMyX
8Y0dYJOBIKM3QwhSNixPBoreS2osaXF0E4Vj8p9Uz7cuu716UnarnGhUGRfO7/oU
indKkLpPBd2GHd8ql+T7nLFB05xpE1rl+OD92j1xeP9iP1XLcfgz+7CrPjHpFUG4
GPcaUbsfQNTuuUA2RJY4wTLhJnu3DotmXHf/wpTcR5DgtCpgMhxvc1pE/n9yan7Q
q6S6Th7w07+Vzt/6To5TmcRDIMr74zT6Om+y9yVTDhrLVLc/iv0B9EZ76zsmLETB
JNod92NSU74EZ4C5/QZFVg93/KLuAt0XWpQKXkGXxgxqsqga17CtqbC2Lu3g5I27
qh3wJgdza/R9cVoiKouyPZR6kYndrX+doYpwCuHLOPdU3a7ZeOLXqY9jt3oLS/ka
2un4TtypuD8u1gR6jAg5a7JOPohf/2wmfFzeUzm51Zfcep43U3RtLWBAxRde1gub
imjI7gac/XouTXbXtzFSr09xFi0/D/cbuVTD0m6M5tpfPJL9Ra4j7Vj3xsdj0Mkf
OQN8BVmwmV4p8D3m0NPYT+oOLXgSEGB0F4UQOguy1pOe1YUZV3BvjiAatYcc4DuO
yXbUWmCKh7uZTrCIoKR/naBJzaboD0eSivswArJkGK62sZh6SaYOvDdQM8TArunk
+bV5f9/hj2nFCVuYyCQX8manbbzwf80maVXDLDn9yLbhFv91rRGdjtZP6ctIHS/3
2M+4Sybho9ePmByhGAcTJcGfT4Ncl1BOYkgLOQA86sfBMdl8To/DIiX6g9cvlhFn
iurmdvAN1Vrzd0J/X+sn51E0j+Fkw6Vou+CkYHptat6E+A+CVczF5SYZFDfeEWAO
cK9dJxBkysd3iUbw5A81FLjh2ExOCZX2W4IttoSml6k1M52/AerLLIrLCUE4bQF2
bm5vNgZl+cK+Przmd84jKjjfZD4sCZjG3a4yd/SqafW6Lew7j/BteYpPvPtLS9H9
F1ipi2/ewOPzsbG/OKRviL5XZu/6cPrsI/3q/gI8LJbQxyIO2coeakSOcSGG/Y0o
Rfem2xgtNOP4BR46u+qJzoJNNFoaCei9Ee+zYSwjyBj+5nwiihyFVpGgUzodhrZ2
78jjxU8NZn7SzWTMBPCzWLFe8KM/hLafU+Sc3PpHZxHx1XTd97+/YfN0cWhfQ2NN
rQwmZ9ywacjVPZrnuVZg1l79QdFF/v0b/Rd/M4MjePKb40Q/DvxNGzd+ZmZ25g2Q
USFcaChoIUV4G3j+0eQuio+wSdt2mqxxS+JrOXodjBjoBeEl0q9XwU7l0gsurCll
et/MOUIILOPJoJmd4bls5fP3EqWHMKGJk9VTUKkqk/b50oLP1FEE2CTvogA9D8HK
BKseF2fO/6x+sYBC8bWE6NKCybif6kLFicfjPci5IEkdfxA9TEaq/5PJTvkUkJKL
ywkuoXoUks05xR9FTYrxOPhR6qyMNL+x4enUOiZ2aKQN4Ap48JG/HRmZkusz8dSj
gtCHeQnrhRdmIv3QWDKXJ869Bvc0bYd5LoFKa0AGCkVzTciARkW6quoQW+hhxYvU
SmfQbwZiHaY9wXFvTYP07ZNmqtgUpVh4H42JymfZyWwl1zZ5aaUUAQz3WiIAgtW2
dzzopfp+Ry/JjnPgEJz7W2++KxOyZiDIPS5Q809IA7BTKyoX8l7GKb3YvzR+QaEU
56ThmMxEdCkC/rvZtQJNLqQprrG6fvx75/agrC54nYEBNUr/WD7KfG5M1U5VbBGs
meMCPvzVdWxvBPJ+GaV9IykyWiSAcT5Kf7BAsdBcU6psBkglBsZ7kNssbTopVcrq
T698SCYCInmUXOXSw6tCIa+h8HrqkiJ5+j/Uu8bS0hrUCJ6G1E62UffJB2fkDQSD
gw2mRB31R1If6wzjKd0hqUKZYOVogpwIL9KxcI1weEbGcvW4PvG+jNLDa1XWytEq
4hCYQarEhjm+D5P9f/7xlzpe0qoznMfQ9Z+tVsAJ//w0H9qI7Ra2dpleBRgXfMDY
PpvP05VkJpxGma9y0D0UALPz1llyeVhEWgjDlGJ05VPj4b6hshfAxPoJK01PkBvQ
N3rchrL0amQxEwbzBE6Tl7N2OgNTmDMCykT1+r3g+GidhNoK2AgRy0Pjh0M0K90P
LSSPiCqpDKTfDONBYNo1nRHLVVycJ8dL+/MD6Wthu2WYTWxOOWdh2Sx0vw4npRq3
7F0eFg6g+OGt2tg+OPE2joocd6j1dafcESaPXqnjyEJdZps2p4o/y61QAMvJBnPI
SJHIYKfQXaJyh8uOmqrMLFsrNdPp33hoUo2Ry41lpyrM0DbZ8kDhdPQkTuCCMjo8
u+H4m5dEQ4WXY/ZcnAyDHgjlv74OESTI+TA52OrI8mNr9Bl+lFtbVnw6OpPcNzQf
Km7aJ3qykaOHc+p2fgO8kIwxpRoEKMqlst7yE2jFmgkoI+Gn6bXXV5WP48SD4o9E
NgKqFHSvI6+rCmRL20pC7IUYGSzv+I4JTepE0mA/uFGP9j8YpYzjhnoRy/DDpler
6TDCKw8fj8v7fxDBx6y2A4vrcDceHt5nsA7BAy2nbLsCSb8wrFDVGJYgcwXNQBB1
5S+5TgDtGpdJ/pQM5ymM1xxMIcWkHMb8A2L8T4Vi4qC2fhydZawcaaJykw8gklZw
8HCwe0QexAKC7/JxiL3EbTAr/Wf4FXOMnrxsz3wq5MISv7YsoQvcP2ZFDtjAGQ6R
KVbcNGGibl9vYS/lZqpOtyAx4a4pow64wuKFMv6VGzu2g55VKeGtzMKaCtizDY7Y
thOvx8a6E8ySrPMk4uLRaJ0vB4nOZYgzAxYsWZwKfpSOliIbVM1I4XoIoK4i26ZC
u38Hahf0x+bkISzzHhr+Pv2tX8QktAKlN7vqr2OVGMXZbvkZipw8jiPeFecjW2BB
a2rmq90JRM+AiNeVEj//F9JLuEfvNpm0ghiPM/dG0aJVfBDIQ4zkqdKXbkmfLa7P
Mvmc53YDEDh8E0QQJChfhALJh5cihnSZYktlU3iCcIcjQr1D9FA5mQmzNtsql9nq
fvXgx5bOhpDSwMGhBxHM1vc5KAD+8QzH/KtU1+6vo2OG5ud3b2X8kSm9exoSU2oy
8RM8KDHoRyu40hDhIhtijkn4e1nDA10r5qm19Oq5SAchNZL+c4OOV2VL31LvIxqP
bMJQOYm12dwPugu4WF5lUtxMCrICMvkEdb3DXFkSrfxZf/vqi2GG+CMiQL1SKYEo
jNOqSjVpgEhtxNiw2PnwllzgEWrF66QuMJRhs3aCUCgCVpMhzxpxi//8R+r8oJOV
7KrzMghLkKZpYT1HXIFVtR2QUfe0BBxkMG6vpcGv/c97XNRqXUwjXtvEttiUAhPh
8QRQKz/oQcyUU3zl6hYkh38ebpBda7cPcFR9sNpmWBJV74H8tcio6pCbp4PrnMVA
l+yFxD9KxUMh+3VDmSgoad+kerWyTzAeDADHGHDedM27w3oB4A5IDE1gKCLUp8gr
hmT0kDp9cI2kT9W1LeSe+bKif9fKU58jIPiexSDEH2eyXsfzemp8kFiOaN4BV9iC
wxsKVilRRSPbfCyUquQmILkiEvLh7/wD1ulKOV31Me0LUxk6y8GTj13AmS8SJDtf
UNQ/pQ0qSGLNWyXxtT3cWkR7AIpWWpi2aHYElVg1eSZsUtXVghSpW1VqXWYhU+Fu
gbF+OBKDwoUv7h4ZBGy7CpGM+N0IgvM3zo40L/CWl/P62PQwjDVlbZEoguQM7eof
SQFbxpSk39sRc0xiOwbT4Z0xPfcBaTRBhdZs2EgsfMMGdP7RHLBIkwMrTFxZoQ9E
Xmeb5wHbPeQhQatWUWah6kQx9EIq9HCwucGCLkbbK0Ue7ZTUSUdyhZZN6RwZlPQ7
wAZE+aC9f9U4PavjOUDYih5GJmGtM44xibKdpVgykP3p1KY0PSbwDakx+3mAl1E1
wbAyAzyOIX9IsUnIkpuZJxLDYjYL27XRKHiX1PzGS9oPcTwBz72MiA8ATwwxRPfw
dkXL2yQMyh9EXh8hCpW4g5Yib3T5n5NLG/TwA5GK2YMMbnfwmQBwB6nY65xkNdgb
XVE5wMqjoj/yWCn8vtCVLelHTuMvsFlQ84oZXuvcxQ1gXQuXkLwQJJeuXEbv7rdD
Bs3np5jMYXA/DBqM0zakbjCF5omE0kB1xREzq8AHog/4RDxoKGGp7ID4qt8aVG8+
+e0sTZm2qFAmbHGYTC2GugAiVnkdg2DuPJs+mgMqIzS6tsJPHsjjwRGOlqDZ6YBU
h6+ns24eZtyidFKqYGz9/nb7WwGgPCo/sMqMYfpuvdMopQs4JrmW3fSy5Rh9aNaK
7mf/PCVAtlZoLPtv3KcBPCm+ear8A4zbUXku+yC6fmvcR9yfvnC/GSI/skwW1NqA
jY7NUL3hb9Dc2J25Oz6QYDIbtC7axotg8Ohv18UOYS7dEWPgRbEqnxZQl5owwMcO
BkLRntpyGAEfHE46odHyoSVP/A4P6oPMh63bv2KHLfWwcEFbHgtGNNhhTK5tGu1K
FJ1l3MixT8hgfYVK21k4IgRYvNv/0ib0S5ucjiSd5wUSlpKqKXGGomhegd7JU4OE
9mVdPXvq4w8FMVRzqFGw/Mi3mwsPGbhMa98Hj1tce5P1Uuvb1SSDEYqW9RXonqUM
LAH80rAfRQ0W50SqSd7wEN46ujQMk07Pv74BtyO1a/4UB53gSN9ljm9Fc2ApS9bP
HThjs0oq/h6CRcFU/XxuYOkXAGlrXXyat60mvF8xsPSJV0u2wsI6sFOqzy0Q45/A
jFoIjW4T1Rx/UN1L35wxNmyup1tR+41fkD8ZZxWxUsXC0awZHvL5VpuGdDX65r7+
NpdiTABWMGpWMRcjRqc3sdq2FleDpPXpbhrwfyJfC8bG6ofntPIy7QPx/wG/QXLv
p8m84VdliAKntj72X0h26nDMMkYQzMf+MIDMUex9R4L3TAUZat7vX/gRH2HiOeap
N3zwN97N1sQd4xFh23uz1IZAObYGuaSJANSib8ButacZ0oyOCnLWOg+p8NRXC0/L
50LZRipoSJQ9p/NU7v7bjJRjiUnj5b3E2UaaEtRtmmbq8m2gaSgzNILGsJ2LMiv9
p2fPpn9Nh2rktB4FfuFZKYGGWVCCgDQnHqJL4AxjV3eVVDt+jw8nfUVexmwrB2yn
7X3/ZIHnViJoXvXNfd4m/FgIi4c2i+WWg5f4QL+F1Ot4WefKndHhQO0m7LGiI0TW
D9ZxowgZ1NQa0jcN5TIMLTuyxFeB+Na9Wpo4/2cfkbIh3m05LZT28yA/3M996t6X
Vn7lWfPviqrZW7IfZSs4AEoKNTL+MNLA9nYXHaiiuDqULPAo5krrAHKs1j6fwaMz
lJweQ1jaocMtuVkyvKytP5thlsqsMhyDn7OhQKOLHInauOe8kRsFfntxMosrnN9S
IAVfLlidb86hobzaxAMsoKQnhHPWkmzUSvZRUZr1KBG5jNkf95LOMkSI7zMnYOYO
wsb3N6eynfjNdDFSZwr5KIfd0D6Q2/CkytHpUUrBo3WFyeJns3SHOIQ5hEaCclqO
+KxyeDhXV4HF/N5sYtzZ68Y3Zdx/4drJ/5YXQ/PhWNMvAttuS2tmRH+VHo+LvgBh
9e3XFrHt50PoAHzlyTY9NmHc6S+vjkaX+NAKM/54zRBCGtYHMYkRTpmj/sWnN6u1
oiaY9CVYYzLuI9AW0x+5M48i1dipIxI8oE9Ff28kYd7YrEvHGDJAqL56PVw91fOi
M02SBjzPIGqhDM9DOiX3sXreYgt7UD+eMuG/TRiffpntm96/b5MuefRe1NqJzIG0
zRdFbvyxzknRtPRpVncnZQp+BZbdGvYoIt6MlSfmUSrC+8JS8n56tcHq6CH6rqA2
Z6x9IOPN7a90zvNK74zDoaiu01rXhog3BdLeLxCLzoF4bfU8GQ9ne+rvZFZG7dva
UGA3tfMM3DMZDQiUm8JtxU7rG9dppIHDeK5mj+jMyD4OrZZZWCjNY4pl7hho02On
NQuiFeJroJC87IIoWLbsn48AFnPTC12ieOr9KUvgY5UyhrmCutp0GLWPlpOKYD2W
/iTg4HHjfCyw81V8ffeFksupf0AWZXVB+w/3uIv+QDItk1lsfYdSjvLaXLGDCqHS
RXBgsyiUENPkqU72/0sEjWYscGk4+pmcls+d0xzglZWABN7meT4gNzscPJqoReFO
f2p8NKzygOYk7PpokZS6oYJ5tNllfkFiQcL/o723qEUifNj1q0Kzez3qNna+dNuA
19iYxLFmVELJ7hpICDkh7/UW4vH1LzmG6Fv6O6N8qz7eqoCcdVN4sZJZUGS3HbhW
TbdLAb666/bTm6RAXPY/NCxn9oCXHT1t6wvbdFYfXBpaqgCPwP72H76vVxNZm+GR
VVy3WZ77d1aahKfTfAlIaz7uq79HYzGSYXNisUctYR+iJmFholQ1oly3cgjjxUba
4YIwyZSk+Gz53xm6BL8uGVOV5cGy18kFJpJXzwEFcbPbFJDKRaiZNt8LQIolqXA9
1LA5+QxfbjO4hke3iF9EYt4l1qKkpldXZUITNPNFSPw6uPgCQI7sZcqLjwhJSrXK
ahmlFz7NQUjzXFKZcwDDMFkpnGi7CO/hTtsAASySuie2Tmsli7PWbQaXWW3AXzJ4
AEa05oPOx/+fDTIiY0u28dNU1zonmUcFqlmIzRrhHrzt7Ty2HTs9GT+qXQhXP9eE
10C5dOzExBmV7ThYtTSVnBeoqYLDLPwzStx9hmAZ6exc26rxk544kCQa0qiB6VX0
wKzvsYa/wGYQ2dwlVPZ1Q8WcINKYJZ+9dy0sI2hQEwAlBrJlLFvIW9gGARDBF/ji
vyNir4AT6x59jBL9UBp+8aOMItTbFF7UHSoNVKCQlhLtdh5ErXInoZmRANcIErkX
0uZvfzt9EwI3kROy+agul9UTsN0ZdmDVUSi1lYxJKDjXRQY6zkR/6VPQxlOcYwmr
ow8al0SDFtnjgs6+ZtDrDUPNZmMIEUiauKRfwGxN5i4sLy3XDtQ98PdVIh34q2sM
s3vAVezvVZELYhfjgztRfBtbRzDqxhEslJWIqPsbq+KiOC/sKLTIjRDKlvz+JxNq
T/KV0fD/keZUQxI9padg1HNohOxSmaDMQY/SY1yDilKe6GOIVdnpOCYQ6eSyd/e6
zMHIQ2JpMWG77Kis0VmW553urhFcV9TGrV/AtJM5Clg21JFqqpwTRBhNrpViqlBW
ATEuU+NvNhSRfY7Ttd0EuA==
`pragma protect end_protected
