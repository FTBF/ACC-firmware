// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:40 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IDDrtn6BqhvdzdHcrcTErLaRzXe4Ev+WQOHzgeVRkFrQIYuvIyhFf2YUbmIhcbIY
7tfYP6tTTSVP6qFGa7JEuReaq0eo9qAgpvPZm1G+hzC/Wq5dzczA+z0GHAybMQtX
YpKJEaf/4iJUHHcEoOHko4FvVRXFs3liChjN+HWDWtc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11312)
oLkVRNuSilLZUFeu2uJbO9ECzvCvytmaoGGPVjsoEyLF3/bM2Vq3oNgJcL7BvkQY
ojbS5WUDHxttuO67zqsVwjXpYK69r71Oyc/CJu8U6pVSZGRQDr6doljXKRNRJpq9
+L9CLsZA3pV/cId8nZVOx2QtwB16Z6F90PDweIODr3LYJptyvZ/PrmzLPv6pTy8o
vsNWjFW8wpIk8MuTiWOzH9/hNuFLTk6X70YYpuVTGqXOI3d7UJeTbvniQjrXa5FV
KeMhEXkZ3CmWk3V2t+WtgPw4J7ZfqgVnhzDGITCNWOV2qH+6p2JQvOrziy6yMCmc
7lTDSbcBHQv3h+G2aaY0Gc+hMkSDN0er3HgxwNOd4/yKfxiNTAT82JZseo3XBHHk
PAx+XO+8Llx6rnDQ0/08/YQG/xBQcsWFvHHvqoP1SosREPBgSlGMzSvBzPOr3ZKS
+49qSKv1NLEALgUSEpYR0zFmYdVunxVr9Pq+2NVHyxMJBKgzlZ+69S8lUS2SXnin
SyzysNdL+nLNqVsMwqlBpuIzdT217uSG2Y+1QH6PwrMlfQHN8ZBxJWERHCOwgW6J
lz4WmNF0QEloF2lsly61hlj/b/jtkkKAmAGtM1qPtAgBwyuTOw/9KRHyjxKKQS1X
IKeWzoysmAmm2sI04Aq4WGkDAkWHXGdbhEnRuhmsndC/+6mx9j7NW/DpOcEYbnA9
mPGZqK++NFDdQ41kaMWkQdSVZzxgalL50xY63dS8/Md45/YRisu09TUaXcna7k0Q
8JPi05RAK5nE8JuA5DlhzfaVH6KZSU8pl69TJFe1igrgZwG0zaqeCRrvqX1W0rms
idGhFVSbeAss5nmUqdWjVTE+IjUWzT5o8jOx8OP9Wwyd901sPwZc0T1adJMy1Pfa
IytM6LHUqft1SA5ZplgDSJKH5+BEDB69W0DW1zdCTn0UMWGzy6yggESmua7ZgZBq
hSXl0LTj6fYAQSM8K7i14XqPt6YhTG+WCntV+l0O9AuxCwKnG4nzBac+bfLLyzXo
qja6A3FdbKzKlQXcrxDib1VGNQXT2AHnw3vPfLHb7ZHRwa8QNtDs+igfKnf/afzt
D46owmUMwN6WQgr/nzzZ3VF8QHxppI7Mpcpf9YoYAvOpr1TNCb+8nG2zj0B2kXG8
ofy+CNMxaDxzvaAqkxmSCpH4Zc8q9wGbCU499t3gznWrYY1eBm9RmPQxvG3v4nNQ
iK5YHNmOjgJLnH3++vVkEwGV42dSkrPPn1klXMD+1qUHxwJFHv6N0WOeYE0490bR
xaI89OFNgtSVSQdYaYH7cl53wAHza50bU01uVHON8Wmb3jhUxPDGtvoIhA6LA1Xu
2slcpTAgZgfr5Xhre8muEWZpUXEt2IaQFvkocs3DBSSdiSrxbW3lul+6cbeqJEK/
0Y81gHfO1KgbU5YuXV6Cz+I10cgQNcccRFs4sPL8Cg7Y9+QIp7DU6xDo5IRwdLjQ
s7QZyQK5Nt9qt3nWC98B5/Lh+sifrUl6U0gWSQwgmgOU9B2FdZs+RY+K+kwdOaBt
plcjvqN6JmgYj9ShNQHWgE2M2jYlr0XZoyuz8dCunm4ZLMCj5VfB6fa2XhMEDvfC
uZlCMpm1gj7/CVy6UkMjrSMCHJCbq+D16RQOB/lpYWFEjCiRWUSoTs2dPW181iUx
CoCgNA6Yo1t88mdRtSSxZz3jkAC7HO5ENgKgIPZYSm7Vug0z5SIf54SyKfeHaV/R
Yfg+Fdn6gux2LlypAuzL2Ib3hAnhBxTbYazgIWky+/ddRX0ktB1YgdktExLURrj+
DFSkQ+FfdoQFwTYV7WWC+ezMV60eklqN5YKK3DlWCQKtppC3TYa1D8IkNzrv74rd
ZYipK2qH3D80GqIcVFjN1lnYNymBcJuGDiy6MhN4VAqHN6n/srLMNqSIXk0oSVya
k9HzMMWc1Tx2uvEB0CsAOyho3DTITL0xBVHh2h9dr2FVCZwHRj3VlYi7ZsFGo9iO
MWvZvbzQwxPhfq8WfkGPnStmme1fdE94/+kdkKvRfBa/ezSzxCK6bmGgXLgFwbp3
NiTSqVSFwu8UNMl7mrRby3DeYBWyXsVi2hxiTFRKG4cZvtOS54MplRJwbsVOaaRc
GuPWyAtGmKUEYZoWTKaQIjW1jC8cdQW356y2Kcuzf+Zg8pgjEQSUfsygSp0uYC17
7W3KtgMLvY2bjAKo23PLnsc8oWbrSEKlFdz392XK6QyOT1r823XaQsPKNAFtQofa
2J1osDTjRKLwwqKoZnEw561gggpjZWn22s36GMZozZRroqO2dcW1BfgRkCjoipQG
ytVMpw/f0pFuud57rjgpyccOqYRjWQSdJF72UQ3+yl8RP76+e20b/C5j+23LoWHE
67JRhnr53wXbif6oHjQp+WSbzkHQ5CZbKYSvKlWXCKtvfpNN9I0Rr9c+gpaydfZp
2TTWdVsKTpK1jXaRFb53ieFogp6vXWsvHgeoSk7C9bo6GJ+QM6Oklt0WCcoKmHCL
qa7GipPrJJvPVT/AEisUdtIWfL9V+srCxJ2/v2iaysKPM5ZaCbcq3tZIOBJkFvd7
TsN8qAZfW8SXhqB7VVumU9EfWkMPNRPWXjuf+xZwN86Aki73cY5LwCDGn5qfUdP6
H3j5IVazV0We1bV7jdstqsTZ6sL2vn1YzlGu9Fl+PrRbbcl9jMx33qqoFxUjlmdq
BGaKJzy0HujpeqDMk4YoLgzf5T3VYw9ftC/AAyac2W+mTFjXQQVv0jKNaMHiezzW
zEzOtB/9/VCRGcukqDAjbfjoQRFLXCnaTRF2YreK5okUMfBGksZ0IfVwHN0GNJch
mWMxliUVi0TAzJ0uAE28qrvrf2vehnROIAT7hJ6XIpQKrf4ha4Iy66b7e/MLW3ax
bMUrP3L/08cbonaiIBsd0/jWYeJ42W52JcKpam1SpT7MPx1NbMhrLjInCAs6ouwt
aocadGuVnvoa3PNOFIt1PtdOXRysQJLHqXvzR69bcA+CJEHekHChQMsDI6FNJ6CD
4vR8WFpXBPKn7mF8hE+4d3ZSMRnKAB23kyWVvbH8NPVUYRfMNMkFIskBa1434DKM
GCI0hcwB4Q7eUon3j+yUzls7z/0C5wdaCnyrl7t7u0yoABFYF2L0zegeEoJLHqJO
CKcc+6vAiGcMyRwLtpPHCd5UyQZNYWNcC6EDIKwNisEqhzC6u2Tl0UcaEKu47FIL
Vve5p16ATWoQzQ2sA9p6suF0gRPtUFqDjMQUd6MZ1MUc7NfK+tVZXNdZEpr4kp84
TWP1czVKRc0OkjOV9Buaq6bf1/D1gfxfLWY+vn9Cdmz+mdJ8om756g0vf+eq6wIx
O3wwDaqXm0gcIxzRqpra9XcYumbmNZ2y8HxQv6kWYRXmG4s5VP9+ZmAQNZyNF8uu
ncN+HwZOgZhsTxMsDaNzsqgysiv3uOTcaGiRmdruvSHRBNqH2xTNtiSQIyClI5Gc
nvBpWtoJYA6ywY/tJGIhaxQD9GzP/VrHZfoZ5VZxzSE0TbvuBeFwQP3naB9gHxM4
5AGDLlk1sugbHbr/QAk5lm4fFNO20NOqx3aOlTx2DeMwDK4dXBX7iZMnEPGQWFsa
UVS9dc+nuxoNzOrDhokGuiGhKRgvz/RXZcfgvM9XdS3Qq5cAuSKxCKmkALr/N/Pe
pGi01R8DIFGoU4meb9O9QBLTYeSkAZ0r3PvQNB33+V9tCHBZikkgJy3cv5l5UOm+
/Wf3zZdiM9bPcfA/YPA0b25xodkrcyPG8OZe4IraCNnnBY/ZD99H25Yd0Q/4XYsD
k495Cs5jfRPe2IU3CQuOZ6CjZiEVfXPMgz36vOiv55A4DU6F5UFYfGHgjDgYnFMf
IsBlae6f6Rsqhjp0XE9xou5kV7Kx2dY3cjADh6kNPr4w7Qlp8qFNc6QI1jUywZGO
HJFLp2JP07BF7avtsZWeSIgJRggeBsWg2sqEhJbuCmja9UmG/gROqwNBKcag9pX/
6vC67rXrcB+coGVwsrs0RxsMNJkM6ZZbZXUaKLoEipS1H3wwDF5nxXw4zAeY6CFs
EyTqW8nsrMirUqhnkCUlbNpmJvjtRuXZU89z4JeWbGB9ct+bE/esT/UOmptrRULM
1Lo1eMt1UvZ1EmnJ1JT+s4Ocv3rmWmoydhJ2PA5gjriYL8vLfZyljRvLcqdRVDij
0+KOnf/WcbRIc5HqEqPDyBAwI/nqFZyv5a19L/UyRDh8FQwvoOU81Zp7h/nWm6Rr
w/F3iIWz4eBVGP5hYVahi0Lh74DLzF2j5/bUabJ3/m5SIhfsAerdk7wuTOKYDKYB
9va8LHOuqtMQ2SQ+JBucGLwRYsa2jQbUpp9863cBXrVZbgR/9nb4gkn0UwtGv/lr
OMBa4j2sXoo3GKsUaj/YnLctdoFux7f4n4ThwKYKjsnlplEWyLCBMg6gLqowM+q+
uesnDQxiQmhKWkuv1y1WlomOIJIhhqQfcyjULGVyw+CkqAgEnma+rvhc604dOZUT
ZttD7ufdReWrU63LLkj/2CgqEXUNBrTfVyPZ8/5/Stok6c0Dz159Ra3DA3W1xHOG
DX2h7iGDHpGEuCSCHyZ8SSnMYpgx0daOURFHt6zZsrfMrTAst2DY9rxiHn0zlZaf
rFRUU1FT8Jxrln7oZav6FVOIk3b66au1mO+Zm4qqfjlR40VvwZKQ+jWEUlI1fkQW
pCeKHhh2m+62BSkEVky9Klsg7aRuRm+4xi+wzQ6GspB+CEUJ1ISaN/iDCI4ge3MI
wfjQk0jQgBhGLKbsZhTbiLPzKEfKm32MMSDtNspWd1T2x+DtCjZ7ztL9p4+5TDj9
86Dp+pMjUOtVUu5pBdjhADAbOYHr75KXvkmnvO+bvHPP6iy5k+cjNA2dkgLBbZWC
6EBneT0LMcwmjc+ygRwcH0UbE+19B3iWsr5X5OUVxdCQMl8fhYekPi32+u0N5b8I
y0LNL7xLTfb9MwPZvto6uaUQc7Q24L3guRF/0EDJXjHthcPFmpPTPuKvBVwbPxvt
sq7kja5ttufL5g6zEkNYrxLPZK5cDv6hu1jb7nuHIdrXpbBgV5XcAGllsHFZp7VT
EI9ageYQoT5ALsjRncgK6bKYkDeKN/D7lrCt0lvMRKQWNr5R63bg5PP2uiOBxTdh
QN1uAN+EdxL1ojoccaCUAHyI7vv4Dxi5exazZgUvYOrw/U4Pz0wkl+m017Qgi9CM
YMEE5PXImyPzD2ZJFev3Vb+gFAPtLIAMAF6KjDMLwOHIwbTCZCixh+wBQNPvp5X9
eaqryOPRYUgt3kCOp0CtRphgRCODJJjcEc+qKzsyLKGChxe5xBrQpWuGTAFddflN
cD7PWGRu24jU2qweYG+1Z3CEnbm61sz93z6BtVUIjS7M/AiZACRL/5fx4Y5X6ssn
/iJHa5LAgz/1E0ZNkZx0MhkYwyPlv1jyN2q8jIscVIxX33DbHyL/FIaQvVisSDNa
p7rRvHWh0oFLK7FH9diPcLHgmNwYHMlRYw2FLuVqijl9senK2Npo0sPLd2vhFxif
gTsN0dpcVG7vJrrJLTLNMyA/wl4uqK/BRl8yzL0X2ewxvPxfNzE6GfH6GFX9RkfV
WAwnTOKGF5Jrg4uWpjMx8ha6+N56RVXkoughEoV+DC57zs9YIYWRM8+MlPLMBacn
lZkv0Xpq73PtwtcOrfBQRdEJorhO1rqG1wZaQCeS4XkPbi8bMywzMr/wnLiFJTgl
nsBRWGRjFFmAjuZr4OBilqIqT1GdsQoYa2YOlxIZDdlJnRa3XPdcWEafrSwtnTfB
oLrp6RoQiMC/chZFWSE3+ug63X5W57c87BNccSJ3D52l7b7Zwn63Pi9CJ9DOBYu8
JKbqA1FGQtgf7jOj8423O01A9yc/jR5fFqeXAmgr6B2uBzKmBG8tXYlOBDCyvfyu
xRbtUzPKtoVyUy1Q1ku/GBC0mXqcovZhR5djBteQ05fCj275Sy0m0k59xYLAwfW+
mWNAeQDGRWe1Qtfot6WmpjpOzag2/fkZyBF2nXz6sfoAq/k/1CLsLaCVVWkW39Gu
n42FSPfDsKsgGIQdtcbahYJ4KQI4o6tW4svLFDJgoiYA9IrB8INc3Rmf5+F9/jD/
qe01+rIbIyVYvfknQn5xrYOnqEIi+Gzw8944XGrumGpR8piySFvtldfoXYlQESih
L5pTWUZyTYgQB01/gyShRCbfIYxmIuz/ihjN8TaDCilKFJs9RKTErY1mkOkvTk1I
q9RWO7bNj/L+f4bn0PQ+mtJcIPvI8kIOFFu3lpumQgqOSqXytACAbOdkhXwF0doN
XjXHaMJjC4f0r4r8sYgvTCNlKyhQ+uTI98LlxzbaoXvOGmhTXGYc+fdh6L51muMl
P1jlQEre59S63lR8NLnmS8nLYOj6EH6jgmMb4gAAD/RBzUkd//ynPjVYSzA/8kQV
+5qQGuERZAcHXnNwStp65eRKag5BU+3ZU4PIg+RvgT029SdWBxbflyCTFUQHMNUQ
fZX9gHS9M2l+b5E2/coaut75DdDhitSaPhHV+92Rf73A96sSSBHFXIBmcT1fMUAJ
YdMp9e3xR8SaAgirF1K7lAm1rleJf2gduuFP8nic0YotnpM6zropdptgJWq1Sxjg
oucKNE5LQzUbBkIsIokuMgZsw/frnCd6sK82/RTjXtRI74AJkSH/am+F5/ueiP35
YAEPnVGmd3SE9FaEuWPmGWzx5i1MV+9ISvsLH1K6+x5Zq9FVySpjkwYAhgc7OqEf
IuEL3NMcSnTjW3zMXAcVOMIVVL5OXHtPyl8XWzwF/UuGVZ5XpuBXifq/tMmorfVA
dSsj8dPxsHheZL7iwPn9Ioxg+axtUreqy2rp6/eI5NmOz75nvi0ZjXM+kcvxR2Ec
urX4uMPoVTcgj6BpsjXl8m70DClzctKIJZkqtRXrsjOHoG4yBIQHspQsVO68hy1s
bkShmlUzB18XPmCGhT3/OaHk0ZWzvQ23iTQJl4uiR8EOyX4AcRm+B/cT0QbxYPc9
JZv0E80R1PDxymlPcg0Dicue0Bc46JuPHAx2u+v89rJwi4Y2kooSa5Xr8rDg2oKf
shhS72b86IU+q0MtJFwhHivW6vFEcgVh6xZIkAtvsWRPCy07d8ZzYlRIu3I9b4wu
7U+oj1dd2Hvswf6wgHO8aglm16nDFacGrFWBPp7f0kWrkoyk/xppOcb7NuMjS3O5
xkjxOuds52CLsFB8UAQukxHy1MH5VWzC7QoPGyEbGs8ope4fwb32Jse+kmO/ifLK
u4ynrH3f5b8tFRjpMPfmQrGD655fLcHRey0wQL9DCmabXOj0O93efbHc9Xj/R5/u
agna5PEkfGWSxOXwR+GtXdMZdcUm/T+avgE3r0mCoJX0z5sJrrcS3vt6zvdWGYqV
3+PnN1Ongf2sGNSX5RgU6WXrmqhhX+h+CxwoaQnBaeuJxNSIMOrKKl9k0QPQXD98
E7ZbBRzyrHxtZ1jOEVpFwP56L+RZryOqZJLjOva+dTZvwhZkG/S3xwE/BO8nN0Ux
KH1ArApPDegJiHAy/5ST1xaFRC/2y1mQghlaeF2BQQJoeQI7zazOEwpM/jD+FhLM
R2BwrXNvTJIx06I8WsmwJTnn/1drSdvWyeQ/lvvR/Jz3JsqBeJaken+7Rp0TnHNf
wLWlPb+muZ+V5/+fZILvt2FAu8oSezuqZNK+wD0WRU26PEmysBROPhmls8ubdJ3r
aWqcKlLG3aE3wtmvGteAhfvuL1SJ3D01UM2BfC7Jx694rYsOTfvoxCoD2QPB7b5D
K+ATb63smUX8C4OX02Nv3od+Y2ifCxybF0kBf8wzuXbABehi6RWpjmscnIzTn1gP
KHXgihmvVGyCMHYl2VPAmeCMB2oM7+OsByFpPYCfyV1YHkMJuyoaqr3ggimqz6Z0
sA30bhH52KjFSfyweehyHJRbsNwE6QUA88VCKrbH8su/V6l5NAxDAmqMpwBJadT/
x7IlpAxn2yzi7df8llfD784HqUXS/zyeTj20GLrGGBYsPUeiR7TLtW1fVdvAHD/m
Xis2XDIUDtdIyAViZhPQNhUnLMbYWpcMXpSltC+r0dzTv6fyH8LBdjzmM1K/Yqnf
XARHNrDX2xPKBSd1PDIElkph3uxaWeZeSfoDPOBQlmBrBktwSeJQa+TDs/kjydlY
6HPvzUlhkpDI+xkvEiZXj2mMCSYo/AIeDMs4gjhVixagFF9EmJQVz3MZ9AVaCvH6
KLlY96776I25QTXst4j6ZYqHAKjMKNycIy7ZHic3+2d9j7N+3/4FCkKNW5o3mje2
98YQlgiqRQAOn07MFuTsvoeYL3l+TPccJFFo55hlTfuWs8TO6Zz3BDTPA5hSe/Fi
RCvzrPYUH+F0joN0FbooWVM0WQQkdCo745mALp7eQkcmx9AWuPqK2VNEOf/qTS09
A0cZ2tGgvmWoP3vvGu1BKHnJg2IHkcGrmLDpm+6Hb0PvpjddRtblr2jmCnuuU4Ae
FNAqm+/NKcvxO8RfnuMHxAtgsEf+85SF5KwxpaHv1DBuk6txn16BZrm0Y72gjE5g
xgZttWr2+0hLd9Um9KF0i8OsrtQ4cpxfF+tATo8xeaxBKgJsYTcRP+hW1Uwo7Fkt
0Xsbu9MH9x4kiayXOfpaA8ck8UuFQkPaSKz2WECKnz5W9brjNW2rsEq8Ncpu8cIq
ntCUKoEn39Lt+qTDAa4GHMKgOPeWHP4k9UE13K4ZXXU+0t48tcOHX71ZcuQWdUR9
dv9cpKCio+a2/3vBEbfRCH4otopLEsCxtT5hIjpQElK6sQQ8Qm4/xUIOpL5xSySN
0tYSD2kz5FAWtmkEM/PkVWUf2PTtPK7lYgq9zaikEW4TqnPtKRP/Bc/6KN1yABkq
k5EI1bVu3irDIpgZ34fjA3N1awbLhLIuGcKi3mzrWc0IQJfBWQ5QoIxL2+IqCfW8
y2Jlm6Dg1Kt129N2FWpqyDzf9JRL4eaFyZdHjFKHId9SXRPLJG6UAa15mOb/HEzJ
hzEpluojhA+pf8vFuCcwLPQd/OBbz4uyM64Ze0BZJT3j4DP+RENRg3uCV1GLfhCw
9bkeSpibb3vO2GyFLmKklsLe050ZmZxLHkJAFnqevpqQPz0Z1p2fVMgVlw0uRk8v
bU1ptqHu7uBnAKNdu87kYrL5fHOGEXBWtf4/phK3v0Y4V8qKAhKKGPRtnZt49uhG
DTztlCvpIELwWUKXuD3q+6h/3IyJBpyZvKb7FxgRtM8QmoSrkNyzV0wCLvDDGXYT
m54v+Z/1QvUm4kAVCTexjjAkETDm91xEG86zjsUzgWKD3UguMeAp7HuMXO31DDPa
3H1l5Q9nslIxO5VH+8I3BGzSkY3Kf5hxXEzD/uq+5o9REMOzt3G7aoFdVhXfow9r
1Ad4mKEAHux1z9Hm5t4ey0ACZntxs4aXCcAKgLRaz/tIiDo9WVSK/U8VsLt6n2g7
lYZawu/1gEbUU0rsj1bh0pnjZHK7Jzjw1wiF3EM6STKDgR/ndN7toeUBmZ8SbZ1b
b1Yc5mkwi7ZDGLZHu0Luyz74DVQEK4KIrACRbiTdXEmXLuperOR80Wk+BTfncX+b
J/Av1Rxk8kfDwdKyXAINSQBKj5Xh1YwTHxZmGPRfMWSNUzZNcRzHIMfeS9nOE6vH
QGydglHxU2Az3DCI1ugbyrtBA6FbpNWuvRLMzCCENNYs4Yay0j2cVGN7auiOaLt/
bybP4LMn6y1wwUxOEmMR8dPGbRl5JnIbatlhifBV3qcQhC3EiXxJXN33mL+Zm99c
MegQIaalqzQrmSzw+EdW56m3Z1w6Adz5KRPJGcWFfJ53jZbP7uvx6i9VlxMGRLQd
GyZyohZVsb5hoKgWQ22m2H7eU6dgJAQCgttiXdUPi7uOA0uybW3SDVg4bOOWdnjV
k8w6Sy1X9Y2j66NJ9C4wkUB+BWex16TIPSZlrGvpyiOMySl7cMO4+P6p+W8IEkwh
F5KxNGAnZJAt/10mZUZzkcjkTq+jQU++Dtp41zRw7NoDMrChpK2t9pnhsOsknQya
HyQzgFtz+NN5YCA29vFRHpDwlOt5lLBHjU8HF/EmYN2sjh1qLG1LGenepOVh1SXg
ngOE8SeJrpIDLvBsWBbWCWFEVTEOoYevnnLyYaNcUvikviU7kCqqrOUwppYtGjmY
M7PjIKAZKwE7G5vQEeKQ/7n4fDZESd+D1nLXGOoPXcLU71ya5wgvFi1tnXEF/V6f
rm/dACS2zoYAe2LfPFknwyvPu8kVcQaDRA5a52CrTfNYAMn/6fy/373aihbPxHhc
Zsph8A5oLbdHBwqGJKfpoVrg12MK8HCDAdRaYWUtWnaxBKwclGMBLUzKlhpX11ix
CxWw+jjyeAAbGGOnRExUiJHIIzwDGI3ob1E3JKRHJYQYt2ToDmOp/Yvb0BefGpK0
HIfYjC+1EBejKuRGxsJYr4RADH29DsUQtaScff6m4DmuBZeBJCnjdYithy3pvcx+
9PNmKJzHjtfqAr4sBHZ+lMZbv0kRSOILTxn4ILjUDIfiqSm+JwcQQHRp+ZzKmBX5
kyrEs2s93PzrOoB2xUu4iszEVdXPIq5NHwZxHaoawY4eTZvPgNmKhltCVXrD6vgF
71pwSaGFPRPsqhGwxiQeAThhYKkvt4mF6WcmRId0e2jadwzefaVzDjWeIOC94ecF
5mmt9bKQvrXHjuc4ffBza1za4a0PSeEKieC4tN2KG5Ojhvj2Q5GquDmtBEGtLm+5
Y2GhhKQ7hITVjTxlq555WYQUv8fh7ZBgIIHxptruIPu9Afe2kJFvNk+i934ElFw4
4JMOW+o6Yu3Gphd7Frc0b5eb3D+PWEzTALouPNJ2zqrMLwzN7MSbirBevgxf6yUu
r1tYEebNfVEu6hW/0Wl4Iuk88iQaoHaS6PjwMkujD25BRnN4hX0CFE0BxbgSATCq
81XwHi0JNBTFAsuLxCcX8s5icCRJz6lsUJy2FUQKJwCyxdCZVLbvdl4rqTgKfBG/
j8yqba5I3TowHMnqtOm3mKcrrUdwvcRB+2HGAD8D/6pjJyWEWIpZvTtF8jIXk/oj
On37nQIggoGVyAaLmjqiayANLC1N89wAdlAiIIKw3K6WY6uwcgAMNoeR9a0+sFYb
pu5Ja0G+zakVMxXcIrZveLyTVYD67f7Pkw5xnAjuf/uOHanXSteysplSt5tRWY+R
c+KOg8fMxrlrYObj96rqNHUrrTP3vTQpsKnw2zB8VCGODvtkhvliQwYXRjBybgWS
j6U4aNiZwZf2jk1mllDfnx/YAhCCD26odVTJx1QPxi6ZkZc9un3AXc3Jg399ix8P
TERKwHykBoz1miJHr+Orv0AvTSoYMbuDBFRUptJPLDKpCVolcaZWTy56uu1AXOJd
WJtqrHwTaJqOLSwQtKLEbCN5ZD7xK71v7KcsVRH/o//xTNoFCRzM7AUzMWzOcNqe
xiokEaK5bSlg9aJEy1SvBUVQ5Uzz7v59Q5vnxPl5VAe9ZI0beqxTba/l6ly2mnrs
iTjWRGRsy6A9604MIobLXsbwEAIR+1WSGcgcKyHjs29suM6obRUiukHaI1p1rvtQ
KtJSZ9HtZR59WGWJgYxWwAmX0r1nKNC64wXx8YIU2IXU/pqmMAYb7AUcmf+ZgYSq
FvQWRk8DKr+aQ0L3FagomWUHDO6yblJ/+S5Ma01OBItXtCheAu9+1rNeAwaNNRKN
JjNhWK57CAYIgWhZ2SU6/OtrlvSOWVc+dLc/gLqqlV+I9BaCaZDfJKlZCejNRXSc
o5LmuznQ/CmuviI/uv+FDpcI9eKkY65f+hPdw1yU48BEHHI1oZTv3S4QCl81hNdd
XPV3JCWUjTB+EF+Ffsp2sBxUu5g7MMrq7v+tr2uuyJaKhYV/MErckX2bc/Nec5Dn
J/1rDMaEQKsCRKJNGV33VurF9WxycVqUlefcXbu33qH4OX8ZmIeXK77APV1jfWBJ
C6lryVhgn4z/ry4ECPxkgCSQdcOQuZKQ6o/0k+BXSg0Q2YXOnYJn7LqNXiAu4WwJ
lvonY1Uf0Ei8dznG/KBnBGcPCyj5irGWkx9DtOTNEiqWj3V/QW7b0HAQXwAGDD+I
8IsNDb1lCI7OBt99kxB6EmsbijxbSn3C2WPqZLw0Q2A13jGnrptteGNnJsYyU1Da
ju88ZuM7CNdn/uMIYgTQH89wBKZlo7V3B7nE0jdVOZNvkBVBUcuWAIfVyrDeFCAM
knsFGnkeHyejzO5MsPXr0m7VsIEjUzOECmudWnMtDjhn6bXG0Jy8H9v2AcbjoNnq
RkFFI2bZeIx0vRQU7qtgXveKLg/jvIAAfFA6/520bmAKbL6/McWDrNgX1Nc47MlB
xMCF9E43kh49DLWqWDFdeo+dKohT/o8tH5GBnh2NPfO+BQ25umC+T198HjIQXJLT
yam+mpo0W4LdeTfmE6OfnqslcBgs370Q03/ocUDTr1Bs4ueTTF+8eDRttE4+c7Hu
+jOL0PHEVIdBYY6ayVXhMelcNeg4+aC+P86QaJLXBnUBCAOH6qleq7Hfu973buk0
t/Pogp4UzOFmJi75OzCIMkoD0jv2irZq32T8U2u3RcRM1ijv3WmI6wD9iXPl5VVT
lcPISMMyBNPHTcGvRNUyPreHm83oF84WUM+MU67l5vpeHI71Ib+0CZMYxE9NVy/U
LT1R4LNt3/CXwZJuXT4PHKgVcyVdYSWknmTKXBPGNAgg5WyuaWCMTIKl/paYsKvd
OKXs++jgZpl0kEl/6uvqBuBUZkGE89byUBuRo0N4GsdQWvENnnPFfsj6gWfnF3kO
b8ay+i0d58aeD7ZgioHnPIZaGnp3VbFPd/2V+wduPblmPcDn2faUAvTNhQsHfBWc
EemgJ5Jf6tAOfR8XqKfLonS3QB9NsA2tXMXvU6MgF7qXIRPZ+Vxwz7VNoLM57LV1
no1ZKxk7IpqDsSDzgDcRHQxaaL5bRqnq1gMCXiLFOJyn+YYoz8BVowp3JRXg2KZm
q03psTx3v98a8Jej8ML+POzoRlopj2KUKH6DRA3C0/0GPzwijhWskH44nr6D6Zv8
eOGR1fVK8PWhzDZYuFRAJGkI9GO2IMI3tr+Xk9U+ciaKXdlh+d3QZaFTNneXSZ6K
Jy+EAXL8JV7QhbVqmGHrA/X4nDS+aafmhRian0ZhO3SxWWS+S66HGgFW4CO3mV4z
cdHfJhJEcmywqEO03dzWgX25MI5GGK1ba3sljEWl74Cmu58rpDnTMddbA5NTsvAc
7PRu5jESEO2FjckGZr2UVrFB9SAXzF0nYMlbHCfHkEXeLnQJCH+oDiKJFXhz891h
51yC3mjj+M0MhZYIwYD6Gx7sAcDSr/sz8aZGrLllqKnzPHRUJm61AkmHb7JTVrwN
qzMcxBg0TcxbGHaQBZnPBFIXID/DJsd3mgsxgrbx6U7+0kl3DyjxF4Yqs6mDlLVC
WGkOTfPSqM/MJ4wQ+YqFgv+vDQHdihexP0bYPRK2MU2/u9Ekvc/o6lxii9GiilEV
AKRe9MOBH7y98Ou7h5HZEMXnV1vKsTXECFJo1l7WDmG9HAeCsDv+qwasr5URYprM
Xab+nljhSZoa7D1zJ4nDxq5QUF+ilQ9D1+gOdWMYR3qqS6kVL+ZOMwg+1U4plzfX
/16K3PC4BJT9CT0r5SxCB36jGZokhMbR5HUFey45qwiv0nJ8R5LiN0lPBc4TxYFc
4eINUGJvf9YBBCibr9IjxJxL2w8rYzK7lUb8V7UeXc7XoTc0g94tqvo38K4mZE1I
eKRz72kghtXtDljeGpxMetz0HrLQwId3XYycAeVwb1lZtPyu2bJ4J07QKLjIpenw
dxf3ePyZnt9mdQay6mRfz0ECF0em0mWSKJnqwZ5y8kc/KyM9sR3mPamP8PMZGfGI
psEDlu95MqVpoHUY8DBo4r9yavuuQN1QEtbtot4iHt/TPbnAGoYB1oJSmcFbsiPp
UGSRjTImR/h3fxqGZBZMfAxVIK4lB3LiVlduAnL9p3zR5Rthhy+RcrySKyebVRwT
TxYVmEbVJ8w77hJeQ0z5V7cWiOk08G/Nr5bqJmXa/o35e8by0wBLUwWFPKbHtdst
YAoODOiK+uy0YygaTz8B7eFo5k3fB1nCI9/AxZQP0sAh0+bpmJbQjPrD/LzzaXzM
pACkoFSih/ZMYt1OoZ429z8rO71uhjcRQRI61tdPsXu2lx+kIxJ4GG/gVDvyckpn
dNwFbWBA68d3ohZsO5HvByGGxIRBTAREMcl11usmR7lWJ8+bcG/WqNrmfW4uml71
ya16hgZgGUF1utKOYTKp8oj+dbL/R/xvyu4RKtQxIsVxvkfNiLgthfOh9VlA/O37
ZtBi6i76vnBnTW5sYtzbSAU7wFn8f/2z43tQYNS+mYNSJkJpj3n5Z9eXtAfLjuN3
jZx25DemWPn1eK++uX8wMSAAb/oJhtMUwIqZFZF2m2vnTlORMoG5rjpSuKuBzVF8
Y4xOkWdkhCxb76yG0qz+azD8QVhPjGkSZVOoetm+uggh75k7jCt1BChVLz/ko1n1
GeG4aZxqjk8weS9LIA26kCd1pZGednntioiZcWd0leK02LEIJ5JLRnQaB+cFWvlI
rmwlIjtv1ZMvyyHPe+mlmOHylSuPhZKJT1tuttdwvrR2rqIYplSHzHNcZr9VY76B
/GVtF60M5IoE+tGLJr40LSnwBnIIDcsQJ5p11ivRVRlmd8YJm6cKyHoKovrKlaFp
5si0e1fPTqiZafwKnbRSLuHMWp5Br9TaOdoo48fSO21eDmqzZb45aIVMoaAS3jTb
5eM8MD+l0v0xgaxiHQdrwfyR4QIA3eMJTnwSx85OMsxo0dAAsMU99LHBcp7ymv3M
QePChDgl0dRAkZUG2j0ED2nIHOPzwv7XLqWXEDEnUvCxU0e637nr/zy8kYHYlCa/
733wLAEiAlIw4GZg31iwMUWoO7jgP5yfxZcSRq8iKw1JlLkYtq/h+4CujB4iB2yh
vModc4fl+aZggQGTbVxNwxtY01BbXrOVNy75rT2a/EQLcahtXN35wIHgkfPk3+fM
Wi3Q6KfTdbnNwAFU0RW1jNDi3z6MfEUoRi4C1WHjrQwg/gEiJ3ZX1ZDXOwW+PnjK
Rx75hrLJ/u5UjX+wFvERfdelprsaz9i6m19xGBqQQik=
`pragma protect end_protected
