// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 03:56:44 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rzqrYCQfsedDRB3MCc++7zsxTPUuNHgiXb74wK+351obHzzi8H+4Hzk/zbZHzmsX
TyDWGATwvVwxj+wRbu0Nqt/UQ33fHV8/s1dpvJyQ5WQiz+hUQV+7pclcna2AppAo
TmL7NdkYQqF//vYS2fuL2HYNlVQ0oSDpKEm4zlnxH0k=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18352)
Rt3ZU2nBTYy2MZHjsvFVR6IIIsbSxw/X8/m0VpIroB2G7NvIlf50Is1i8Jj8UmiJ
pWFHgY01GCgl+N3zG+LEAmWNypagnW2P7enVZxl6b3B+oIOcO4WFulSK3jRQKak2
X8K0fcdWRJ8z3ssOhqoB4skd8EoiVwhCRCcHBSZqpjG7kKGX2812KVpOW3N5KvHh
su684C/sH57uaD7hjvnTXbRW4xLftYH5SFXSSxpjqdIi0QO8OcV3czbmoN21hmfA
CIv/cWKYGJmyoSW1AUQHw16+JatK8GwgZcuvN9CMPdBnAXuT9a0pGc8oCkNF2dgz
2PJB7cOe9ilAq3jhfXMRvd7nvNtQOG4yIEW0J4ThD1sLhmUFBhzSSEQmjn5bikJJ
8+hp/TlGQGLbMfcetmvwm+lIL6zxb2UJCOZshVOqTwoiv+votVssc0E0a6xiI3Qu
aErM013UcN1L3YaMZ3AF8MSB1NWRQKZr4bXRIEXe+l2dNUUU9UM1ob8ZceMIytqB
oQY66V2auK6IeOg7W/ltyGmREDstvNhHNdeaZ/bWDOQi/BlXOoB+/aRHCusvTJX6
RQdjOfAsuokllWlj/VTVkkhgrGQhPfZ+Mp8lzdIUXfJqtsczztTi/a17MwUigsad
7V7KdY7m9IhpLzvB+okh/k2y5msg9htVHIV5LxiCfuzxjdYUYo9AVIZleX1lfC1/
yy4WzCN0n7H0ePKSm57mP7IDdBykYUzA9XJbOr/MbWUeDpxDrMdVjTgZExMZvmC9
UUnKCmCpoczSjB+419Nj0S9wgUqgakHqwQr7mEU/3DVyySiicuAHqTpSqvoQMZWZ
eF06zD486Phc8l4YsfqDMzQiBTKBRT/XFO2Rl9kYExbqrAAurGvgY7mYCp5RQF+B
J9FG8+IjptKT7zPGsuhJFsa6324SgHvYxmO+hl19V8zKgGmErYQpxhEdJwNHqYNM
h8UJgBTkoFGgUeJvmUXvyOHBreodONCVD65PAi5H7CglCpwkS5HVSGDCDHXjow1d
lzQx4Pjd3V3wPZ/bil97q//r+9Icq90PdRQ+fJGxKgPbe0fHxNNpFWmaruD4qqZ8
kNkyz1b33rdDv87ERcFBegcSzR9+CY8j+sSKhsQptbHtOiWPiMR+97UBZLa9noIf
t2+3C7D8baaWUG2kxT57wywlKXScPh1UFAFOhrY7eE1/+EyCfL0vgwKgofmQIOs4
6ycxkFkA+vBAj3D+0FfVqZGm59tsP0I/ZbvkeY1D8CVQRpTS8KSPiK3ildBBXLtB
JrSFJ099OZVGTYykal5K7gWV3l4KRi3U53ZFeN6WBlhJ642G1fZHcpP56v5UCd6u
5pZJ1BWA8Kdbp8OrUb5nup/Zc98rAhKmqCnlGRZPnoyI/epR6BdMY3+uhV4wNvdb
8A6eDBy4BEi2IvZnZvjhV/sIQO/2JsBCR6ZataFVln5RzVQ76hLlU5iFkaJImy+f
C6GBr5fMQt9lw1XeyFRcPRScEqHXTAJwr8+xAQBSf6RnyFk85NB7XeHrqftGLG1s
Pgg9IP/5HccGyfIb1D3HULBbMY9XN0Duf4Yy5CiANjoz/04d2/GuyV0yt5wEu3Zb
81rr4Yt7zpXShmHvxWQP5NUkWZGsCliBbYhAu+gZ8iyDI4By7rGLfp4vrtYXe09K
EuKyPf6BESJveZln6DSiCk+93Cbs4eDyv2Tlqwi/n9B5LXIlE0xAfT8WyXzZ2Cva
a8yZyw1xPABNFAkTdIZzS0XiToR4B8TLv4ja0xm2AOriHO5fjQ1ngcXrPhlxoCkn
bbZQROGGO4D1QB/9azCgYwRQVpx1ImjxG2W6Up4Sl0k5YB2OQYYNXLQsrY4ON7W9
O/nrGlQ235PIOTd2qopuHUhcfKg2n/vtUnziqpqCoEA4R1aSRur0ngonG/Gdqzr5
T5QS3FMl+JFG+xPCie9bX5ccD8b9oD9vPym0c2gFSLNoIy/w45Qob0UQRHY+6qnN
vE5YbvtVyoetMhl81VfxEJb2QFxctJadVIo3PO4EIO4cymFsFaq7+lik+g1qzQZu
RaYAfWYSi0e+gL3MoygvUXH2WLeHtKuRB0mjBTi6dxSbQ+wtyhGjoOwtif6K2YN8
bmsdy5iZIv0OgV9tOoRchq7K1rl1VldGK+34fiTHwVBt6pe8j7d1VgEbJe9VvdlD
R0EjO/p1s4+5dBGXSOmJmBIecqdGg/Ae10dJsLBfseuM+scwhbUZNlUDTzSLRxe0
coj08epZ+f7u5HQIV3EbgyGg7F0giBDJ/Bp/Ur3WqFhpO5G6AcWx9mRE0zNpNmsC
2vDr9BP98OyYS6s+dfNJXQw2kJjuGpI7H+1tDL0FTRWxs1sFWFlvARjXJK2EwIK/
jkb18q1Fw0iOq7mDACmqSwuRFw2lUqPyVXpL9FYWOOEZ+Rq5lqwJmtZv6zh0s27g
eKPK9q1VqWIdpje37TM/DrzpbjpKFc9iLUdcWnuf0bBf/OtY7FfGiDNUk38uSAvz
X88/p+HpOiU56QP2bwDFcUdUtSkSP2hmhDWZl7g7/YIs2pi/rt4UaBwb2GfA/HzW
BMj9bTRMNTYLHlSPg/Ibicg9LB+x9AGdItb3ohhdIUgH3CwKvyn9OP6wzlQNCGYf
dXJmrMM8k9+l6Q0XJ+zgi+VGdj56SuK5a6dfX8cPwX9Gv+FnF/6jVFI58RHioe7q
oBZucN0eP8NkQZvrgiOpPU6ZfFvP82OeH+qJLnxr5X3VgXQmj4qLVreqv4mbnkul
wvEA0CIZ4wISLIAYryyeZcprhWJnEbBa5V1hufaKS0EF4bqI5b/CNWSb6+nGXQ/Y
i0AQkVGwjCSI81dQPLAK2X2HS224Pbm9KKQE4G6ylJWX1M3vUDJku2ZqPsKq4AXp
XPABVlwTqGd/AoH1PsAA+4Zr7MctmJNAYRlszTuM0wpAu3RdVSlwCnYjgK8/1FcB
CKE8u9HJRIzdCJjKFKuboWPaHCnY0NYqaSf9o4oE2IEBcVLIxoauJZ5NgDGph9eH
4jdGyLZZCwHFKg5LyT34Gvq66dCoH048994Ng+AqRQUUYebpfH6al2ZCEWilIAkK
7laklthHs1HL/AWAr+CN6fjkq41OPUAHAz77vnMR6GmFuw8y2ztN/BGcADmo9wBL
1Bwfizlx+LC+VqoGsvGwMnCRgqy8vFeMO19HSTG5nD3Te4ZPZrU++allEjD6Wvww
daHnVGvnR73mVtTH+fB7AxcB8af1bTzi2mjt1k9O9s4O425Vu5Zi4uD6mPmdwIw7
cAozi4p/dulYwnIuvt/r2j47jiUaOSbXZawfR4D972ePuYnFzY6Vr81fvsA1D3fP
8adN1HDxLsxoATRBpGgnn5ZV8JwsbNkcSI4Y2CeO3OT5/YDP1ndwZsi+cbvf195j
PtlrmrwueUG2zDt6AKEh3m2sYzeravc/KPeWpdRhzv2tyTQWDwAI6omOyvg5HZ1e
nM/LFT5vuGEyhnO2iH8SdpJmL1iRBSJ+9uR6DI2NJchdm2GTysQUtAU1nKtZhzmY
JU3h6v16FhTcWfjllF2B4ARnYsdX/BBRPVcfi+p8Qb8ymyxjSpjex7RFWs04aAAb
/dIjT/p44fLBVhfzI9ZDKSBQDUeSHq2AC1txMmfwUhdvNK6rVSwOZmm9bhb/fXSs
K4q0QTGm3NO/BuriWhzrqGkbMRjvnZqnEyjKHo8TvbiGd8QjjwEmHfpvpF8z6az0
z8D2VyJsxZlawdHxG5fWZIW12JteYV/8uBbFxN1Vcu5gWzoRXucUsQnph+ezmX0x
L1qv7HeCql0OPxyYRDHmBp+mGdYrJcgknw157dYky/T4LRUtDZwSbMW7mw2bevdE
uLCOFmM2tttgMnwdLWPP6EoQFg2c3kmkQpzfO7y8qddGIb8CiWtYiKXSNsvFXkPe
wkOl/l6buHgP3pF/mfP6rRguD9twju5cseFZSvID56k6Jr41xQLF5Kfv6y9iEm8Y
qe0L6T59Z6i+X0aqAXnOgL1ylE/Sy/vw7iBRNjbg4qezEsfsT7x16J9FMm6AKl2W
8NTcBcnWVt3Wa5t4ZPNioGeX7K3p3Qw3qUEO4WOk9ZmY9SfuT2c/RBQWvatFVYIB
Pze0Wd+D6Y36c2w2okkl1N/n1TImEdeXHmZ30uk7TTLr611zqTII+BeywhT6YR7Y
JYEwJ/mOkiHDH42m+poixDR4gEchABo9+aIglYUlCIdwV9ygnhnwUAHnHUDqwnQx
oLlKKWaCw2/VRrXUPsZTzTgaU0EYmayjoMwRUP9lwa8O+jd+rreNEc27bBCTcKRH
voLARyoSnBSwEzue8pIA0izUDwVmisBDlzZSrJv5g5K8cwPli1RPS+EqaoA4ZVGA
VlEN1hGV24r96ukwSXLjbWTLcqay+4zKUw64flwGiBUXurtCxNaTJTUruicCQMEq
AUgRYZSPrc8EtPWp6nmVYaA3Z9rBcULpuSBpbF7thUM6QHdd2TUmBc6AgHTSP/e+
oEandJhhzRpKVMV/DO8XfrbANZGjXZpMLyFRed+aL/Cl0RvxZ9fL1UQBKXpm3W5Z
RLoN0tKs8Drj3/bhGPT8djpJNC0RuPRtj2f4GkG2YzZi+Tq3IUHG2WVr3o2Uy3Bu
GAXo6tWotMzwTUDj8X2bBE1DuzTwMGaYB9Msbm+JsmtK/y95+w2tfPaG340nKbQh
tEue3FtkGt1CFGYjxqSg7kV8Vu8TDU/3B72y7wXny/9I95P0dpBKd7rItfBXy+1z
jAGcoYzRPa9so4FD/ivhNkqwegb6xrdfz1EpEKHLHJUwjYsOAXCJIYCJsnIe4w5r
41dRp8IcWAzXP0uuk6dHfVWq5kCMuZCxKqWCilR1wPUzBXmLxZ6Me3XH22hclq+g
erlLcuotO/VlHS9kdPOHixYlRNJbPi3SUWOZ96/AkakPINTD0mJ7B5aeNZrRlWnk
XR1vNNpxeJMpJEgnrhzA/2Qog4cUXMf1LTSdSxuza3vxBHF4Ei9XFwKL5UdxBx26
JtZ8XK88tbizMl4hRqGFKr/dVXLaXZo4TjWjSfqF6XlJBhQe6Y2p5wuI183vizGQ
T+9IsJKESpFwuTq2HxgYJOLD4Ro1PVh8QLKEY3mMEk6ZyZy+LWGwNgeS4Pwhg53C
+AdsGS7AoIcMWtRqdpqgSW+mYwIxg9dMN8NiYYymFJ7OGfSI7XcuTPUiYJB9GPib
qD4SWe2lirWwP5woLwIzbHDqz2oBlsPgWPpuFTauetAaFJowZ1BobZsBc1Vyz2jS
MnjDjUk2bCIAYN1gfNHSHyWdTad+ShCDrwnf8y/P+Bpo0nwplVpedWaaso1etfvI
0oFkZWkXVqxpA+CLMn83TQtGjw5f0m+PSLDrYFUWIufvbFQRLu/woxxxW/rKAY+z
91O75uNE5Y0BBnqpMc6sGy4T19ADqMsqgGEyRPwwOScsY4dpPFeJF1PYvvFl/235
CKwMbAXbUYwdfWx9WnUzvs45Dhbe929d41v/ykqFDlDiBrsCi68Jvfdwybc3/qA9
7aLgaDTp15jUi0c194PUDhXrN0giDXn+aMkuxoWxkyK1ENNtPPJzArlkSuDLPVu4
8KJMBg6BHC/flCvHq7iwQVsFXB6WsYJ1dsR+mouedyFHylNOKiQJiN3MkKWOpV25
+TJVDqYPrkVVVWJhBVxzzH/76y6h07NM/EygmwIb532rYA/tubmoces2FPnccR7a
QuhHvdmS2WL2c3Low8QEv4uU8xH79002DK9yRgEoU+5T6eosx/rChYjfwxqZNGWn
6CKN3D0uD9iJNWeYnIfb5n6gkXSAwPq//X/vxfzGD/GSJyKSHbhKsH4gEFhSS06B
Cfu31FhWs+VcVi7v2KUkKT1ueP1Kl6AI6TxjP1rWISu70fXi+PxXOLTyqVoakc3K
zt3TFyasjbx72L15pXIME5CragcQd795xBoGpJez9BUGpphduPG4wFi7oT9GbzOr
eSfKnolhN570A8E64m9aOf2VAhkSgLNGshQY2MiRabjbXVpr2ec3ielj6A40umgp
S2WbqQOvuGbcnf9KKfcHmZkrsO+tXtFFzTSaNJjBiOYCoMp1ss3PrRy7vZ5PJP37
UhKBfJUdAPEr1ONoknlqsD478SF2kqNDDECuAs0QVIPPZdGq4mCWhDXxiOzk1DQv
ZfitFe43MJQZO1QJPUwh3z9H4HBPHo9oAHsTqQZ1xCNJWEv5dM8g5fHGNMP295f2
z6GZewiJVLkrrp4dn8xI6EoZdJFncDBQg/kne1ns02+SIOj8NKXM7fiLtK5g8pWR
5xDoGpEV72VFoGNH4s6ca7JXhtwuWYdH2x2pj3R2HPjQ/V7slSTxddZyH4q/o7RB
PuprLCsE2pXon+MEjwuhjhkFI+mbUSPbIKlLXEoyQBbYIG5vuDiM5b14lfOJ7Trs
1iLNaoksmjnG7LvTtdbXNU4+rAAPvV+4eALhwqqrmrMbdLPGDKqe4YFnoFYzSWiZ
10R7i+OPhgyV+4Y397VR8dIpXspm0HpT/aN77r27oFkaNZCSKVxP65JfhWcAtZO+
k4fChLyG+LfWjW6lb7N/W9BBMoriwjkombvBc+HSjko/rPwg6Io6SKri8EFFyLW3
4WprrhGMedIus+4p7g40eJx0hdfnc4Sx8WMQc7lGcpirUvZql5Q+4HjHtDpHkccB
VUbjhbvjnMhgzeL/yZnqZ+W6ZfXeMk94jLwk5Sr4aNhZFGG3kiQBO3y3sR4smr6b
RK2+KZyxCAxNluGQM1Rkvli46OXYypawsRtH48uJaNCfqcvXxXn1M/yQ30pZG2+V
FytsKtbebldeiSrrKLhMjbfJpAwKSpzLGsW3+hQCkPmqEdDNonA7GI1sxBWEwfrk
4p42+oI1VO7kfYxxB1krHFCcw/Oqpbs9C9Ch16nxdNAS6vHIDIJn1JTH5AWTBQsd
34PElqB8E+hdwGyRE32t/KppAeimoOdGu45KeYhqCeLML415u5ULAOVvCC72XkDt
2gxHNYSBD4B2LVV5mqOpdQXC9EYpQNBHNSAjaIEoFSBszIJ+lu8QEJ0XfAhSydO4
Mkq4NJSsyHLKGNefZGPCj2OdttTrwGYsapibqgaxIhwzpsg+D4870P5lrkaqWfN/
jDC0lTwY6x6Ra782ft1rSLG6PelbBXvIB8Y+ZFx0I+gsh66KgyYgkDZcH0i4erfm
Rn6xdBpelk0cRuf8YnnSSEoO4MPnuJ9zOz/LeTr8k5F0d8gJZRySIZnFdSj/lBgu
PYJIyuxSGTCPt1MoY+19dz+rN95emWtO1AfPXL/Jhza+SpUYtzjCvF57maFyRnyK
Ia1Yvfi6rXuPc9ET6zSGGQHI1UcOeEJiSt9qEQ9Fpt0/kfBE10IYSa/qwzfZRMvw
tICtC5Usdl28hMyaIeYJ+66A9P+VcI0O0H7hcJjtjxgNBf5rWH54xKwC0YbzjiLJ
Ve6Zz0bgrMqgYTglMj/zbch5+ea60ybRN3vhYzjbtrVPHVkTaxjAa3ey10tJPDsl
F+2FYGNwUcQaMd8PJvX9aj9LOVdCYd1gRC27r8BYRuuQIV78yWaKykRDQi0yqJFA
+3zUlLrUuMFf3t+5PsPGgauH/IcehlSFMQ/i8cbTRkb9+JAZlB5NPxzpfnxu6kkV
pYTh0oV5cWOCCGkaDBUm79cnnDBBaWBxiD9ZgrYHKDKmqg8Vn9HIJuK6gCkck/NE
FvFkxBii3e5fhKLT9kdS49nW3xQfUxiHjUyv3t7A7jSId3YRlyAdAXGyJQzRpFAt
tO248jIUFHLKrCOkbWR8W3inpPVevRhEz3qSo9L8JwjdRzUypEtFayAcvHxVsaDW
YQIi056DbJvlhLyy1zd9b+s7ApD717kmBCGJmE5BlAYZ7mOxRigyjhKoL2ApU/Vz
aLr4asfBKeHNXeOHTIREUflu3Wdc1YbjVDdeolPoAjxclXuFG0XCLeDi20pRmURY
+6FKsevKLDB+3+0g4j2lZRNw7FsRl2dbsY4i22+UnHs8VxdRqyKIIAxKLp8J9lhl
+8JFMhmuEJ2vzFjsj4wQWOkPTEuIzCZYcTj510vzeF+Nvot4F5TM5LWpm2pxC+DH
incZh32c8dC273XBcTScDP9ay5VNNc/KYCaY89atRk6Q6HoQAHVzRkIun9MzjNTu
TQNymyyvD6CXMq3Kx43LoP/1bMZgCDjutHfRKScD74EdXFAEiyuVxVWrJ8yJNACx
wznmy0tObbbLp0ixn3QyVs1LU6OvOcM4weh0ykl/U4gYcQHJM9h81IVXKbwcDfOP
QnZmkMzgvfSAAOcsdWW8wH2GHUlJ6i1huqdJqNcNkxwa1HEz+a636RX5tal/39wX
EMR/HtiVn8dktAjZLTUokstqNU21C8GRmIIaFl6U9JCYABXEMt6HiASUjVWnGU60
kWtpYH3EkAiWW2C02Sepd/zbqJKC4CzpRVOH9N4hEzPzqaBwXbL8ajwJ6bUHwuej
c05QiGGb8Rc5L7Uy4l0949KbALK2HJ0KWyFycD9FmVIqjLklZVql1pJomhDfbgdZ
UHOHgO+afgRLJtHDk/suG55L1eUGpxEnJACR27HFjAI1gK2cTDocL9HyLFaC/9SA
ivN2D603K7NLTkgYf7tigEg77hLIY2b/s8t9e1gl4VG/G0T6CjWk6mqaBG/7kXDh
tnZoW8mJw9bVdLJlM2MFHadUGT+vjhdzB80vtlpyQXTabPLf3IQEcR2j6y/v4iOc
655ytgXKaM0iCqX6BAubm0/0wXH266IcB9AV52mjFSnE4Vqc6SC/CTOjIu3L4uy4
h3eDGU3aSnrEZnkBL2LwoMB/vbDAdbtvT0qf/7IYsXzEeyVNfh3ibazdciMNqJBX
IeGMw+0kfFvtjGw1SBgP2ev53Leo4dh+AGrSxZU56wKX+La0U7s1HB6M/2z82JJo
Aj62MUM7Ewl5mUI87suQ0vUVlTnd2M2SRKIeaxcw5y6epw3qoGOWZQhFSFYXp4H7
y2x6SPZg+4Ik2QbEUSEP6TPFaYI0VqsXj7SYNRvy3oXt006KxW/NKPXmPXH3q+bz
ojAga0qY88xywjjByoJ4UFU+OscSy/U5c0Jpxp/8BSFu7x8/tDcHXdPtZbN2sODd
qqWSvbwFLjguRReYoYCRuy5BbVrVA4LPeMnxbWHeFg3L8+vGCPHh46UagKUDtzw1
T64iprwA/l0QcEl0/C69CJzF3M5ss5tdmQXmUr3RS5lTuG6+JO7I7wcrQd5q7BI8
t0jdBcStCHMTaxknians4yN7F5N59+cSQ2mx2V6Pg/TW3z+MV+ZVNlZVnjXL0j4T
/B0quAMQi77l2wjeigop+LNTWoV+GwCb+2rKph9hhei7QAXXo5M94/u+5UkIZmJ3
s95LvLUeptj4hs7CsvYPiF2/UHuvaWsIdZNOGaAj97EiRr4xkgyNyvujW7F+Zb5l
PS55onRiGLvPk3KVNYITVCgniLcANo0xL3YrV4+oZAONIxXE+QYAoRceDL2DVbTj
WwCtP20hKCua9g4Ulblazun9Ur6JBL1CYFd3Wz2ZfmXUNjl6Jr1LevO13lDhViqB
3YVPOPK8J3IrG2IlHPL+lWXmmgRRgvTOYs/q4WML5bGdk2v15iraB18vQw9bAOjI
/U/JvjNGqiV8cj7OBd80e2s9BL+2O19EQQMfX28qdtqhomwF9ykRn+7lwJXIZT6h
qlR8hJLIC1gMib9q5XJFgJlUnQ5K5/8vcrnQS6SKmKWCcBYVRdYlO8HLMeY2j1qw
ihERKN83fn95tCwHv7z6vtbzZSOg2uq8PV70iCkG5QJzl8Rk+FeLTWYgKl30sPMQ
4RgUf9ilu/zvQ5eZ6X/SEv9U2Nzt4uq8pixWNMaYzTrcG37xSa06fEjz47gfmaWx
BEGpKQ6osy6pgZmb/Ah+weG0LtumQNGmUNKGkIXSxfJauQkCiakg+5Wute4ZJxIc
oi2WMYTi51gw43b5qpFg7A6t0NYhMDzFZypzVMnuPdhoXDCmkeXnozkgV811USZE
BkiOANoA75g1GAEzAPxqIUez/GRo29u9HBdzJpdtU4gnQ7MJELmExiYsj6Bnlwek
V05agZClJ1HVupQ7oUqn4bljiqHmCL9KpJwDDRFdyMYUjheFF3yj6XG99xKpiQpe
2OziEBux0Cv2Ljqt5pD2wkwZ2adkcbR7+7skgfudlPYKySK1AActLtEpbvQNEHw0
KqiXdrj0adDfb1DzFUhBsEUwPmmjeYyShV16EIEESnOaIL7C0m7LRcbFJmNwNZ8/
mv5oIhbriW68flD23vjmFPIsjCbHsG77nPh3OPeQZEThGxuafF1F194qDEVa4Bcf
/LD1WjbUS4hQ7vNX7p5hdPcCarhomRFQrk7R/LCva2mgOIg5g5HFXsHUzRytjOsk
fJrdxK0UU22ql6o7TluoHFK82V3tmXTdkioq84qnqeu/2DKtOvzJEfDq7aF/bQMG
WzOLICKo1RX+kezXHXPgSTZ5PXkz4xBU5kN15qlcaMluRKZS3uzt9q/aHY2X8LDX
Sr1Do4D/WsdiQOYaOuUs7HMzmfZqWCAvNDuBiSDgUFg4blHp8D1zjQzmhaw7gucW
AeN/tMXg5tcVW7fwOPaUVPxW2TBJ1v4ZxCn/DrEdeCfXMqu2nkGt9PCcE8HWtlU1
GIW1d3n+tTN+xzgrUBjLc2f79mJLSi7hnZSOdgOFCBR1mA+VTyZ53Ex/rREDQKwW
GTVEOihYkUG0HWuXjX4Ma64ocVmFs5QIIwbHFdHdkaSS7+BGfE3imzvwKQ3+p+QL
f3xRMXaIZqR943SuLiMg+LNyiD1RhJMcGlQr3YqWltullFAcj2Dr3A/w3JCbHvok
2Tt5tSiA4Pu5sB+cHnFcRyMR+cAQdaULeM8hhW2+LecufJ5GSijqV2gPey1Q7c6/
GMfQ0Ct3NBX7d7FvX0rrMfQR25wAUoW4Mo0zNgky1XtsNWb2aRyJU4HVHxwCN26q
9wLF/3jIbdnp90iMRZdk4yJ6lh70C42TM6eoWQmKA5fPkGUz2YurYDTIYMzSb1A2
MR6qfepw+xLdxzXbLObr3+soJOj61778L7lR66rS0cLzn2+CHKfT+jP0jAaoOWLm
2mY3NhpaTLjDkezVLeVfxor36DXC8kcU3uaFcmb7J69+lglyH245OCBIhokv5Mwb
bHRVdmaTC2zFzVH0SwCyfRPqd5UIBo9Rm3Pomvak3x2eNZ8MPg7f01oe49FJyk0n
j5B4/OpjBR8iRGcmY9cfn3gcRrBiW0Dz/3GlCavRcb3n2CB5gIi3nJyVL5Cf6D0N
LPxvfNXQDpTKhtUpR7yluTnMxkIb8mIGoUPt15AXoQmONmwq/fU7/Y3vPr1a1BOv
1DERm5koclCOG7NJUjDAYmKbgmgwn9EVS27u+tzMN5cm65VfFs6t6gMHjepWqDnN
11nIolTe8qr9ZWF3nr4PXm9YFVB5r1mnEskZsARLoj2RJk0FlGKZwfifiDOTNVcp
S6OecCdS+JtZmLHcYIVADmfCvf9EkxfUeZv/2uOq4SGCcMsYuLZlDUpoDFBetnkP
FI3nhT9LREHGG9UR1YhN9aA7I4s6VWzm0g9pQvqpb6Ou0VPxI4ym541GV75R+hbp
3RSrThI6lQYi1ML2kd/2XP0SBmMwTuLj5UCK+aU6oe+ODYkFmWSBxtdzUe6HEUeO
G6j85HoHuTVgfMR1UYhEv3ea/HxUGEIGXEBVUuxR/aARIxNB+ZGl9QgmIt7/h3jx
kTHFzusPzbGUxNuO2tK0p7aiAGbGXJStz1p+r4eAZQ8Gh3tMaZLSTddw/DPlZx8b
r4ma/idalv4q/LY57LU2XS2IRw5biUUK8SeQlgMlnodIzFs2LGMPKcBH/Xa1JyJ2
nPrDa8ye1euahwgTVCRvXgyF2hDdC02RJDXczRRgk5BTvf8n7lcMJWDVMDgWkOR9
LmmfxqEuPFtfadfmAZMw6ST16P1M+5+eHkNO3SxHuQXxzvKVfdU38PqY/KUH4LDq
30wqkD8R1yCJI4laMlwbQpjqTebJeV4W2+279KAwSri6zaBJG1J6R8XfcjvRltk8
n7gSazbIukqr/SwTYtSxLMELowvNOTrb3HUoQl5E2nmWJaFwPauaJodyNgraYdOD
G/57g/K9viwTSA4b6uHzdJ94PtMbCMT0tSfyAWjkLLl6cx75xoI62vo0sMaYTwTE
LnjOV/l6b6P4XAoKwC8fDoFDzAW5fYJoulvMsJgK6f2sfWNG+AL4RT+Y/LX857bc
oxiNc2YRmxaL2Mw9TlKOP1lgTDiMbl3umJ9tJSikOqY7iQZM8xG9dPmtfHAo8oAU
764auNmkag1ITHvb4F0sQmf8VFN0RZTerkMrLpP9v/wOQcpYKe6vW6ipudUEFFev
FK3KcZ6iJq1fZE9X299JLry2mrGOYze6zvsymjovHgD6MUdf3FsCFJLHzmBUONS/
h9E1GHBxwgXNEuOdO16jv2y5wGX7qWOmXu1GSwAkXQxnRqGVVq4baM+ZW68IOX16
s9Q3uuEECTRr2mzPqD7m6qN07WXmkWEImFxJfPY8D/I/pC0lBagNaX4S0Hv1Ggie
D/EdQmNicFTLO+EqyplkFi7mLUYNscZL593GOIftqnHV/HcJj0CbO/+9e1+tijcW
XL9LE+Sdf2jNMludThRNYp+lMoxvEJCzTzwUmYaA4ONeNdPGG3rhgeS44RsAYF2b
5Q2SOin+gSZjhAgDwoEOUJ0MXDZ7hiHx7Qs8ADNi5Hg5hG9Aoa3Q3gYLU2QBd3LI
lsbde8ExZAl3cMxEYfIQ0dQhpLmW2sbwPp4404iMMmLnsmJid5upnC1LBl6Wu1hS
nIZZkssa7ooikjZGocZMx9O5HbR1c6uKLj6VKMvuqJRe01wwP4J6UIhTRQUHJ040
nJwCEaMZ76mUp0gL5bNg6i7fmks8EnBlmhTEySbY/bJTOTYD5GvZosBlfO3z4D4+
UrBhtMewBjqiiWbzvRkONcmrLwRQT7UellmjTzWlBNODaOcVVtJztXKvRuM9gTHE
9KEHNoKumZZbDYzFGMhfg54CIEfXzPasghlax+af+TebAN+9lQt7CD/QmPJH3Xpy
ud+VJtrbnhWCl/Tf2+9CjVYxpW+P7HTN1KVkvl7cuNY1Tg7UIhULCeOm+iZVo6Tp
tA9vd/Ge34YutQ9rxpINymg36NV7d6sD5w6flXw/k3r0UPJEC5b74x6qIpW6Skxl
98ZmsYlGA73lWKQZ7DagOCbgLUIEknwNBI4OULh2s45DWsrfhg0Vy2cegIIwoeCn
H00Ev7qqdUJBAQTGehDexFCg9frIHQRJ7acnCrGGSnQSNvG+u6SBZeQJDqOqdD/S
C7I9ScMvAf03pPRkOus2K7KxUltp7uGlwxECJeuhm1lopzJeX7pv3P1SdXEcaFnN
tdjAx2QVsFwtxNS2BQQlcdoWOGlzt93Ev+ofpS6gKAKl3utgx68l8QFtne6MlFjd
a/0ox2o7LwVN33xEFVwaV1ghRhSWvI5+iAeelY7PTHyLIKrXnIzcG4ZJ0qv3Y6PM
RavbqDcO7F8tfAze3aYfrtj8zFtI4Tc3hUWgd7LDDUamka8lNC+7h2ViZk4uiaU0
ShysDn90E1u0dGKH5wBqXS2/kP+1LXzmSqHkp3PEP67Ny6ov7eEub2tvDlU6Yw25
PnLG6qcNYuqBfs/UCl1E6SIvkO1W5kGlbVvYmgIrW8FE5Pmh4zPUIkk3CNFc4QTX
Hfd13+r2B0qdChoWpwfFfnREcUqpU5OYMeE9pcC6bz0/Yjewa2R8FpADAonBrqCx
UAftHnqNY4cd6R0olPWNqyv0hkOapvTcBuYgciFpJ2/MWQSIGD4BhVONhpUQ75+G
B4ugpPkyTLCzTthUws0fESLylxOlNxHwVl5aP/yjxLqglRfHaWTo5QJw1f1JMOKq
JAaoUzK5/ZohgmOuP+ztBSvw3Kdb4bDOrdiQhp4SPexBan0cy7oZhwKLmJmX5dW1
pCk1qAgzQg+X13tJzvMwT2LEEe/30aFSM7uUkgAK4RACmAhsI2HAXlt0M2c1P3jD
M9I77v0BdgO5LumP3iYiNYj6tMCrUBV3MbJW8zGNIV2iBHtJx43h9zX7H3ug3bEb
3bf2QAoGN4BtZJhe36VuKPvhNGKU06KH6nxsr2y1ZI++q7QztQKubPpUVyeIfbW/
X/6HM3qm0fG87d/J/Jqb6p29brAjmbzpai7LL4PBgPTIOp1lhRlJ8atv0RLciC61
51kpgaScleuNn341DIp4hZoQLztF/RE/E2/ODoqxqtLfjpoWPs5Woy23RLr0VOzC
yyghJIv8EK0k22mMRhdvwppYI/MpeDIdv+beWCh/K4MeJVjobMFbLcQ2bLfZI6KY
pMPVDtiSNGsdtqSort+PPoF11JIOIYtRfIn64Njtaa2w5Fw6AJs7M7mbv4CeqfTz
gpnvz8f+HhjVhrkCsOtM9RAbzdisTN/cCfv1WoO82Q0KgFc9pMEgpOGkwS0WCVqW
2/EMuplOupdWNpUySU9ODUUl/cKJCKGMOLB7KDmdAqQqMN4NENwoh+4v+cfNLuJZ
0Hw/1E1rYaMDoRXXouqLTDW4asaulQqxuq8BD3ws31HTg5TUn6st0QXx7ufshFK9
nbLGFlZug+3EapSXedtC5rvDME/54gGqdPFp6T6cUU52NGLra9GH0pe+K3S8Vp1J
xU9rjsDWb2HL35aAsGiFPZQjmCK5s0FIJVy1GKToOKlL5SNImnlYRvUU8xv6GUmt
YV6gqZn0p0huuAegXGFUewEr/fpxbv9h9ohf3uFrNWa9OkdGDkVP/JzvvQh+3xhx
ariHvocCRA801cL4tKjCVi27a35Y040kv2AJlZ4/6MVKDJTVO8E/W7pMjxjS0GGK
MXZQk4v5ZJggtFTIeOCkDLno0TB4B8EDuNl0oaGrwixlqCxuyJ698gjgm2eomY2o
0ZIkkM+Stp8/Azfb12IothCHN9YYBmCFD4COGmDOrDWWUD2mGGYXcC6usZVUCDhk
4WCwfRS8gCzNtba9nDOeA9gqlySx021qlWYlbaO9N0IbK8wz8+wOoJSG1A8GpfUv
MDgCPggsMEqTYuluRvKT2pkfbYMJwMuqHBeN6C8mc2OQKNwMwa7vTwW4JLK+AfvG
j8wVTOBgK2njy7oRnNbUXp5x9n/naVPrua4Eo14k7x9EU6Jc53PhyHqrKGFOD9pN
LEZ3sS1M+NxzVRAitGqIvTn6scTOw90K4zSLZAiwx6NU9oaos8W1hHFX2Vvr3hdc
0CeMr4WzlIheGJgtZbeXP9Nw2hlSuMu+ijM88W8ef/y/MurNfJCAKSnjYmkMx9lU
2jVRiXt4jvvWP+29x3goIF/RRnqZ9oxYJDXU3kSeQ1t6DewifcyATyNYm9zcttpJ
ZiMLe56V3k7uIMyVIr3sao8+NaYuUyxZu2s7i3nHpzLZU8JRj4G3V36g9TpyDczm
PFtNgw7mr5ef0W1r67Fv9D/p6K/3FJamrSA+tDkzrseu0DmnxYTHz0jiG6iwDM7F
8QKpb26VERVXpLEkgDQOr3MYIww2J4h3gLRtPXqh9fC+Jnrzc2AFst2dNck6nOhA
wXNwLNCLl85sP3XE1Qh2ppxdk81NerZTigGgAejT7+HvuzoTsRMClculepWxsoHg
OVyhySzoty1sl676dYnKvFrPq9pL6b201r0gM7kQsYJHqYaSrSUot0CbI1Uc8T5E
gIFcrCK+7ctkS1wr+CnNb1dTcghXpYHXTeTmLVhQsaezqfyi4aN/O8+unaY03RB4
5h/S6Bd/W9CVz+Qhhw9PWB42cTIpZDyHCiXQXfZ3xVzm+BY2Z6WfLV6HDpKkzvKY
2ZTmCMygBLxdIMAMyEIZ8Wa/ryx1usth3ed3QlcwMLb4hvLTPX7EeZY6zEWrb0KG
DX00hCf0ksJgamWCc3UaXCUHJLmKYXDPN3i3458frCMmaDYL9W8ctez3GD4dsfeK
gV5b3cPY/CwMYkZQir7X08vbptoSM2NBFPcbADz9vujoVFn81ZYLGY3PgDF7cz2D
G7zPk26q/fC9s48I55t5wNVO0Ko9Fnmz4YBW4LY2WdpVNCXwCNwP5kcQDdMP/vKw
s0HCu7gAatC9obAvl6JnXNqNn6ntZxr+PGXBkd4MUVgx7CoxjChJL+XN2CN13HEH
VZwpTtkfkyddet0LHeGiuVOzHctytHdskP3M3ZFndWRtEV1NKLtGyEIDRWQu6kBp
Y9mztPzNpIF+HXw8v5lD+FxNZqX69iG22BUO1m8Rfp7FIMJNhWmMky7qZGkvBCe7
3qYEJTeS0lKLOvAus0w7NIhAxq3pxf6bashtVRkLxheGUVsV/6dySrwIqscfUJ7Z
hDS/aQiWhGciRH8G0haC7a1tEGVvlFLNewQbszHxCZbtNRqeRtcs6d+v8Tzl2Z5I
d15QEL/r9LTTmd07hKisNSrdWmJt4FHSfktCr3sfT3sP2sibyO2Dw2HKnM1PFn6F
fvK5pyIt0p6DAZ5iaOiLrLnFr/4mStgjcoKGFWRY4k7rbumF1tDWCFH3qdvqXfFS
mZNgCgLbQ2X0cVkSzv9f9OWLe7EBXStRKfMa3kUtOPc/PX4aylYx36jesns4/Sxg
diQNq6mw3mT9LGE7CR+8UtD8S+hnSaC4Ui9LIAigqPLZy7be83ySLvSP6AOmAoVf
qGcE1wqmNURG4eQyYjnjRxLmJF7slJH0jECeDIy+GpPeNPIXCfc4rUOUJ65AMt4B
XXIu9PkTGSmkyq7n9spFIAY1t4o7/wYVCqUTAFkFQs7r411qh0t7By/9BkH5lhCe
q0Boolgg8X537kSobcO7S6SHVL900XLengKy5EjcE0/XF8b+Mn7QABhWekVFvN7G
9Dg2N4PkOZpx7/X1zdUjMzSCqTw8gzeCrJD3ZPDtOHkcfqc4sYDiZ7bxjc2tgtMs
YA9MS+yk7y/j9RwGwfE2Oesktx/dg6DgLc/5fP6F4mcOtjV0+4lc6UHy4L9N8c7n
kOaNSy8B25G5oc46lsfGMEsjfeP4zghIrBpY+PVNtwmrWDXsEedCdtN9RMJRo5Ut
nt+AcqS7OZ4zWjCzwkyMEcjgMNOK53c0cpm+d3vQ8+2T8bZI4DtjAAM5KBh2cIxu
a9qZVtEEXGzrctvPxOHLppky4ZtApe7GPmOS08T/j1QHCZFLCYXopGnukssum3p5
h20uFtexWuE6iuT8Tc9a83rXIgwiPstZ/VMdFqiJVeccg3qiMyFgXDV+S+OIOIF/
99cuK9/V4Rd/mgyYGfgk51yrx6sEb1gu8kKS9btV1dWbT3HdfjgV/tRgzuwDatfc
zjRZ8SOJ9aUchaPhAWb+5xWgTCrDOXaqddKJL7pXiSBEI170vfWWsc9gXrAWvzZd
cOr/lUc2MjZGg3CiII5tMx9e2XDF/Txqb/6YqEApLzxAohpcpKvuU23lmD/Tv6Ky
WDzkna2nUSajrcee0IRNk4X6bLWmNA/zWLy+C7gMPgYA/Ej5sMpiGFaKsBMXK8cF
6PArgvo7djOvu1aBnOpVpfxwffM3nVBUfkTg6fb8xWNbzJpPrYve3z5/D8woGp3O
twNrYmLMyQXdpfAqhXpM6m/uKYk4kuEoKOcEYYeJN4eji/FEcpTcuGfX/hFxX6jc
OuPJRHHwsRNzNSn6pfAVbg5+Jj/OlUEeU12Z4fyp9LT7Fm7wVRHKDNyG0revFjpw
wgGH2BhffIYx9cKprFSPNTGYdESGRNyoPVcvqHxXOjvDuziwRIQs3DBPIX429ptr
iC2uf+WFNDL+QxDbJ/WAngA9U2iqpvebHok/3DH15G+PMvQCuR4lzzKR9rMgmU0l
SIfZm4mUZVjcKPE5eyqOeKZ1r7+0B1QT0vQ20Yu/ERL2V0heBDBig1uWw5r/RNF2
crCwpmk195yKV6tQWu16615Y2EoKsiNqko8uC3WQPRSirAe62Q1gBMTqaNEn5w0O
eM6W+rummalH84FBPgtS9CcMmZuC5ejETLhEvYjICp0+yiK2fb62sRBZv5VZ9L26
HOvpfumKYuzZUtywGJkZlkdNFU0bzFSRsmJiDauWF1/JUY16dJO3YWsJ90g0v5eu
KrPT/C4K+ac2ER0DI4ezZqYF3MfuNWeVIjw2Gd+PbQPv7AtAm1QppsOuicz1nLAf
7UXBntVGnRs7+5/PkmauXrRmXtlg4JGgPnDWc+cJLSSbMJTkyMxKmY4lAo0oR6+E
IRIEOOZxpMQIRYW5fR9Tku8/9wAg96EQ+Gi9BHOC/QyjCJ597qZpCIvE9I1dR6kX
Fi28p/FnDhNCgPtleDaHXK/yN6iMHcfoOVADfFbragjGODmay3EiM2iHC3eOrKrU
akr/CUaTzgev76JWJ7m9Y5KmD6gnLkhrcogo980RS78CwbU/BRjjsJmwM567XugN
Fmh0pJdwaBw6PWxSopQ9uF5LPykkYmAJSeqLzh47wuPB2x6nJcweEKH1Cyu4o7Ob
Vf0PAoR0wWgBQ1c0yGtwlvFqNEDrzJv0CbqWar9SCZtCUnunNvMcLnl3q7fgccTZ
QbV/LfzTxbEjyIGdcOyakpZYRiBCjq1F4/ssgFjTrnXI8KbwbCBzF7aLSXxF8QcG
yMo0KTarI7i7HiecAgUOikg2JmZKTE+At02YZe5w2XXE07oNQ41AVjz6J7W8rSBb
4EwElMC/e17F3SccQpIKr2nKRb4lygucOJHW0VA7zRFRGNQbZTJvQ0iFWCdwv7Lp
EWW/DUzthCnJUWAwFfiU7QIUDYvBD19GZYhU7Htmb7vjAcJQiwIymJ1RlIsGWSfT
5T0BdY93UkpEqwGQb3p+bEezbRzMo2TVie+fMPz2Uxkl/z10aOay5FIKWGJlDOut
TQm1/tB6efZNzmFMN//m/l5zBF82AY/jtk8Y0S4SsZ8SFm9NEC8hu9P16Er1YxCi
hPn/w4gxxlMdQhUv9goBXbBNF2/I6B7tmYrZFLbKDVmZ7H/KvciDBxxqP3gQUIV5
/N1hKWPicjo2ZpaM6COgPZuU6MCojSYVzLh/WbW40SMvsNVZBJN0TOLHUF0L++eV
t5go6nT0WfIgu8NJoXScVmqgMJPP8AE8HpMbNbCW48Em/5HwKxWoFPsPHt7SM8uw
Opq/2UUX3qA5RA82maeMmM40IVYt1AwCF7l6QXaAWc/lutBmKPbcpIm/dW4pGWHT
PzmhpoS6xWfJwZJfqxPd8cAQHCC5cMXtcaLzYmURsWfKIP4A/9MglyxtzNAv7dd/
/vlQgtn/QTKiOsBRLEuPll217FXijQoXxJYJVff18PTCH9KmRabt1JtvJvTbwrYa
gjfhXcQ5GN5x2DRtmg4MF1XS/2950FlrWk+GLGV5DELrV4V49pepEpA4cHyNNK/I
P0ryRiyYhD918OIATEHkQWyGlGPIPVNpY7WsVEPLnLsTLbY3iuE/7biRQf9VVEsx
+yJG+FNtwMr3ahJo6P69OD5sigghz4uoQKugby9YEUkkFtUzgp3ScMS0qHHJUFxI
HTChFsONEHxuTNFcKkMu7KpaLuVFQxnxsmXzqO4SK+Qtp4KbLhKsUXxTLxU61XJi
XhLjo9Gs/898qlcZhpvQm/b/8ofsQq0b75HFUOyowajk45z0VLyzflIwmNzawO41
aMnJnr3J9zbg8XaVe+GeEsfeWeS6prLpTeU0i6K5VScCnwQeHfxZqJbHMH43h/Zy
RCPxHH/MW+HCMSfi6Rlx7yYvtTo8xuSw5rFNep5s+Hr5tEpInAboOxp1pEmGa5qh
xQvhOKNPQllAauLR/STDlVhC/Rh7/h+5EmZ5dG6qnUPoKKS9JVAC82AbHCy1NHy0
yRcTM7LDqsFqubGUv7jSBE7PjCj/XLImbNWX3ytpNE85MKzrmgbXcMTV2lNVVJCi
CdYdsg091ADPyJrSIJPRqxo5PvTi0hmpJazHfFOmw9HQ8cp9QIIZhUFkNPeFVPPr
IN6EzRG3idp0JinCST/dPPDe26HmxhQS1v6N3OJKqvuDGke8zsH/ORJSZGl0DaOW
pUlpfzoE3/Gfwh8EtplXcGKtz26Mv3MhVY/EEE8bRjqJUpT0w37M2jOFClNt21Oa
9jdr4DWrqHzyo0H/I6DZ/wOyt+wCRADnlgwArhjK2TbfntM2kSihK9oDzVNqgYaK
G01n+SLsaxstCaLs790g7bhkrUfag3jiEkiljI0d1TvX9Uzxg3yBFM7DApXHBmLs
mmVY//TVWR5pc92JIZsP5nNoP8ixPrUhB+Rc5z3q3JK5tEEe96wMzbpiIptbi7MT
ZNex5u0JkuAYJdBuG9i0OnoEzUumXNbWEFJMj/h7ExH41DpdQGMxITafM0ZOde5A
zuX6avl9QgJ9xn/C5zisG14Gzefo4k3ctDI7pICe3egsKaENK1r8pTWM/iNfqkzC
jaZ2kqZt1ij0jQSKHNprsgGTEENNGH/TFceNFz6oa8kFG0ehlDtH/VL2AtC4b2K0
oMxioomjsy+QbByK+QpwPgcZom43/Qym+4mcHlCLXtVnHtPKldXIcKYqY4MuZEsm
gFhfTaDq4Zo5Rt7YFI1QKd13TcUP2OVEvwz1xCCax7Hj/sUEkRsK78qUgrDfQxyD
c0OnxPZ/Dn4KecK1VIAz/D9WtLAa7YBvczw4scsk4Oq2q5oqVXheucM7iQudSHRJ
iYaWEaq4tqvpOfqT1UB6zhYKocU6UcGD2F5eVbktVmHJNCYqWYDAU3zFhk4s7HuL
C0xwUAPvsuruBriM8OJ/rgehgCVMaNf8WEgT2UNNX2EbgW0B8xYnFxjMZlY4HERZ
SFMV8mbJj2ZzvqznY8yVTYyClYwQtbBK3uKRHQsttQDOJkwelokB0mVWL91aRmRN
hKGLJRMj2YNKJbquj6ndsnSHhGYia26YY+kMt5Y2UX5qvcWqS1OnjI5mNR2J47F2
BcTcLJfa6OTVjFcrI+HbgjT/rmvwZlbs6qnDeltMzChIkFogDwfXK61hvs5otZRS
HfrhsaM+LIvu08SXx1LgtZyIpAxHW01QMmlqzbKnsltg0eelHkS/KV5QKPs4Jx4g
aBzfAciLSDI4VEJ/UDKZ0uCSHK09MHWRZY+Y8222vW85kf1qpPN2UyrXRnIT1q1j
qQjciT4izvWNQ8cwaYHVtcBj3KAgaZlkUS/gwROV7JyhwdBo0rpdCAw5HFUDIoNO
tceQDyGGpcqlUSvoll7NGR3+PCyqwo3lgW5t+irJGcDRADfudhZA4lgQ7rJ/VkCw
RnL8IiDDERGkUxXF+68+moNnkfLEH1eZwuyrKxlReP2t6Tyr81xiHdeiyeYoMBLj
xxlTkBU0P1mNqllE6cNThnExmL2EbP7sVrYMBciGCyX5rMKRXYETtAP0P+T7R7l/
B4tFXovZr60iVLxvyRuNEyp1AOATulreVZyxptceGzbc9gBis2rPxiOMMqa9XEK0
lBhlUkIcPLtw3/3XCg2OY/k4tU1IhnilnQ4h9sr4a9aF5jBy8YtAXCp3sN+VH/Jl
nmSIXeYqaen7Q4296PnC2tbjsnY0T5lIOQ8+RubnfCtBHbulnylVCLpeQZOx3xjc
0G6Y3JkvuAUJUAd3hgxTX+ohYuwQL86OkPAFttNmBANaM46liOx0PtSOw4uBdFv9
Cq9rJiJFgX6JFVYII6idRL8GUjEMlRTmiRu03oLTCVijiaSInipFs0MGFrolPZu9
biITshGHBw7luu+kQlrTD2ggA6KE0ChvXrxS+WZToeg0LykGl/t1K22Ii/yMM333
lfOVWt8lNGfBmi+aac37U7n2Mf1nZ19uKMH5XTxlMbY4x4L4LZmWKLDXEb6GQzUr
HJX+STFjvkxvAU/wi7nKuvNuNlQm1FijeGLpw7OM5IZfzuwQyC/97WBfzfaRpcR/
DUharR+ZTWXqQCCfE1JkQ8gaxaGK5km/AVz5i3D2uWYyP3f73zSldLYdQpOEI/27
RZCpLvaXkisfRR5vmO4+jD5czdXqUsToylveUwk2prankMizKWPwfsbjM7AKlCUU
q5kXWExzWHJhhGhtuKR7DSIXvcbNec7/wT6d6ZCyJ23oZnlAvYgc0ASIgItfYfO6
PCLqvQLNLluDuc3l/ibzY7GLonZTd9V1PEQaVzwp89vLWYwgcpGWkHdHr+sCaAGk
y0+t26+ODM1LMivKvFLl6Yb8rOk2FNcXwRZfKBOBwvcfwzHEm+Tm5UudBkhBmpkK
liA/8bHQdmYXa8b499FPdXuKet7DzOjgr9mlDke7dOAmMh0Iq1Eo+JHbyE6/sYUN
MiA4C3EXIPOV8DhSJtLSFGsOlm9UUlIJ5nVEf1XpKCQmZZxM+eZ5mM5kK1LvUCmY
L+PnDvy4VwXrylmIRG887W+6ZMGBBoZjk1BQsnRAF7FnX0av9M9afxHs/lt1JPQL
n9a+2pCZcaA5wQX7fKVZMJUK+4BEvUJT8wx2DSsgAV3RR71CluW9FRbtlaoJzXMl
Jutr+iEBRKoDVy15dmNJ0oE7rQIRFDetMGOhcjQUU0poMO8ufvWhPfS81QBlO+/l
5KZkxiyq5nXSOU0BiU622wF946wO+n4cm9/EkdDLrE6Zk3ZZRajNinL8bs3Pr/pm
XAggqF4ILCvI+my633Pv+n+FPQpXG6AnnQ+/7H/nneKSjRw5NR4+TcdOrG+iyPmU
MQ7CylrMMn0nYVhf5nhcXshal3McPMqP/YDZEKkLb34MxrHcJ+uKJ706/s7r9+vX
RXvOhsUOAMKh7dFIQ6sLZ87CB+B/FzJx6wqKz+YhqYpm4gU+wzCVRybIOS/C/5YL
H3vE9+644Zoccke9dnqQnoEAzqggdOHoSxaGATX+5Al/cu+JQfZNkRZfPJ/2alm1
YBrPeShBHoui8B3s3e0fYqHa/p1Gxu+CK5zjsdxITaBGAVWFZXf6OzjQFVYJUnyT
W9hVj1s//At6TRrVB22ie2eJCMO2mwNfRIFj/XdqgRtC2zjZXhWO1sY2bgB07mXs
p5R0cF+8puDGPk1X4zffl1WZqvaT6H4P0yYwNBv3OzHJqwv1/cc5VPBMFCF2GE64
pk3/4/szbOpIDhuL2nb1LSWiDlF/TrGrwj5hOanRjSbdOgN4dv6hkZLwOpC8+zhy
7GS+0tm+MeV0/3qSnUneaRxXVVqNhtBcORwuzr48cKruKzkp9v4aporaxCDiWNew
gSW8MUPfusQ/tYNJc6j3L0hkN+ViQcJuVfZth/f8XpYkcf1vg8t8v2V/vp12lR4Z
gPojSrZ//pV1OueVvmFWdOAC2OxG3KJgkfDkN+FMsVA9m6AbhS+eo2daWsq/5Iu3
2gtYPkF9JNeYR9qAdB2qloVrVMWWwQnrSKA6BSTS05+I4xtv56KU8pyb41hyoafE
gWMqvJcdY9E9yvCV+o8kxqUB6NX/YivFSMxpWPNJcuK1lJRQh0WtdGkLk34lPPB8
sWXVUK3mW93aF4RGup4puYF8yiKCHR9R9UQzZ+aj7cXsSo1udGAzWUMY5b3zBQ+O
p9jwpV6K6FRaWyneMM8+jacg+ReUaF4dK7jDHQAohaB+2yWNCyA7aku4wquZjeFR
MHjDjqzvfVrgJlMXfZMoQfj5tbZZxS2DfsjxItP6z8WOA6hoBRVhNe6hw4D5uSkL
+Tnlh7sCza/pVMUQSjMFOw16idAyO3H0v6dA/Tpl20T+BuVCPZ1f43WdT42oxFjH
SDatpZM2UbwL9d/MJyZutNEY9PlHxSdzFacHQz0WCJO6oxSfLsbRF72O3ShVDQuP
EUlPhh4ZifnICNDM6i5pggWWOGZXJFHnCqc7vx0uH3wh3+/Ft++LnU08vS5841GN
lPcOlLZkFCD55w59ka8sS2++PQ+SxLRPXimWZMaRtMAOcQypX26hIMSxlyDX1F0e
nMysNc8qGlatSIKEjRH7AJN3SGtGH57FfrZjzPgMIc4xekbxi3kqe6B6a/9T7Rki
lvTgnUNsc3J8MQU0z8akZzeCwQYWxrEOxgB1pn3QWduQEU3o0dO8+fK+dx0+rDGf
MjzmS4sOM7mOnJyqIfccANRaehp1wkr01LcqJNzrizcy2lycZ4D+wZnNmgVQeeRK
l+MDesYAfsyTDp68/L8NuCDh9+S8qt7wfI3FXempo+JLyqhxQ6xqO59O5TTCgT4K
9gbXoG1Nb95xLBlcuVRVRXxIGgstwMPycBekSdDRnYAIgY462MtFn4sNH7VAFQNZ
wQhuGG1dK8ZRuIE3gdFmFusZtmFZQwQfr3KpVKNl5pMKE3mPQDcat63/3RQipElm
67OKr2sJft90G3jZgm5mukre1/53UOfXZ1OVyxDJo0KG2YwxxLgyoqBxqyTsEHi4
YRsK3sc2ACa/AVp1yLej5ulcLSODxgYKr233gsbpjc9ZAJQHSwBoKZFPkanmhHU+
4dwpLFSA63RFbOBcnOT3+3rxLwybZKJckE/MaH+7+xhal2Q1fau/ppPiANL3/njV
d5z4jA7gvrrQynTyyv9rEgiVnqJqI8C+i9h8v4c4t9c5FdRTasFWHHGb7OhrLu6L
P0OEX/Gh2lBIfrh09WR3CQ==
`pragma protect end_protected
