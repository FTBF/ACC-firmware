// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 03:56:36 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
F6Vwh59sd3V2VCSPb1k9eJiGR1oG5UXrzfLhA9hsmt/5sF7cqIe0FVfvr4vKF1q9
JbTeENfQak/WObD+kvIXP4UcsPM8Hz/gE6wXydsvvGpGmXYxyFPdBE8Z4Bmuv6/0
xxqCDIjiO3JRGyRqKokeyIYKZu4nvl2QMQ8SNcAInbU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12336)
X9fiqrggTMxwAcpLnBAHGQB9OX0aJDbXYdSLtW/fg8oEB+yo+cmt2743A/2oBltM
KgftVdoOx69o0pIH5EQ9Rt/qtB4aUiK9r4pAbkY2mvw8q2Aw9HvDh/BqC0d0qRqU
jmZocb8BI7QJU6YMU4BQqvLkeluASPJaHT4LDJhccjubqkFQOfJR4uwvjwyfjoEF
eIvbUilf0UgTbRFJQYBPGEd3LWy3dT2iQyENXYwZGv7d/pzSxtn0cSvcw8x9T45E
TkiSmnKoF47eVwED0Vv3SpLzYRmNKl+6fQdOsZV1uy3p06dvgAgX3J/EmXCKG8mY
AvmWLQXLE7da7qaPPEr3uytzL7q46UUst1Ig0tu6JBsSiGN6J40tR3XOLhNlg/cj
y9D8uiqi5bn649fNjfSxqzqP7SQczfByLX4y3B29WmTkGWJm3ZRWyamu++AtTdgL
pCMqP6HUQWt9K3LJcKuRVwzh7EiLYx0EcQ36Tmm2/8AStuvLSm/HawAYSGHPvQJn
Ocaw4n8CQiBOCWqWJimS2uHOVWZwGHDrOGzGtQwkl91eQha8hnb/tjxd+aKvxXay
zrzyoR7Eu0yr8rHOky892IPHZGQeOL6EU0Wt8nuXCcgc9e14xrFHv01DMB93oTOq
Ep+1r94oX1kP26ELWgIXX+WHL0kMqev8fmN3Lf7PTt+qWrx/0PhAdr+nXjZJreed
3AOJvy8kXPjiUiSbvOA9SsP1VnY7o6lpJ1EGd5FxGMbGa2gpCIcMJFAiwS6RY0j8
Q94MpoxNXZiLmjoiAnexSV87CQVStXLp8m1HWL+Lv386LaZQL2nLsDla6T9yJU06
GKh9sq+GzUgPQpjroyd5zerMy6GGUND1C9M5eXFWsHVblAqIA4dBla5jR2NEVYfG
hNubSm64NIHIQhYExbiVQD4Yan+8sJFDzsiugyiifEkSESfMMUb45irFiV4BckSx
xSJk7rMs0iDtCG/RL93Q8KP9tSi8lzrt3qJuqbybtj6XwHQie0MuhvYbkjOWUfBw
cSjW2X/PrEqnjC6ulp6hQILTvCyrRFVFkscXpzuwa9aQrZwriI3l8p0s4KuYT5T8
KHt+OFtFJXV1FaojpOha5mzF97/A9uYC4GCUNzpQCCClqxWcBtFdNxcO/FYqfMHb
HHSgY3w8jUh2m/EQb01QdH7WbxK1PTXeF5Tvanl1T88dXcPJBc9FuByzYnnIIDhQ
FgbRvIkmYr/3QVJKeoiFmMcMj07IxImvftni0KzNd8nDlob7vndsh4EBqtm0LeAl
yn53kOB18FuZvcQ7m+ldNVCN+0J3ncW0i/QpBkHax2y2TMSzX7nB8i26l7ifqXSu
f/dGoaBtyMsTqi14O0MYMy/boPSwZGNEWU6z8/vF2uCCvsI5oNUP40gp2hLwXLKU
ijFoYJE8dKa9kfCMiy8OUfZEaZ4dSdO6BBS76rAjVASv8eJ73pgmlaYNr8iFQ6dr
pHxlUmNh6AEbbJg68eemEOm1FjJwUYFEw/tIwU791lYdgivPf8YI+nDiYO1Z2C3Z
EhVmYLtW2pmSkDZplGnRiDvyW/kMHR5xoz/zz6horcazoRsgjrOQeKMFvY43Lht5
zQEbqGTneyMciuFXZ/qQi+IbR3IzXTo9VW14BKP8hvgaPldg3BijN2q6ue2/w+7G
vmGF5edBkyCz1iYHLsFMtURB5Zr1N6G1YeJ5wIOUi0ufsKHTOEAO/WCM9IADbERp
YhJb/kWwnJY75ZR2Wf1GgsgZS2hxANwvC2Z7zp7lgoilyKntas9teoER621d5Oku
Rf8L3bByaaZHwxScUWMAHVkcexVod2z6Gc41VQiMOCvCWowU/dkdvv+nbHB1jidJ
P+DLeoXrAbns0zUIdlwsiGyVp/MY6EMtQSBaNJGQyTu51/6ODsv2/8Rz4LNWIS5i
ptbybQkeFy0Z/shmBv58cZ8uO/RyTrpsYZE+mEv5Doaqg3btE1EQJd7o/2gkifuV
DihiNog8epC7fLi10ZorJx7dK2/7HeZGMxUMTtPSiPWgzMMLtPZi8ECqTFEyxDTu
tmY5N+Ou9T0vsAmKWK88O0YoTxuV2p2G+9h2p/1w7VvloigzwsTCWcl4oH50jnd1
S59iLu5yvc1YRRArz6ubI0AcWtDbHMkK4CYaKa01DOdX+UNPo2KHJyJKrIMs7EJU
8JBqBd3bD38V9Ma2uRYctEuRSTjJ06ERrA3cgyKECgrXCxXVP3PAYkgxNpwfqI3y
/K+6Up3adg2/1pXwMB+DPmmeCLFCYbSQ3A19WsV/kTHGFK/USuZ/6Labq6QdQn8q
YbuT8QUUMNULoA3lpws9la++x9ByZJKkUVSbZn+foQaex/hFAh/g9YVoQ9DUPMCs
S8vh1mES0gusaUB2qnh4DC6AOMJtZDERWQoFPUXjhPPBv8RShvBaxCk45iPSXTGr
XX7p1RS5bt4ZJ7rUbcQynntPqPKq8nN79suPd7KNgluivHCKn34Lg3yCL4KY7DpV
ir97Yrx+zPL1LNy87o9eCt1OuKomqnuvvBa74Ya1JfMDQT9IejH/2Hzx+guZ2s3X
JFcAyE8ymRkBGRJboQD+s3Rec7tBVG6yvjbUCY0li75Cms5dG6fWip6bZkEK52Hk
k+dZIbz6Y1eL7fEeiOBT1utBJLA005CcLRyNimh2hlmaJGqKE9kz3S7L/SWghGeb
fGGabSVQk+GhjW0ZTbToLirLLWU0z5AYrAITCVA5A6mGB0JNZrkaPKd+tCpaNq7k
V41bnXsf7Uoh3+Kxe1aRySaSlfXRLyFtdZa5QHWh9Vhrdcx4k1sqo1xGP20N3d+7
UYhaNzQMlTx1kJahauYtCJe0zI0pbGZZM5hQFdzsOGdPBxZBDQROFp/p3idCaz3Z
qoQ2Cj3xOoEEa9o26ZZO3ZR/s3rMiVDwfmI9LmCLOqoPuUQRUBSOh1JbXGDUAFVc
HBtdWqmBTAeWc0h4kXgRVLiApgU6kLnJ75sFXy/n1aVhCSg6Ic0xSOlaIjnE+0JL
nlJsLOUkGBvVcfyV9E/K64MYQFtSsUHQ4YaxkWyvSg1433bj0gPiOykQXoIy94eh
l/DyeR6C+UbG4KLESocd0JW34ADoN97VQtiFLfQB20Waxq720sFuGV8sIsoVFLOp
40WUjtstH/KNkOEA4GAn/5wSjJ8tOouBR2rqBTfsiMMU39XAA37HY2xktl0joNdD
sa7G5lidw/gssxnYpIr+Jb6kwN8xqarLj0dQmtQC6Yc4uqnphyBxmXLyX94/M/p1
KTJx7/6hBdSb/1WZKVwyUlSL6JGqt2FLp5c3JN9ghg3NqUAysc//ZpZVj/vL1Mb8
qweQCAMMy9T1L2Lne7pvyUhCOMzH8VyY5Kk9TvDtw8o4aAknWDHILoU+RZC8muju
l9Yvb3me5EpczAmB995Gt1NmXEwk6YOTbndLxTmUanscroN2ljcLCz1fGB/S0jKX
cOJ2URbzzvNI9axichxqgbnr78ZG1XtVLYUvgGod7efyDXqgj9CA4IUWM5caazlm
gJoiQ1gtAT8ocMp69lc8NPGh5s7O2WTPZTlz0DatXDnBdHWVyMTXSm8QIWvgg8Nw
Vhs2w1LyJCGTDlMqs5ychek0qZViKqACU2MtWgoOG9yV5GajFK4/vMW5+/RE1YXG
8OMBEEiRGOxMefIR74UMs95bvIqvIaXaUnbdgi0EYecwOW1WjYHAuEFBoOppWRkX
vw5SLognJSwsXaEABVA8liEoK8/jok8RJyam03gwJaHl6eENsVcMLMNPcCOjmkGm
WPQ+9ZNJfKcfu3ZzNJ1woe9aEGqdWyaLdDf/X95E6qTBpR/B1uZUrPrdKIi7XZ4s
DMtFw9Vh8K3kbEx0dpqel5i4m93i0SelX1Q8O270WlO8xFw3J24rmE1OihbuuFIF
iPWuz5vAZQLLR+dYl9sEJiu0P0lRKoEYhzsTPSQgN61vrTabFX/y1Qez6tlajxwB
ntnO6DHCD8uaUbKU30DT+t/ymptaRCQMpDUvgr1qRwB4Njue2DMEU2frgBOyOPPY
bvY/aKCf0FdGkRVvua+PQkpUxYEnGC4i4wrze18vamLpx+xZAh11v8pIRc9k7+qO
gY5O2BPnQFe9rYsDASVfH7JV+MZlHnDfsk9vilgxPjSMpZKZvqeqPV77bnx8gFcv
eC3+DD5/pDhu2ZuVhQuzw9qjLu4gYCrVdhksz5ru7gNZ7RqPo1oX/Bk77nCLWWS9
bgyiO+fKdpjTNOAR7vt8ft20YjorJu3TRxIVfGVXXkoEiZok8cfOcRdD4DJKx5wC
od93lplu4UpXRZuli7wMoAEr7oIVzK37w8IIOLrT+L9jVV1OZQfpzHBhkriWxYKX
ALxNxemqFS+h2BcUwLwm+EVrhnswvsrzDO3l+TfTIwyCh1RAakiuqn75oxzMCLmR
Frd5Q+hOtd3kUL1EJbhxbHpFqPeR/k01qodMN5X6RDRldFs2HzzKSV1OnAu7+zZT
IKGvstbe9fnkmzD/B7BsziAfywn+ysGxCnARByjUCy76fzYi57SaGTYE/K2Y/hE/
bAGscmVfm2vW8WsumQ/Z62lOn6KWsNy1EBQL9w/ZJF1x1U82ffE3dcouwhxAQfrg
TlARBkzl6VAAoBASw6g+iXAzIeRXcYz9lUpqrWZW6o2TZI7tdurCIbifpLMh76/C
FxxAFES7GkYed8USLIPWTdCFa7BHt1uI6s66skk5frd1FsYnXHTrr7OvHo52Lsh5
o+0P6ulRfxQ8qDKQwLFR++hDElengk1hNm4ms7iXCOpK+QzeoN4utX2/yAA8z2fa
BN+W/TUnDm5yGKEluPfL0/TtR5zBkdMaZtk6Erw0klOtWYU4Yl/YQlnZG3DEqrBe
0C/Ff6tIlq9I/r6zPmrLXVTbIkG3jw2DM6/1Rz1Nb8z/d9wHh7knubyv8gqmyIsF
2/bthqUP6EtsTAypO+txWjW1Q0S3ZYID4emBGuH5QJgdVZIvHoCsW6675OyiU4oR
ZaECPGMoYGbyQ5vx6FHx8tLCNoxyf21czl0Yw1gjUTq8w89ZslDVLfmvY8kceX8x
wYsCBNopv8zeInPuY00lZ3q5vn1vA6H66+fdC4GkzArP9ZbBRpNcZvs9xO4oLMHS
ROmLZwtCwOMBVr/4aqXM+rEo4dllOBeXsoxBfEdPYSpaokG5j1R+A8wSu74fqMcz
Vh3/GF1rLObQ4WYQ0aCEhB+XFWlnHlAy7PggNCo/6GD8Z34qlNwFJ+vQ+BOIORGn
NzfH2JgT/6fuqFfneqUboYKidGqD7D1ySbd1Wq1hGB636wnZxkQx6CnueLbivYkU
S8bFP/b8gqR3GvaN+HMYWtZpDVzWna6RfnoiB6jwZU82rcpLnC+RfxxL0kLxZu41
XtthREBJnEzXhoKcVTO4xzHOfNvJkA40MLF+HIJEpfWm49Klkh86A23hkBOes8i7
mYGzbZtu+Lq0wo/TfXgMgtsju2A4eI3S84HLNoPvlndxHCt7AZyYlJ3CR4AvPZdM
l8eK0FCRrMS+OBgtsKJRUQh7WI+AO6tzowdhyWV1izzJwhiyjUoa/6ebrpkUigJG
gvGmnNv1kErrwDC3ElxXOC2DLgJVSDNuDN1fVPnSzHZFUsPwFeo6BL/dcbc+MFCe
HBvhqxT9XPdcOktJJX3ogDiX6F5HEfZg9orNb9/qMPFrGblRO3t+nIG54sZU7RKh
M/kT9NF0xYK1xa6S0//ShKFymAV7fRy1mUe/jWzcRpiemY3trQ4OwPj33m9BtORF
uSZyXCfLkPA7PKCTrEEuSRjgq/U3gpOCJg6ZVopQjg2etx3y0CBdf4TDWpqb6+Fx
hiLm+PxpW4vM+AhS7Ec5balcwC3x5JgvpIXdlh/sOXqCjdZenV/Jamm30fa3smtP
GxXAMMK4hbMD9oN+S04H/fNz1RvpCJ1zGuiTXlxr7PFh9EeXG/fOwLFs3CcfYTCp
/dq55EGuCrriluyJS99Ui/j1Icg+PVzZiEX3BTm2Vr8Yszp81S7mF0MBr8iCjApe
xQuHB6COgAoZ1uyy0HtfZzQa/riJ63uz570GA0er3zaMSVm3s92zFSW6dDTRifXV
o9zSbKFata4NgfF1bnk5XFwKmaHRWY5iwxA90kBK9DvYPHrRuN6xoqnz9GeHaopa
iZEgW5AkHpKtCwcbn43YqjAqd6T1ChfLHpjageQ23Q0kco5QbNs0LWE29aaZkYyx
wCXNuacyiCcv1905AojiGIUIWUtUoFyE+PyAJjRLjOniOPqVvZs4ka3boUWDuYye
4iw2nHb+oGUZ4h2nXdQt0flL+mfBnugcOQru+s3M1Xmd6qMxgHCVBunDNhabjuD8
5N2pu5rxI19c1Xqb1071FfvUqgnG/HDe7ABdWrOf4dJxYZ4iSnXo3bI4MXYbxux8
L8aZl7aN6E/lD3irf4ZK4hDmrkSPLlTw5A/LGZPt9aDRXv41U+9IBQl//WI49AH/
rsNw3v3YJVo1pIqlXIIpXGsVgnda8TZOMqvwa3CpmMyqXLtFfM9y9G7ErgbpFuSn
qckA+MUid6eJ9l9dKKjs1AnoVoqB2H3DnoNCfQ11Nx3fXwyA1JRPF0SsPY+OYAN+
Kht6+E1QKGggjAZ7tNn6O/MLCuZBobapVoEd468pI68yhmCzr2c+kaWJeR9Ex5A4
98gwPaaCJjt5qxn1V6f6BIm6Ty+aoUAU+X7f3kJ07/1OPUspHPH6wwUcSeWdo01R
++bSY6blpAKkCcYyM4hx1StY4EhqBVta8kJRG7p4G+xpr03KaREreovP7e1NERNd
OyHNFAdO/9K2R/buj4ZjAxBbNAaqRuM6chhv6CPLMgxdk44M7iCn29osiry5uMjA
5T+WwDJlR/wJt2bxrgJwPeLGA3E0SiLICBlxradCIBp6vUdshqT70uUUL60OXeoa
Y2K0xOHsdK/95/ACX04h9y36yTqfnUvtT9nsK+XzZbYk1YiOrxCsFmlt+qT9kls7
tBArQcYxP/Q7tI47mOeFfKiH6zU46tIiw2HyGigayTDkNl+WMyv1oxkOoEM4deQH
KM9UzxyVr6ElX9XsNz4cTtTeN6xTPUCbOmnaOnfToYKnybr8H2C5oRRCwmOHTKvF
ACrxHkXDWB520XJejVsWyqGjvlXoJtOjSbrkRuv5CRxTChDDw8ok/3/hcCpRLayY
dUZEHoVcmLJG8bSZ6JETLDNkS4pLWrZKTPdV/arnIsgp1IOwF/87CNd6RxmFgA5L
Sv9G48TJX25RyBOKGW09NbRdDVenBZj6xh21TD4MhWR1CSvyVmVNMBiJO69I9LgC
UMvotOyH8H07Yc0hiXY72zFxnDqEStrTvIQdPITQBr1UXYfF/HOx3oks9qy8UWo4
/I+y8GBR4n9WVzlzeVHCSeEtev/swohKDDdLzomOFfhujhvkJzE564HyweL2BKew
MMB0M0/jdFy5Mi4HaEGxMhNhcRQNpM/zjwaBIRV5Og35N1PXb0BXFbCVcidKxQ1r
/wdagZ1nJ6PZ/rZkLEbdmpYH2YPu/FG0kDryC90mH4FHoNqJE9+UW3JAgHjncwxh
5bm4/BdNseASh1OpHG7ImNhPN3xU76t9UTplZryv2+WU7CTtN2ZVphieb1npEgaR
gRO3Db6RfeySulwAGTFCWOLUIOD6oFHaDNnbJeA704D0C1WREmUZAjAeTp2reI+/
XlpmL4p/0RwlMkr7zcbpgwvdAwIL8rN+NL1ZqvCHWErmrhRJbdiq6MvMCDN6wayi
1ZXkixYlpYNgBOPiQbCM1eLW1kFgbMl2VmjHYbYvR94NmWnZGjj7mq/87cGDVymP
J68SWNkfgMHDjhanH2K/pjQhINjcxV5N3QOBH8ZoLWqFXlHudpeJq50DeJEJ9QUg
kbn8uoAjVR7GA+TVOwQoexAXUKaiSizHg8l+qjuXQnVhtv89fRB9lVmJied3YFCA
fYOsRLEAZjSoXxyDKqbSEDdSxE9j5EWSFOJqckI39B/jiiJ81Fng/cB6OLRASuB+
IestwqiwLJtUbH1iChy+GkkNEGOWM4USqmv3Ez7PtsVBBx15HXdZWNYVJX4QS0Fn
RmHaA5LpSUSeoDGI7AW26gBy+jRK5BoJuJZcq8kaf7yPEAn7DhScDGxgGlzOtdIR
fTichl5Jd/Ol+QOXTC19yWadgJrowfzUBWJI4Ln4P6ZXclzWQtqYqxa2ly9cnph/
Wo5av69UpGtT+ciZWjH3RsUOb9XUxKOxDeet77bZtmbMVG3vxgJmv+VBDTB0voPe
doeJmgyrDcnIL2u7l3vAxVItv4KkfJny53MnTuXfYfQLzGsDAKTmA6qcoEvOmN8M
NJ7Q/cjTvLna/pCkKRvr9fRXzmNLIHdHs0n3HrZLDcTaPkBA0+Tk1WIDT1S2D0o+
EAbmj9KCLT+qUYa4JZesxrA9nWuedm8qxzGiDi791zreHrQfvIMXrCpAwxZtHCfa
MprKQBcKKLs1cLgEZoLK+SLtVfa+Lle5yw5IiNXD4pOrj2rSMsoIMykgO83o0Zzn
k6IMGEvs3IYdfTztAyKQS0zZ+nbJeP3Ln+qyfwaIy4gcaB49ufd2Y1YYoJ0PMD97
uCS2mHBLtggcDSPUve6zLbySMgVdR9vcIVOVDvyqg5Evqq5oIlaIczt4LxR/loRv
lFiiL7aBrbTlOQ9DlWma/FvHP2a5KgCabZPTiDDPfVRWTEybcOA2rL06SJQXXM/R
j/lPBM+r1ddSOmu1AERZZanrlHY5s4DOT2wJM+txb494gf+3CXs+HOncIxoKwP9l
sxXJuAvn2Vkm2Sge/bwOBRP4xMymctRoYDTBcmjItnhcVdNersxJFpri9rxBvze8
zaIcGKbHV9PulKnW4RjlR1SO/KZ5taikmCv/5MZMATUfFcp0Rii+hRYdiMv/R+2e
yEk+mpWm2e/d4V9GLakhwEuCJQf2GBHw1Ya1q80rdeV3jFimT2BPnfAwP5ov49U5
YFLtcOfURg8mVNRvmJEAxJUMKfOPyUvCthHzOBoalIIEr+jfC1uWjEiRUlHh+ScL
0Rb3iy1skRhvUh7o0L7tq1pE56LixXdbdm20ecc0jEmKlOl5qznpweV9p3M1V+zJ
VJe2cNDCHuoVM4vYGfKno0cqCtLuF9a+MJ7BuqPOLNsHj/GnYEs+OXffN6r+FaMI
DUgTcu7G9IRih7Slr0+5cB7bRzg/VQq+YALafCTG7ZIhU7kgPm64tir5n6tLREoo
4+/4K13kBNPO1Sxs1MkqAFL1RuLzfKWXVfMfd5D6VKvq0FVE7t4nPIjVmYubLmBm
5A1gjdQ9f/i75VtKWI8sAL2hrcIn6JkDpcqsKEREE1+B+pJMi/eID/NuBZTtXogT
0LxmFBF6lZW9xjp7UrSKDK8X967CJQm5rQ9sH9au7FPItDOZFmZqYmdxZ8090ocK
/ZbLqLrfo6ofA508p0OvGog6pUkKaUipt5WQ7LXzVWiKT7kkTsOwT45c5PDM5zSO
BmZ1HereK/V/DUx9Qt9sFMW3ZZTurlcQYhrM99bhbUQWxvRrb2abQyeyKgtUlfDR
xm9JAOM7cnTavWFqD/JczrsWinz9UedARBgEq6O9cJS08iO+XkIDGTP9/1c6sNPa
4604kYzNjDYSvd/NlM6jxej5dkL6ArsNRnUXS17uDky7Mu8ble3Oe6L1AGl4M/FZ
MXaLkUN0C7XvF6XjS/i3ImprKzlGvjMCJTBrhNL9qHGKqYRr+KWOCk6jEjFzQtCn
JyIpWzE6eHwaAFBsRJFaRg7BIegQcHA/9WI/6pyqt5nAvYgFeIkkSwrisdT/XqWp
HlNm0myz2tw2ff3WUOzmQOHWue+PvXKmF6G44OrRnB+s5SWucgxdmakIy0Xpv+TF
whKTaUVX1BaxDN6KVYBp5baYSWQ3ZkTlBiyOlPHchknYWxW+y33Vd36fNEcDZAkF
W2gdeTgP7q1tvl+GMonmyOlniHJrMEofcT6EjqcPCn2H6y89g/zZSk5raN6K6tgp
rZ4A7wj3rMtTapfp9f+TbQs5h0jbOJRFthg3VKXUQLWRyvH5Uxy46Y6UOSSR584b
NXZD4mZqn9ypI0Mn/+PAj/tYMEL93deUWk8cdXpxe3pPn+qItLvRc8qprQnb6jMA
3DciRhshPre6x2W7bcQA8F4IxeKCzpwaWkc/nq4eQSSmnyGuHLSsDwsuCMWJ11Tp
afb6CMI1ZcbEURDT/4Bu7OcTS6ZH//n+xdOUWvt+TzR2IRiUsShfwCk5iTaEvRb0
+ROGeEmcd6Fip3EeS+bEIqdJw0G3awQ3LEwNBhryxQAi74pZNvjgrlRupJ38OPoh
MdTm2csXA1Nx+H3Yf7rMZJ5xCb1FzdUDFsH4pQU3gxVuqOPsvQOz6EJxcv92w8Je
jMjAo+7KjnU8Eawm0x54KeGL3nsl2LH8zQqikMuwZkarp5Al/K0F34ntze+lcpgq
jDXu5fYND/oz7Ah7kTkkZtP+iaHtpfR3idAfFbGaqg1rJuurG0o6qENrQ2lJop/m
RhctkCbm4HsJ8nNdqfAhu6Bia9sjMW4+UA777okqDroxdVTPnMmxba797fwJEGe/
zw/dZDPFqUpg/3qm/YaxLH4eA9xnGTylhqFce+E9FWR1XscVb6So1F/LWR4/yl/q
ckwpM1AgFGp96B0twPXEhzan/lBP1aVSJX5Np6mREzr66khs6mQWdaNJ5tcjl48R
7bgvQFnVnpdS1abfG3qdyvBDGdEMTC+GnGo9J0Bs0b4TqoaxmFwLvJhVgqMY90zj
QmBynkTj4YKLCvKpAQiwc1OGhpuff790scuf4X646ij4FqpvNUzA+VM9ULE58FV+
AXLulgg0c+00vf3dZ3viMyEBRZUolfRvkRsNPQqsCDZ520XWR1YAV6e51hcbxFb3
rvm7gsDR0wkCjiuImNgmLvysdDKxplGaCC19ASTUGz96QRA7zpt8dS3mahbeUcSV
oP6DWmdDAHfDcBm0xzSeEA+XE7XQmS2S++wzcKe8kIV/jVCh79nfm00V1Gg1FHre
86xF2B+IUyFLl/Q/OCmvK2b5e7jAq1G/K2IaePemlM2Gej9cUEQ07DnzPqLHLAub
84qTnOPYYE4fjbXCFF3unl9/wEF8GkNH/LhqR05QWERDP09j5rp47RSIMapXIztL
aqYo9kJmd0Koq4MaOMFYm0khAc5qktivCvK9jX+1mzRc15pdJXTOWtX25uHywkPi
XY3lIeBIjmsdsbTsK7W5T0wPcIis9KMQeJOEz8yXxuBToUW5MZAfi5Il8rftTjeq
kKvAUxd0Hc3Rc9/mxefWa2J1rgkcxkA8BnqKjjE+EbBkInYV49k8dJbeXf3HaWoE
9GjpG4P8YAbgI18HaHqbS4L8ldDTwN3SsdZUXwj+TpoyUkdz+RJ3dHgB8PB9+PlR
5A32o1V/6DHvkQiqtLkhdcmW9GmgW39cesrFUXLxPe3n5ZkOGR+np7dBPItbBfK+
7Ab3PEwUaOaGO2wR4F/3z+i/6cPCDiTrFpDofbRmP4wx8iCws7X7MwhNXCZbBvQ8
sndbU0hK+4QyqhKmjiX1Z/iIGBcG18co7eYaZYMZ7MHMjP2MmNN0xo+EmydV4Fj/
12FOMvP9lLEuDN5BlQhWH03WNaWZ9DID/yXYbhQLmETb0BwUwqUQe5Pa+tnrDgOR
zZPR0tgyOkfvthDe0SwmuSOXpLyhN283vXL0DAKfxpmz0X2Y7bLtP7r5M9Qo4Op2
HJ1sRHXltwaxrO3xRgUFjciSBuS5Qb737NPuUQgF8nhztGtt2g/VEMrlbPYJgL6z
OP4+Hoi7paAdJV5j2iT+VniES1gtuo53zV4cgKkFq8qVi6rppLAhiopu0zoTlUgK
VQ6QzryoWkT/6ghoyiY5tqaYtGuHiBKKf3PHparTxbg5keU96hCHS2UPZTIZOMPL
qeZ+JsAWx0YlyjpWO48gjrF1Dx2HyeI0HlnFLYjZf4hbdrDbHKMMof4c5id13EQm
vBDqXg3VBNv4ZG6NfXgqObSVRJF0TVBtfQy3zUNAuHFf+7u00sUX+ku3N585Pxes
9mXI5w+4vjYEJms8OxzWOe1W0oK4AG4+dJFmMswmceW6nFggPYkrEsPOSE1PCNu1
Adaf03rSZpxYYCCZ+ideI9BSHLF4LJaoc742qFfu7revWBCrsNWjuvrjwKeNAWJ0
/VD1YVkvwNYF8G6HrbN8dEVmWvyDW9sja3iQoP3JdKXLUMNYVcfnMaTzYyNKnV6i
h/1qaPNi6SLNYjF82Cw4vfL/EPSPwspqCr8bmj3WTQrYlnZxcW3iBwYcIBBy5TRr
1C1K/3v9bG9X4RXBxSCMYESknjQScg7+JPJpaEl1c1Hpk/4X7HSFzRNKgF/ADnfU
CB0ssdVn8Ml7jcDngx8dV5tO3e81SyBkYMH4wYMSPu98BoJ1/NE4iHcOHFZ8YnQu
zqihUuoth++RPtZDG7qzM86H7eM6+qWQOH4lH6bgxC03hym0IMeAjf3BOoXMR9Yf
5E3fd0uvavrpEKHEbrQ4nbbq7xy9/nzQ9oJEW6rjLEZzgGbaM+eeLhlSwJY4QtiS
4KCzWvungsTKTz6+rgXgI9+YNoPPGHOoQ5f0dZMqqaW35Vr8ugDSviFi5xmF4Nw1
lzKXyGVWZJo8rdiTGpYl/UWkbbyscdyS11lkTA9Q0S1oFfxjkM9CSpGQcjR//98f
wtK33NuBab8lf53nm3t431LQbbMt6AL8goT2KsCX9mQ5B8HMCiOA05op3eIiSZSY
hSrR/SZXaLw4kWIVD3NhD93KN1njUyaST5whUwVGatQe/duUuJrVs3Cto9uc1F4y
JwLjo3Auz/R/RMor3otJ/MuH/1AH40QcK0jsZP3xqE1zeLrTkGu3ENgrisWAQiUk
L5HC+ww6LlSclsD7/fT7EmZzirYbve7GsEVNM48ZbF6aQqzWYZzbjR6eY/MPiby+
9mycZO2GK7SXZtgwriicOBXp3B0Bj6ewKm1AOklAQ+74/cQahpn1dIjXwd71uYaI
rgdz/uYsuDgOgZWKnydIm3hwWJ9uSB/PYwfmRfW7ZqYMatPrDLQvNUZF/XUkwS+K
HJHVvoiwOs1I4hwSbPcnLHXPPj/2L4X+rmXPYdVPwCxQigdsz5DjGW87d8sWbEb/
YUFW8iVLu3D/Pch8XkZYaAv93Q33fvl1DDWGId4ChWUHMjUI5F24aZzhO7lHI2Us
Lf/PvhEAgs4jsAwiGxe2UH4NP/t6HLJ/0O1CqmIigH0ymfqKy3Oy/ZTzFf1OyoQj
D3cm8m64qw8Xuay4g9TrUPNhr7r1NAxaECgKb3eRQHzLwjdoNWINzOQEITnevQFQ
eFzCtfRKIhYnOfgJlPXpclXHI4x5F7KJsjT2aRGMFl2UiOeyvEpf4hRHI+gtqMEZ
JAdrmrTNHqBu1p85239q/u7EekBAA2NwRdOa2zrWErzg37/zoF+UzlkQ2S4w1mWw
VrVI8e4yZ33qqfVPTtvI1PcgqLf6Ka+Z8WlryiAaKGultsqPABXMT4wIP8KzNssa
kl0JLJ5VQghiPBMBfX0UCqoGlIjUDnidGbMl9WR7Uord1dDTHEMPsdS5DEhb2k9P
jBW3czOF04PiGP983FEHbFBiQbNA87vgjCiLSorvUYVszr36O9GGEvbzSJVOS+F8
YqEMpTqtOFx5ZIAaW788FNsgEkrJjxPM/NJR/nOpMp1ooAgZhRnY/3a9t9IFK+BA
BDBLpukS0UWDxbyBkIRXZEPfs/ZdsYLkkJlZxtevk0m8KUqz8v2EyZR8lFsixlZm
dibf071qmdp2WuR8it/8WTj5Sk5OrSY97k6CCNLocVdJN0uN+JvyraZ1qClIb8o2
8KRB2Dq7UQCAjWgbmDQ1ia9GNkb5MpA1TR5dEsIfKImXvMSgjHAHFSJ5eh4J8tEU
RAzDza6MNE4YbKhN4V0+iB0UznC6BxUwPRWb25e0z0mqR2plgeJLMDHmDHssUAuy
d0tcB8AsVRUkzFb3o8HGsmKseleTBG43XEuHYR4j3cAjaY0mkXfe9qLtE0GYloLc
C3kYnnS1V+tI6u44ZNIJRIbE9XMBlk1tPtc/qSViBDtMjfsq6uQ1Fr0SmsjLb1Ee
M0SiJW8EveHtVusZFLfJCaHVHPUmKQT+Ux3C2HW9Ffayq4YbSlzqdV2JkbR9iytN
4FA9z9TfmUiftYrLAaEYf4GwjNUK/lWBTS7tHxi5CuwxqOHdHJx4owGraAyP2FEe
y2tJc1j9GM+jt5/DY4YxbXKEwd5ujv26wPN3VKm2n0JC1J7QWXt3sSqz7uvU6rs4
0DB0qqbqKlvu5bvL6kYbEg8RGpt4CQ5rkb43WY++NGtLu8vtxZvP1UA2wdosj6Ti
skj+FLelMbXxTD+0Xk/XHd7ZBdrVuNseOFDo8XFwryEDltRWeSAqxfKRD8Zjdhac
5JrSsBFViRpzftWV/qMguTmId0jwUzJ5mqTS98igAqTRco4R7w2EMl5HC7ybN8LG
lJVJgcvCg92FHiTwL4BptTR+lHebRR2sMHhNCcwF2aUxcAPznKxdEKxBMujzdTXa
QPbzBUfdnNhjKkfnLHAEuhgK7dWvRKZThkZtbteHRrpeQGD+vqU/10ilN4+pbMgI
xfQngHvLSKYs1FowceoBTPJcUVmii+gIrBDZuZlb39qoHNKtRHdO0yet8Oi5XXVY
hBPZiaw6dzpq7+7BhEkzzOGUfJpRIYhMYhF/d6Kzz3U5XWWi9PDml/Lde8qkfsT1
U+iWDvtf2JI6mYFHJp+I+0NRASQV1ImJL8StMJTuAfn9mVyVCrXKKrz4DGpgpl7r
BiwpniLEGCmBGUJmWHbIoMJDF2YU/NtEopBV7WRvTKeS3Ge1LwWPLtEoz0xpgdG3
SXnzNiHq7PMAj9+mY/iFdWQ8SZrQIuEoqbumRzzUHM1e4uLYhNloBiGaDxbYbQXs
qVvLGJwjuRbd5bdnTFI3QEFDg7W/dFHLYN59FYiXc/lG/InyOC+e+TLJ6WZBJwe2
GIAonB6PCw5LAEg5JN2xbxGgCFw+3YQ+bBP66Ba8gOegg4ymbIKouLqy4oXf3WgC
pCemy8cfaXR/vnAcjyhpt3+O2BUBtHZGYY7LOAHzmsobSSh9ZuP7kggdZQlu8srr
bQQp0GmkJpQI83vlA5rVVxDiJCet/hsGrnpll9GWbZ/2kjCEHxi1hbsXQ0wS5SL6
g3ZqhQjGZK/jUfIxX5HR4plt1CKU4WbeC0aChMtQrY3k03SEhSvwMMX+rRo++EpB
ZTLgOh0EhKAOB8lsuTXguP+IUSQCvb8XcYI/BwOIdMglIGbg74qNJOeMehhSqMcV
8IorWos2UBBcjjW4WfxDYN/QxBUfxKmBstm5t0OUjYkInzvBRfIfFXvQIqljuet6
qz/MrEfAN3cmu6wwUh2gjLvLlf4f3G3nu24akZgHND71tTckoq+41+WVQp+oQi/1
Gp/+I/q8bywIC509EuqV6u+t17Wlk3Biawpzv8D2kFUy4/2L6L86+9k8vII/NLLu
yfjT/tb6qU/mesmwa0qhFacQf44qQf6pxwjeCd+fWpPDnkLTLSgo/b9FYATsiPBZ
tMAOOghpJTdg+83x6IKgFa3UhFHsnN0ID4AeNwkOU50zTX2rD3h0AtGMDFRMSx4n
Wjv9QSh7VbascRekynhlhvTY77nnlb718C7iwGuPYcBGoD8o4+rM6lo5GpEUTApw
lyMHUzzDmDvMRlZhSD05vg9gUfccRdaRcuJnsoyLWnab0SoNsVlgLUUzMkMNQKPH
iWx8SpWdpGFNwug9ZoEN3ymntsGqlkSAAb0dhvd3tRJHYqvgeNuiKuDC6yRzhXIo
eKjh2LllNxDXvmuDaW6msduT3OxBnMo317V/YgrFsPnY9ESkeiT97B5t8prSd2fd
F8n75WgY0512yXtX7SuMGcM6ys7TzEhG7LSGq3E1JE9UxHltur2wIxI8FriWllxX
dSypM20VOsTRAuz7os6mrHinIlQ5JhI+ZBGqwohx2C87bYeDv5id46QlZXbQo2rm
niesMhoysq35HiDNuoXFF5M+EheDTgNb7tumOVwmx72S/NAJ/hL/manIfG8r2WJL
8a2CEzZ8M6iHW33Bm1qsa2IsXSYceXpDxujYe+T/uWZVLohTotbjcasvRGXixktc
u72gHy4PsL0wJlqktbrcqK7hwccTd3+zB2df4RTIcvC5rTwJFfEqQ0jMI3qpHfqr
+FBanuzkO0MHVH3hrEf7b6oebVeFIdI/2/+EEERJBp/Rl5dwxgPjEL7zShJiEw7l
SU932IHMWtgmccoJfxIbO6D+frPHVHNQ+WNMsJW6PordlkoZpNHbZJaqxMMD0dtI
hrLPM1vs89e83fxIEgcYFWv9x9Ew0IP7Q1ElRr23zcAWfipiMRx/s+Zq3C3YIlUs
DM4W7Dk5HxccQQqBj0EI0EbiX5FDS7gzCmf5NTK0Q7jNyR7uLgSSK/cHBRSwZdFo
`pragma protect end_protected
