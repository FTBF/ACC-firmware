-- clockSwitch.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity clockSwitch is
	port (
		inclk1x   : in  std_logic := '0'; --  altclkctrl_input.inclk1x
		inclk0x   : in  std_logic := '0'; --                  .inclk0x
		clkselect : in  std_logic := '0'; --                  .clkselect
		outclk    : out std_logic         -- altclkctrl_output.outclk
	);
end entity clockSwitch;

architecture rtl of clockSwitch is
	component clockSwitch_altclkctrl_0 is
		port (
			inclk1x   : in  std_logic := 'X'; -- inclk1x
			inclk0x   : in  std_logic := 'X'; -- inclk0x
			clkselect : in  std_logic := 'X'; -- clkselect
			outclk    : out std_logic         -- outclk
		);
	end component clockSwitch_altclkctrl_0;

begin

	altclkctrl_0 : component clockSwitch_altclkctrl_0
		port map (
			inclk1x   => inclk1x,   --  altclkctrl_input.inclk1x
			inclk0x   => inclk0x,   --                  .inclk0x
			clkselect => clkselect, --                  .clkselect
			outclk    => outclk     -- altclkctrl_output.outclk
		);

end architecture rtl; -- of clockSwitch
