-- eth_clk_ctrl.vhd

-- Generated using ACDS version 19.1 670

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity eth_clk_ctrl is
	port (
		inclk  : in  std_logic := '0'; --  altclkctrl_input.inclk
		outclk : out std_logic         -- altclkctrl_output.outclk
	);
end entity eth_clk_ctrl;

architecture rtl of eth_clk_ctrl is
	component eth_clk_ctrl_altclkctrl_0 is
		port (
			inclk  : in  std_logic := 'X'; -- inclk
			outclk : out std_logic         -- outclk
		);
	end component eth_clk_ctrl_altclkctrl_0;

begin

	altclkctrl_0 : component eth_clk_ctrl_altclkctrl_0
		port map (
			inclk  => inclk,  --  altclkctrl_input.inclk
			outclk => outclk  -- altclkctrl_output.outclk
		);

end architecture rtl; -- of eth_clk_ctrl
