// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 03:56:54 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
d28AX6VqxMihKcwoCAmlMRUk2yfgYloK7Su/f10BuXWK/QSPBINU2CXnLxiBeQy2
ogNiuWpvfm61n2l6qMCPwCQ8HWRkABiM5DIFX4u8Mcvaxgdj+AJXGftSLI+A8f8U
a2xPkB9JkZjP4PJY5wJlc6VTRRcFZ8KuZCcdlIGctZ0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3040)
mEkK57jhuQ4HWyXm5cQYlKYeETcPmG+65k31yvNrisC3S2Uyz///wv55wnKygoH7
MXEBwTZXfLrm+f6UZOliN6EufogrGT0nRbB48q2wXaftTEmYVmHCMrizA1Qi3/Pt
kT9dMrS6ngNHSDrb+6qZpQZxnSgSQX1+PZtdl7tBsZ3dSr6Tz5i2mMgjzk1MUQad
Mh7aufY3Zbd7Fzmw5xFpImFd7hs0qkOavGAzYT9xPqSyPeFcdtClyq4uumrBnxiw
bN1qEzdLGsm/KkhTYw/fEuouZtjaRBgyNW1sirwor4F4mqijig/2H//G5GCO3vfr
guVGi8TdnGjefety6s8ePB5vdlKduNFzpjcahRpyd8oD+RPNi21tSInQF3IBS8iM
hNznpbKuA95HPCaUA0tzfFhzBN4bzIlFXCa0FKUhjTDc2UhrGW+TBOjaRXh2KC36
d3hRUmcH9ssj0Vf8EFKKNmJgP5vYwN4YBklJwWFqNGH0xnUr/Viqh4CuJPET/glb
EpyPvXKzusBD9bd8HcCc8BVLzkL3Dr8xByBeUMypwKzE9lu9YxTFLGajUEromsQT
o94OgZDcWdenbMShrup6vPP13Kcz5RFXTU0/sdVd06U/s5sjl4z5R2/wOmNN9dqj
hTwZXkt9Sk1OrXe2GOMVz61yS4myAQcBHim1cU7eUNHi5shhvWRm+EGV2CIqJ9/z
cedYlDnBwt/zVD2lD63vXkVU/jYe0hEraA+02vhVzc+x3lxATxAYAib4P5w69U5l
9fUPD3uKs1N4GWkHwkjtqNhtzNJ6KDwakf8dUAgFCoMcN+DLSvbmSObXrt29qPyH
s1de3LKv14s1lIoiQw4lAFOyQ1L74k7gWeBfVeiNUufxVQQgYZmiDxOeiLshnAnn
NLAT3JDornRUQ+n4RumTqOac5onxBjj3bk+FeCHorK6ikwE/DzMbEstF4Z+5wnBj
maga6+T5xhrJYU5FuDzmzcJb/NE3JfUJ2EsMPn34NniPJmpHSoycq7qdShlVHDIb
39fQVZ8psAoRfSDIVyGL1nnURaubL/b7oqWxtZqO6+BO77bq8sRIRJPSXYbxy6vk
Zqd6484613nnYH1fQWstA71lOkVnPjrFM04kB1lMld/YkcXX/6yr4YlXAX0W3buW
uiVjnwKHZcnng7E7ma2IjChflHmFo+gZw6e5U1Nt0CcGklzpGFRjC+mik89OKAi0
zlTEsIWXLwmW2EzxZvOejgYe5CpyFsY29iLtIKPDXGi2KNypcfAJ+C+a8M5rEH0T
1K6b/5Gtz0DUI8XuudTGx3TtzMrwWjGv1ap5McayNWqFtqg1LtFhaWCr3U4eRUpB
tNcKrWbRcIgSPM1fRvHkhPOP0a0NhQY3BFgq+ckOFtACd8s6vbBwrUyCJo0qrcrY
UNxcy0PSZzhnsXIQmmWsJ90XgZWWemq8rHUkWQX0UOcBD3LX+IZp4dfVxey8OkYH
hEMGdBgnH6zDi45srbxCMhePej5s0VNSF6Z8HUhgIKjasBEYVoM+fj4alDM0gJCX
86m6DAfZH+Mz3/uKeRZmhCrl/3jhvV006Ep24onFLXX80OlXXAfqmVc4k3fWoxDG
JoSRJOcP6mgctjvcj9nsZBly/iSSPke2IbxQUSAi+f+VlC825npb94XBURJ+m7cH
bkI6F+zdqa9ROdg9nMD6rQm7qv108/nL+MIHGaIK662/+bvQmD/8mQUKK1bIdj8r
6WSz03BuK1plbabj77fALTQDcVK0usJzLVQaBAx29SeC2u9mxveAvvnY68So7wgw
CODeS7nkuMqCfgWwYKcAqeMFLeifgCoxt33tVUHxSVXRBszdWqBgD6Q7yrRsSSbG
vjawBwM8dNOnDVpcjJ00lX99DcCieUhGg4AeeeZXtoltuReOhhRiP/H7BxuA+Akx
vxAUlD7RmCMv+xrwFjUyQSz1+d15mA0G2r4/9dXMSJsoZqFhDtVVcMBZDzoweEgs
RUTJTM5wjgJfXNWqPh0lZcLynqpJpVFWHnTUxRsWMo4MCZ5qatJVb4qi5o/gJMvd
7UgynApzkSujPbFhNtbQs61ua9/OLJmDY+eAt3RANhv+maLC22fxjtG0SxoJ7d+X
7ZOZMkzezCoKaJLNo6EK74V1kjFh/EWHQ+cxi58Hnpsi2tkBN8BUbQ0TAOk6CCi3
mOz8Acmz40ihIhjRU5aJa/aSYIkLdGlqacYfNl8GS7TkA0WsbkBFZWSTcAUS+hYK
H5Bm0+QzLtLueSHYE3DmQn0GxwV82cOwWM5YtU2Nlj8mhYaHXKbTtVtO/mn7i8wt
BewjgoycVfkcL11BnvDhFMGPrSTzPgEv2TJaxvM+sPVrS7xkCx6dh39VIji7lnKy
jO580nLMzQCIIDqRt4hzVHiljN48Roy/TIbB0BHpSNT/tRCA8MaXR8C7At+Rm+LN
SlIcswCNySYg8oQlW0Cd0DLTgllpT7XeBKGoj0x9e3P0zzg8zpR/bXHVZSHgj+2e
S2lixkdWYgjsSa61+j9B8wnF4CKIoXdkJD3bPU+bOuxqdB+h22GC5mQuO9wvyyNM
/cQ6WSOD30f78XlzZWZFQCYlGsUdOlycQYojhlDKeIEtzRvHq5hUc5lHCzOvlhPY
pbpyMIJrf/m2jrfyWG+PMFWCOyprjrOd217bZh0YAyLpJyAgQ6g1SuDrTQA+H/1W
ThOwOgoLfPuUEZqxyG3Dl8VVf/y5dVDglKlUkzjFAUEjtX6McFS/lR7lUowjnOYg
mOiLsRHlx7PBFpx7c94ZpXnhm2+mIoP+m0dfV0q70jhznctkxSsG4yL5M5WvLFoJ
wYa5rmfj3pXC5pJLB+ZFaDLgEzFR5G9bzCVd1wz1GN1lhy3HB8vtkGUtGr2Z7IXZ
03cnzmv/undP6ScSLw/cdn7271ABv5QkJkys5etmgvyjX0K6hTTHnNNHJnt3xYEu
o6Gq1VUSPSZfw7Mp1xRScLvF3rVhi5yakxFri7MDmW28AD1Aq+mfGUNmCpbLyX0u
WzGp0XIyQlai4aRYg3S0du4fYblHCDY5OC6sh1sXSXy1aMlsCm5Ilo/YKhtxCoD7
g52Hc6P9b4k+QAvJUFRa9yv8NdYd8HbymmbaYiPa8qM5Z7UWWH2WaJR+nLb/zY9G
AySXdOZpEhYYOoy7qLYrQFpnjvrOw27AM1T3Py+b2pp+pTM5qSP1nGbVhlO9IWc4
Li6WWg2N/7dWbYtW6wNe2fGJrG7eA1z30cN9Fh86NZL9tDTvf/kHdy8VD9l+mlWY
3Z5+gRb1ZZULF2hrMnDUyUbLj7aPzC8+OPL2VA1W355uVDkkPO+nggxEMgZeER9b
F8BxzJcgPo/Qlf9PRNcYNWRq6IVZUAVwYqxgflgOhUAfe8BIJzQ77Unwbbh9srZO
QuzY40TQwYOOrjqFogCWukEcFBAXHIYMw5zZBUHLqLZKfaO8O35BCemtYJvg0vOi
3KzHqHSUb8pE0edadqPTdX3f+m8yh8jaoAFChD8huPLl74QtDqxEs/Tc3GBJLipI
3K1hC9izWucQJwwmly1UtNNGMdawXOD5CXw6M804JQ7HdHlu0ferYsErDjF3WvwT
SdvaWiZj0CCq7CbNMSUdAYgbVONRW5M6D7cGbgXyMSPRj/I1A2ql5kVeXRSo4xO/
yR6PhMvommP6BhfOOI8h4aHSA6TB4DWU39rejE/8h9EdxCtQbMBfB6BwAl0eYjVA
HECzWzSMXXWKamkvfs0mpZEwHfFcckELx51QARGbL77RxUUwvktUgTIebQxF9OIG
Gi0sy9TvPOclYPFouZgTaocbMFCL65KGn9Rnr+5LJ32sPusSU+3DEcecMXZIB9CG
9X3sujH3uW5lTW4zIYAy6hdwjmPNaKUNa60dySAX1x5gqKLqqDEazeuD5Y3PtG8Q
e2nbc842zVkjBlDQBKRpgGa7wl87IbtujRdyRFqVn1hy+iea00L5WzcD3Eu8UpXl
YPcfVGycryUwz64zR2sO+Ycq/MoHfl1LD1uUvHegcuo1qcD87LXL3OvpUl3ouZ09
ZW3A2DWYsl57ydTAK01ung==
`pragma protect end_protected
