// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:35 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kvSwxBiZVnnTxd8bK8i+3UwMK74422Lo7p1lyPg5tUBdY/u32vdXRa7E7z4A08yN
fEh+qIPUeM0IjsGqc1qazcA6Neo1NCnSKwKkGRGQ/RLMkJypkgGHZi2EOfDNYHzx
GNnrT/o8WRrSe6x4RDUg79gtBEII19IZYHNxUxoE6oo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9184)
imN9WKsYQb1MEBEkK1CFKU2WsmNB0pjl0SYjqlCMfXBl+Fdo+mAXEJiIYD4CiXwt
2Pnfg0oxFRy817/6iWop4kEG5KkGgpY+eYtxXk354W/I+gmkQ/rAoBBf0Dh1Nmi8
oIHHdcEdnbFz1llFAzvR5dc6EI35DBmW0/5jj80mnMcF8OeP0gepDFOGAnNDNjnN
2W2837NsDwf8t5t2N1sqwTKkQkitlXR7KBjj+bDhsh0fpSc9rMpjRwu+jieb3/BH
Wg6B4VjI9NFSL6/CEWT9+PN3zDNzNZkDFXG64DuHUPMEWrKEXwJOct2z1jiekdHA
vu8VlUfAp0Vcoh5lpUtV9K0wO6m9OHDqd8cFUbfuZYM+/Mi+iNqumAUYOOH/arXA
LXUnFnOB/FESoQYu5MSz7ok2U8d2g2TJYo2R+PFRN5EWXRbg/2B1SkGBlqLBr2fe
XpHj8+xXf+Ct0Vds6ppboSPQ8Sf0+LrajSzFvy2j1iXiGBE/5AigFrenSBOJqOJq
RMmAI+R3rnATD3y9H9tPWJnNe2tR/U3ltKhKpLxgbsJLw55mW1jr7Lmy3z8QN1v9
r8wRIdx18L/FngimEbvzb5H+gDcRmHZ/9z9tHO/vtCMEs7Xgf5sz4mi1VZJjhDLk
SAQQsCV/FJPAxHklR9aqx8plQ6VyyTDLbw4TfvqMu0Z3RhQCOwGErb2ERPYqJMkd
u/7wtoSRp+C9fvONMr5wc4F6nuzSid3Jyc5RcFwTKZaC7xcY9LtMnwaRAdsQZAVa
kLjMNYs1yOYVA5gThz64tzFGFNn0NwJwBiVY88ET1ftxd/GuIeX16HsYPgJWcDdp
ie2O9xte6xXM6UGM9BsMSvZ2K1ALEzvUPd6gjaVscOCun21lHM/3OmbkvFnBJr1q
iqdR+gbi/JnMmZ57tvb/ggI35ad+gpGarwY8RRAySZYYEIrWyRXdROcyBNXJ0uD+
Xy1DZV3G7a/cTbYWUhP2+CG85MJAAWK+Dkvj190/Xl/5/hQkQxAtWxrTi/czPUoN
Umx2+tm9kK7V2now4RRYT8odJIYMysJWXn+rMXKGGVkV2kHPChCefL/pwKTGCD6D
MsK8chQwRkilQgHynlEwYUox4E3FfBoJjTN9TmLke/Wp6eSSlrbfDTfpA7GcWDFP
7VO716iBEITbTRKZ1uQ/sMFTHcsmHkGNOoQmaBDlU61T2IRAZc5Cn94bWslspvz2
xy42Bt7v731fG9vGIpCRr9iMadzzyzHFwR7EoJv4HM+CVKW63m1o8yhq37IWWU/w
OcK6q8KFpDfPS/PVg5Wg7Z4+0kb9r/Rr0VFES784u+d8YJIW7kYWQLymA3zUf4QZ
SlTwdlQ7d3sWhwCPfJGIwBM5NTyz3L2sbIaMalkoElJSemSxTerpWZmWgCUpLgIT
+yrl9ZMQQn+XS+x+uHbf+HgAgpKxIA6+B+hETIT5VIWkE26JX0+YwcqThB18KnBG
NF6ZJ37/c+TWRYLditaC3XHXfrF9ywYzIHaE4yH5ylIu4cp1ggbam3neLmNCqqxS
FUTrcYI6blI4mFZ1/5+OJ9+h55AQRMBe2ZsUxVNpBS0CUw7AZiVrVa0m2l52JNfd
6XtTvKyg2kAoYZZlZoNiijObCyfmRsKPBIUCKclXO/Uz26131k1pOFt6ZOfRaWXf
zSDTG2jnZWyYgTGSkSyDhK8/rTedXgwlV1+kEjMLs1qRSGqRQ2RnA0lO02Gx6K93
5eORhhNt7h2Egb1ItinD732rGtBxN6uU1pw1/YzMvQs4OrYnnuk9IZaaMZluxRNE
appbqqb6GVQpJuaMCn7+KSrMC1c/4AOtGwZx0YW0ZV3j7buMW7/3O2LOqJC6+FD6
3ik2xlyjKwQA9RuqiqciSESVjm9RTz9XLJbVXsMhG4UkOj93JIL/luFRj5sv6STP
1ETxZGgBVp+40snFRZCarrI6OnLBtOq/66xoPOGbD3o5EnUxUw8YRf5MGConVjP+
R+Br7N+eK4cr1C/1uYUU3aY5fZK3pi955Y3QjvSQ7CDnDWO1h7KqMqkaovBH8Bpu
nqizupyg+ByGAK81Rrbes7PSxKqhrNIVlp/W70PzqEpCDJblWOWP3FLIAajaecr/
XJ86lSD1W9sJRlX2/UyFt9JQT00MI58j3znM2TOeWOea9fZMJZoq+y1x/WZazs5l
K7pf48phJTR8ecGlZ+Uawvu1OO3TeXfr6/D1GebBG0GVsBdHKIILzxu81ZlFLqpE
vzLlfWFqnrGYeMVMLIQkvjEaBANKBJ5SQkFqxrOQJNu/xroLcKIVBydG2JuZYzMH
WGDvNXQPhPjgFrODX4DG/0GJ/9n1Ng6P+5qevZRNsWPoVRQNGA6zp5AUhVfyTVVO
F1I3Pwqv+vsI15KsDPPpMhHY6Y0XPCWB8+5SzHEW3hL70AFlHoqMZ/hsokWSlETg
RoRL6ln0RrFKlWyjZDNKw6Htq8xjfbihoSwLu/NgDsKCm4+HjC9jhp4YE/7z26W/
GGml/5TqXo0Bj7NhDP9Rki8ZF+XJQnU5O6YXqZYz6hPj9LNYgEjLGqgxaZsxt/t4
yxzsZWTIdKy2RhdORIrk3iBfiSua0PPqzKciSfcSImhjOTm35lC1Uuy6dPWKd4y0
0p13+7yGT4AWlV3JEJjCINdwAy8JmdSuMY56wgRGnL+YPpV3r1MmZ19/nmVViVBo
wqz9S9W81t5zzPpCJ8Xae/8aQ0Kc6ZAcp8YjaRoJ1hTw2nxzcGwJLVu4Hobm6WCU
pBNZtmo3EOWmSARjBmjW6FoMlZldsSkaWkmUCyegv9atXMfceFPVc4TYvXcapTVj
NAOtn9D/RtvGsOsiLDnORCouWqb7PwevEetX7HFfGcl0aUXslE6rJ8qYZ/GgRial
slxoKkT62jK8nBIa7Bxfl7PzC3+NxQZRw2JvyhL28QAhWE/7HnNAUBt1btJvCVgO
bSM+1Dsym5wTLxUvPMABd55ARPljfWDL5A9e2/AFB6k+Rl5KscuTrno3JOarsJYN
kqW6WX5ro320M8koycsz9aMiGQGqL3tArBJTe/GmKmsxZ+CuFUIaXnmDRcu6cGa9
z4jfbdCgvqYddfk7wql7jM5q6UalEn+gpv3Dii/CCP8rMvFV/7PIGbzv7pQH1Kwh
RqBY0aOV/y2TbGnj8semZfcCYwxTk5l5LuvGjB54LzTj+Qt9X9mxUxv0dbzsSQbZ
YOYPjGVLMmQisNrW7IDcHnzenogkUBtigsFI9lie1t99XeVxkSM8VzOR4AWk2SKR
48m8iQjwo7VXaXaDz/5+u61Ild3B/W+6S5xWxL5XPo0zj+FOc5tUkHn5veccbeRP
6WIDBkrxKnqDFEKCylEIIwAc6215k+OElEmyEjSbhpRt/SmLd6C0T3c4vx9d7XWs
aCYDOghvQ6vC5fNeB2bpYtCI8Mhjsj8sX0VnQN0EZ0Rv+b1II1iSRGGC/j5wIQvf
3q4qPxXT6Rx4IojNlEfdLYzqrIUL2Dih+0xMfztiVvhM7oGmNahZOthPQfIpW02h
hG6YmsXg77P2r6sWUlqYYkd9EfBegBvoZZ5QhI77Aw1kbqLEYt0Bq+Tr5DXIJuCs
axGwfnXUr0/j+XsTIIxSny0+YcM665rzKcq3pvrNu6g6VKp0FzxAoNoVfTzZaCwd
FrdG6p2TrQirFj6RdQFHhNIbdysGxyeDcb/nAaw5+J2DhrKcdMDU+9LWQQvDnaKL
3Fo9/sD43T/OTvYRfvUPOBcDM/mhJwgUpg4eAlBQVPcJZ7d5THBK+i0PgXnb2OlU
yuB/gI9mTu1WClHBYrA3ABD8vo9xguCq4OVRckSLulIkmhFdDWu6gq/vU4Jl6ULH
G6NupOlwOS4uh2e0p83USm855GpcQWaaREy5QyQLWlLMX08D9u0FMwbYtgod3l7b
rOjVWsNavb8uC0C02ZzOMA8RTQu309sq71DtMeIraqhNrdWzfiAbNp+PyIZl8HzV
/axOyrJdktZWuUxZ+3rLYoFmtAW67vZjWikV1uYuS+lbOXkLLqk597J8/YpzboMT
5Ch/b/l1ndSlMRzgVU1HUtObNLXW2Y5R2vDWolqoxhdzO4o7qZxHg9V/BIbRV6+B
9u01oVt95tvDc9tIPipyt32laZWHg3gTng7bxndUtpYifrkIyAXQd3bj7EFg00iO
4z1ANjQZuF7C0tpHdjPXpXpx8+Q2nPsIimUHq6BsykHJxfXuzY20RUuHTPNlW/9A
rribdbUHr9mArh9teQbokUb7ml4Ywi7tteSMSyPRQjZyVBT1dNhcAe2k0/jZnAL5
ToHipdjXU4x2FogJW1NbgFeLr+CfkHJl1t2zHYptC/7jvVqdYchhislpGZCg2YuF
ZYwq81mR6clw7ELiMBViF9G7ZD2E2LO8cuQ8cfRXMkEKnKw9DPOFfmQwcusRN4Hu
D+D8h9ZdCZvWnS6TODC8kT9TEc3HKGIscF1fH++6pSQDwhMdiVtz/QcWPoqd4raA
jUW7vLtfAxWeOUyTUIhFaq7UBNG+g/Nfk7Wv6tj8aAiiO6FOOUZOD5kPzuIE0b8O
RgYAX7Yoz1qpuu9uNhPxTK+4GFVHqEXY2tOILOjaMzsgio+ZXlDSpkZWIxUme2ws
yUkK047YIXukuQHzaSHxKFleYa8awTgdtEKTazuw9uzTPrgCQcA+CyHaavmgtzXL
jZL6UDI+9heP19snurWm9t1DUKohqBGEuM9e5xi2I6LnfyuRrNkgBOAe+CkSZfoP
GiCEx6g0Njo4g0PfaEbW+DjlovupFpc+uYcjWWCp33p2utmsTDEbfEggH+29DRke
XGW44Eet9lzs4llDI/gNyynNYJmSNoznwR17MaITtT0tm1kczMdeFS1D6/09QdJt
47UulhSyAecjEtTIOneT1fJnsw7BPoYeY5XSlNIEYidDNqpjeCT+mMotfMY6EvAA
C3BjwaqpXlrNOY0h+xn6RzyZ5ZUAzi8Zus9aHs3yb1SW3HqQ4dPSg43dEe5y+r0m
USOJQsvzsluVecuT4Mp4OAhj82HGHzcFfDXdJCIcoNGM/vUvxqX4Pz6KEmu/NDDd
u2DomktmZlUJHIG0RrQUrw9l/kCpT5RKXlzpXrKxsfoVp7YoyUTkrTEJ4wlbltSQ
mtuHejk5SEgfOAj13GYBHTEoPVsy+dXnEkOKiyE9xQ4VVTYzluKb0i/yIclJ/eSc
Y8TH8H5Xv2pIWWAUKtEm3eclAY+++kFrPPKDuWNnuDSQbPYKOlYlws5Xwo+6cNMG
CQ8M+2W+myzzb78HJdflJntrS+J7TNyTpcLn8ivCrWVNiqbLavZxTC6amwE4gQgS
2NH7OxhFBX/FFmSSJa/vBojgB46FWQUaDfd7RLV7hyPWor2vi+DwKh9ZAz1Wjdqb
BODsD5P/np2RbBqjWfvyBsc4BOgFbT59F1jCdPstP4QAKX3jQ+nINFXULt8GsXGb
0Joi/isryz+ofQlkCxJ6H0mBcIvvXkq0v3+yRgC/uRCTAU5rwZD0SnG+5zXSeE/4
BD4o+NdHl7wh7dPcgIdYWqZvCNhcSqfv1f3ePlsDYdsG4XPi/5OCSKJqA/xCfvfH
U6PI9qkvejd95derI+v0DzfpdUrq0yP3yAPMghQb9RQNlJXTkyvlIeEg6dHUDbjt
NMithtMMKpspObDfMzg2QXSz6YTOzxMcaL+lPPqVQRZQbnKySXEYv0X+GTIOaHMp
eblSfhoN6nK78WuHA2py503mHohGzg43LJ4B1K2ScGqqSw9TFSWq1QSNhP8F4GF1
L2gUmGgNjd5oUgmqgd3ncnZdNt3J7HaFTFVZaqZC7j+9WyWpOF0H17CULtNbK/XE
mGOjf3+HOSjWDdKEqTTcyaL2flXEjPcdR1MptBID3Ys4scP8wLWCvmx4FpiuEwq2
Xn55HhpYWKzZbLnnNvoP7nL1R6PTNvx+rRF/z+oLguTSU0/6+UJC1hjwjAZEpAsV
o+wOaMIZNB7B1n4qnKVEH0E4aTU+S+zOAycB4adtxC2JtjQcPIhc0379mFgV8mFv
Pavu4kcS7vSL8j7bxdhjGwrlrGyif6hyyawHMI4XGae78SswCjgKhrp5SEBy9Ug6
/T2Wv3sm5xjqXvt7SeLNy9pLDyxLVWGKQMS/Z8Xos0GR7cPbaWyZVCoW5/WM1OFY
ZvAwiz1qGePsGbwM33HcTYXYiwuKLVZ74Kb0bxdlvAAGdSTgOaEGyqfvWRwMYcb7
c30AdelVGQUcwaRmj4Sc96BG0Z+oXobIuizU596Ao32JpH1V0nwEmB6qDLM+M+vm
lX+nw22zBrca/zEVBF98K29XV1xW1wTehMhdEmfhEKdAeINJkjWX9iujEtt+J5Il
i3nI4loPNGVFbTcw7F6pkzRedcAMdmZvdMi244I1ZXYIqEZG/uWtlFGwLfnP1AS3
xd7a0StYW6+AlJ4AYyjXtL/FlJcFoydpFYQnmU6KuYKGvPbOj1SipAKNVbrpL776
syDoWIigi31pxndd/QtL6gq9T3NkZUVu1GOguQ1ML+exI9WouSJZ2neZvuxRM6MO
vLl5MHIp/N2g0ObOhse7Wm8jQseD5lEEoIrHVdpvfVERhWH8BJcatIc/3xzSHPDC
A4+pdAiknrQ7y2BJ4gnA5e3d6H/9S/HjUmYdntRSGfs9h81/eTruKWtbrJwAmECh
egT6FqgYBm+U/DUcKGagmq3EOy2m2ZHDwd18m7oviIcpQP4gQH0HGw5Xh5rTlaiv
x2BIguNhvJSKRf/S2SOU1CIRL11agSgy6ksH+rT3CqVLyvUccpYxTJnvne0MCzo0
VegRByeJWe7BUQ4R0j+lw6WGtNbZ4oRr4vR/CdtqBXN4uTJAva+2mn8p8f7jOulz
XLco3zp+y2okGfcKTt3kM/CRa3OMIt/9QalJgOl2mk9kRTnEc7pUFrOMRTzF9eRe
n3+nwjNx9HNlAZCfBDB7CGdgqqWYSJIFVBF3Xi1aOn91c2YVT6UhFlKHXjyzbpDN
QrninTHy8h6sduBeotJSsM0Oq2hM3RqIvpllPHkJxvAZFEWCFTV5QP2CovnlHDns
DQb9PkX+/sCc0YQBqrPPOPwlr351s7VdVczsFng1kTC25loJq7y7zFpeeAXkQmpA
hcmaUZP2gmQ3+DIZSUKYRmVeeqmu4JqjINL5BJMhjicpjPa2ierUI3ItK0rEXBbS
MzfRwRY2s5Y+dm7SqagOwnSUJufoFTzFIXq4lzjv8Ef/JbbXuB8UCFqEPpREWbpo
bykQFaupYvR/cm9eg5khVfSjF5takViHoxjh3nVOfhC/V1MGeunn+NdTVrhI6rmr
4Q6uROcR4FIi8yKtHA7ySdm1B6hL5DJDXzGBVJbHazwS8eHxgvnt0CQXAeD2Uan2
CrYyTZ2mwmirnfTWaSGFo8WU7Ydg184uPX36s2nyHzQl/pnLBXqdkajkeEPVp92W
H+ix5dthTEgqTx+QMMo79w3mYNQqYdsfomA2KJdflbBGZaiPCL66AvEdTfn/TxVz
7pAGoKtaxZTyrxZ8Vv/kFhHXTPnyRRDugdsLzy9XfKwCatZzr9hC/PL8Pt/foodS
tr48lqQaa0skBlDj1pEHb+gpoLLoPJ5o5JoKO8wENEO3zYGHT8NEHzFSOTyQA2eA
QeP+bl2BRGm69VljvJr0TiibFWjJSKSHedi58niLgQabd9vSxwwNxWlE+xfSbnWO
DrO9hhEMALSFCFj3BlDzgHmds8PZ5KWJHkUUZL20BL+eLvbj/kiHxet4WntRceR1
1Zv0Q3Bjyst3b6EkmWRmvRX4yByCk5DapeyDlPB825H55bZxRSB6BAy4vOHiKTTq
4X9hRMYQc9aMvlhTEss2oAPhrG9LDTPDVwbj1pRYRlHSgFkmLBPc4IkKewpxTztF
jF0sI+sXa5DlGqqxnEBhQVAY1YDxE5ij/IBGYqgVCwFvFh0JJjqRuftlCVuEGhYc
iV6L8rQtE0JJWiupQFiMfAhS9mgwEbPHS9MlZFjFNnLFwZPvfGcm2NY51t6jvY19
IzpXIfPs6NsyDnwV0y6muc46RMHo3srGMQdNLnOSutnZMllatsWLWQLWoYDS1GpM
jM5q37GWFxebVVHirkAJChtXy2YJiouMz3k+GmYuoRqurePE50ee09rc3GGsg/HD
Omq2A6D7iGEMSGDGZNOqi+i7V4tY1ZfSa2Q8bT4EZZNYelqPnaIypzalGueOP8l+
5g83BJNB/HazaU4tZhREHxFdLbdzPnfAdUvDCUREFO7VCb+C4OG4ljF4se6SCyYd
t9+LvHw0e6TMP2LbIp14Oqc0quAF4TvyO1Pli0PyiUYFN7YuT6IsvmCs6UHhHMZa
PvIxu9+wR4vuOzJD/nIeDH/9WerhE+guWlsbFhqN6sjLomh57IY3BPdjmQNZis3z
pQwIxKIgzyLncTWkaKw5+vqhsEJuaCM1ocnhWckN47uB3hENY+fwkFg8+q1ModfD
AnKlCU3gNR3ZAwfdqfkO4pFoYE8uCRNiVupaS2ZP05QXUD0d6Skopm0Jnf4gjq2Z
HeI6jqBlkBspXF4CbeSG15BmLov829UOy74IZUi7FPR62rPZy9vCH5SE1VFywSI+
MhG6wSgsrZzWou2himgSNplmbMuqA0aUVcbKYJeORRUp18tXpYF55SBnjxiQAz68
lOCArRywLBNoWsFMmag8aBaLM0a0Ibj86uxgyigyz+P+kz6d632zh/htb7J+8V96
86kZH0E+VMTxPCS/GfU7W06Wn9IMK0hQvJVcqeEm7ajSObAxG0sn4fYOU3BteqG3
YQ35O39HBJwZgjrWuC8jOqwL0MFHWJEDeliwgAwla5MhicbGyNhjxsDGBKNG7ko9
esLCmqtgr1Oc3TnhZ4Ioi052TA9Upu3cUB79fyUD35Vcf0L42cYLswmEvfmYuSIv
5eEKmTd+yoZYmPjgkd9xuuWP52phs/aV4YRrhUz1Vdqvr6US5tg+UmRvDi5UQqcB
IkVmVCZZCAh7mJ46242RIi1xbmC8PykGD1tBsdfAciOLRF0/D8cEexlXOgQT8Wyf
Nw4SVwQiiAwiOsK3sIm8keeBhYMKJTAdEhfIrdet/O/wkpk2Iq+ZdmZ2mLRnfBNT
WrqqLI0qH/fhLOIeHQOFsz9EQuQG6bjE4MUSFzpJ5dsVQJgwrCS2E9ydoDnRFzSJ
r7AVMVl5v/jzK5d8bVspE8S1XxsZob7tq/l/2MUze/Skis/15eKYoGaKrefyTK+k
+2gwkr7fSvDV99K8rETXfSMKWZnFZ473tSK3ZJsfIQDbCNOmCqWXKiwUDC0fFKma
urTtYIOEUncGzGHzQgyXEbTBkk16Kgu3uzolWUzUz4Dzgioh9C5c86jDrvhvYndO
j1oGNJrVrpFw8OCxefFWgN+oYpMGnd7Yks7RA5wpRFz4GX7nrg0YUhBHIWhc5J1u
DGmTwtdC7hcScqv+y48rahiXmPW9yW/bux4WLdknK/uK1sTetA78PqYqlnVcvZA7
ti5+yxxQb++uGN/RA+SgEvSc+mX5yR/bT6k1TB7Wu6BWbIL7wvZRLQfsJpicfbvo
fqqS/LEA+kYvc38rqi7oDA9sXrDWuCb2n4Tzt0H8TnqG/N395z/vQxZpEsNKiaMD
2aqadlxzGEI5DgEP2edpyBAvQa13vfBG+JVesr2TIne2c73NOQ0F0xnnqvJmqtaP
RyUiH5jZHJeN0wnXzwNzT9VcdyWN7KMIvq9+apHPDWQ/YN0r2wTJzZgxP8eCcT6V
JVINbjd5jr+wbwLAvsqgbT8CSKqntQQm8f0dg1KOmxR9OyxijgCWL/G5l51OzVkh
MwZNe0WOkPsxD5LTWIW67KsLUTNrYqyn6biqz956Je2OzdPVotQ78TyqxP8p8kYJ
DuM4cKx3vDBcwjSStluTaqcfVCmaJ4p5C5pkpiK3iRQ97ylNX1WefO0HRgvDkOOx
Rlgq8ZkxmiPfp7mWnmy6HlZHieMO2xP6GqSNJUOBBYPf7mnEs6ZBQdRYHo/pSYUz
t0tUkwui6iQnHiGTcY+cR5G1MFgHqJLfVItsYZ5IIy4daUCqKF5+TOe6ctCRrPX0
l9SDxf/0tBWtMQCXWvRclT8e0UJMfHbVX3GkFgnpFgP4ePZuHtZQrwcKO3fP5UaQ
uPtAUEq03TN2z92QHA7TMFq9QmYCLjK5UQx1jEN6enI0GZC8Z5Xcq4p2xaog/mMO
q4bhnKPLtJQlztLNebFIG/uEsC1wcGuA2GlVtFbdCdS7kYbzIAXCVe/RYOJi35VU
WcqTeZaJh/DnEG65S3q3nTD8PvBlOT0IMKEykcwsGcP22Oy7pLXFePLGXMS4N7np
4CgLU+Ai3pbR71AdyJpFnFI/ckNcZzbJ6NBsgXqqEc4xmFLxTsIEEMLL/DNhs8e+
YNLpF7JPEKlj1Ga6VM8oTU7m97HQ2OI4dyw7XtU5R05TeqgalaU+l4ncUH/PrAo/
dWpa+h6VdFP2bUUpvmsRYAPCP0BPEsg5XOMv6chZ5NfYHQzXsYo9bYdcGLjjixkb
+N2DWVieO3T6NsA8QiipUpv2fpOMZT6J6KRGMk2rrg2D4vPELxmqWqzpopKVl6zo
8oP7dSRXQgHGvgl41nZl0hfJ4K7GDUmbYOFCxvg4UFPc0pwD4X6xTuA+zPlnacB4
dMDlSs8CifaMZJCAYegjBv8cFhgdvkmT3ZZa7MO2BLa9Tx4hRxeaNkgNaUXWM0Ge
AAaW7J2b10CaFiEPV7TIZsISLWbuflh4u1sWwIwLK44/qqJTnrIYTzvNXZ0tdQb9
h0w6XJMSan/5HhD+fhYVs49sFzgbA+nd0Kl/Z3WBBFAqJblsRaBILq59kXNRlKpu
KT0wSxMy3EsVu0maqTJy7GlHo9xpNtffOfUaKIOkaFBvbczQ8uOZrG7Ivw3of84d
YX1JQBUSPEfABNdvQyp5hqd7CIemiDXrLRaoBlG0OJALyqtF9jg1THfOj2TunF2y
CZI3509V6iNiyXYEcONmh4jPDMj31mrMsRYqPzh5uRBGN0fxlAOFJSLgY3Rk4mkp
pL5wdyetHhhB0RBHczcbUkYqAvSAkgPRck3WYqGBbmDn1O3Rk+7uONztnfjwFVOJ
MvHz/URNXfvL34MMLYOYfjgqo5eML25BKkZvVwNZD1J4hep1AQ+EXcB90lXVeaQb
4XTs8nl/1mwpWF6zlHOu4Dx/uq/NZGJcuyOY/nP/UfFattSP9k1P08EFBmOeOa+I
1JkDk95/zOIyAfojPYtM+MU1brXXXBQAoRra0W+s7+zDbM4p1UZU5n/u4/xGuWGl
L296iKgCw/9pjTeD/5rRKcp4GpKd8H1CIl6aRgVKERj0zI4Pc1iJKy806L+8v+Vx
H6zFa3m171vM/3/tQTzRGBGy9rzsPTR8ws9MM5Rvcm6xwCGr3C9woB1SPhZqh569
/zAO6scc3Hol7KJvN4pDlZghvXA/9/TI+qdn3bO/MfcPXeuRGDeD4dIYbdB6Ir2J
kNqWTkZvhd+p4kBJhInyXYuXkGusAjazGUWHRCXlFszf6LlPZCXhT3hvlGIUmOi2
DzyIJ/5JriLb7iBW7HDmGpuKJhfaf96JCzmVQoYs0FHQvlc/0PFa83ppFaOeqDRA
3NCeSPO7dF3IK68x9F7zLtG3aDb9ofyl4mc2Mf8vMMLtJ1VNJyDgejTx+paGRVJg
7zc6iyEUXz9oAHCPPl/mmz82NSW85xl9I6jidbq3/bVfp6BoC4mFpB5tgBZszQre
rVdjr6ZyKme3YUL4PXq/MhQLKfRrUHnE9v5DZU5OGEOpReVkTWocLslw288FgYmK
+1BsxTJje5AoamZBtBqAPG2g1QUbFuUCVNrxAFd0+C05yXB0KieO+IvqA+CrzeZM
WSrjbBtaAAFpAqRZG6PMkz05+BnqHdLOACiWSzmryUGU6v1AxM31gMrq9rbm45Lo
vFa4+R0fVBTZxAQHUGstVxh3QA33CbweAOeOwhWFIPluYe6IHG7xNlau/cGBIFKs
KL59qZECMUCTTiDj1fytH2nJHG+CulTg57O+VxEBmm4mHyq6PtWvThXw++5zUfPf
wROk/CQwNHKM7BITg5qQlUhi0KKmSOlBtaI3e28ouQwjGXBTpTC3IxHRoy0/+lJ4
UHY1+jDDpeIw55eiA95Z2iix+DNjRfRgDndmPBXwzqcJ7EQi6EliPgSMYhQp8QIT
gpGqI5TvQKbNySYLncEQn1sI22Fo1N1uWGZbWDzJmhvoZRCd3q1vXdUXF8tVO3ok
uVpGgO9wKTqAWiehsOAWJA==
`pragma protect end_protected
